magic
tech sky130B
magscale 1 2
timestamp 1717329483
<< viali >>
rect 35173 42245 35207 42279
rect 24593 42177 24627 42211
rect 25697 42177 25731 42211
rect 27169 42177 27203 42211
rect 28089 42177 28123 42211
rect 29285 42177 29319 42211
rect 30481 42177 30515 42211
rect 31677 42177 31711 42211
rect 32873 42177 32907 42211
rect 36277 42177 36311 42211
rect 37473 42177 37507 42211
rect 25513 42041 25547 42075
rect 24409 41973 24443 42007
rect 26985 41973 27019 42007
rect 27905 41973 27939 42007
rect 29101 41973 29135 42007
rect 30297 41973 30331 42007
rect 31493 41973 31527 42007
rect 32689 41973 32723 42007
rect 35265 41973 35299 42007
rect 36461 41973 36495 42007
rect 37657 41973 37691 42007
rect 1593 41565 1627 41599
rect 29285 41497 29319 41531
rect 29009 41429 29043 41463
rect 8125 41021 8159 41055
rect 9137 41021 9171 41055
rect 10057 41021 10091 41055
rect 10793 41021 10827 41055
rect 12265 41021 12299 41055
rect 13001 41021 13035 41055
rect 28733 41021 28767 41055
rect 28825 41021 28859 41055
rect 28917 41021 28951 41055
rect 29009 41021 29043 41055
rect 29285 41021 29319 41055
rect 8677 40885 8711 40919
rect 9781 40885 9815 40919
rect 10609 40885 10643 40919
rect 11345 40885 11379 40919
rect 12817 40885 12851 40919
rect 13553 40885 13587 40919
rect 28365 40885 28399 40919
rect 28549 40885 28583 40919
rect 29929 40885 29963 40919
rect 30297 40885 30331 40919
rect 12633 40681 12667 40715
rect 13277 40545 13311 40579
rect 25053 40545 25087 40579
rect 28273 40545 28307 40579
rect 30849 40545 30883 40579
rect 31309 40545 31343 40579
rect 1593 40477 1627 40511
rect 8217 40477 8251 40511
rect 8953 40477 8987 40511
rect 10425 40477 10459 40511
rect 11253 40477 11287 40511
rect 11897 40477 11931 40511
rect 14105 40477 14139 40511
rect 15117 40477 15151 40511
rect 15945 40477 15979 40511
rect 24409 40477 24443 40511
rect 24593 40477 24627 40511
rect 26893 40477 26927 40511
rect 26985 40477 27019 40511
rect 27353 40477 27387 40511
rect 27445 40477 27479 40511
rect 29101 40477 29135 40511
rect 29193 40477 29227 40511
rect 29653 40477 29687 40511
rect 30297 40477 30331 40511
rect 30481 40477 30515 40511
rect 30757 40477 30791 40511
rect 31033 40477 31067 40511
rect 31493 40477 31527 40511
rect 9597 40409 9631 40443
rect 11805 40409 11839 40443
rect 13001 40409 13035 40443
rect 14749 40409 14783 40443
rect 24225 40409 24259 40443
rect 31217 40409 31251 40443
rect 8769 40341 8803 40375
rect 10977 40341 11011 40375
rect 12541 40341 12575 40375
rect 13093 40341 13127 40375
rect 15761 40341 15795 40375
rect 16497 40341 16531 40375
rect 24777 40341 24811 40375
rect 25513 40341 25547 40375
rect 26709 40341 26743 40375
rect 27169 40341 27203 40375
rect 27629 40341 27663 40375
rect 27905 40341 27939 40375
rect 28825 40341 28859 40375
rect 29377 40341 29411 40375
rect 30205 40341 30239 40375
rect 30665 40341 30699 40375
rect 31677 40341 31711 40375
rect 8217 40137 8251 40171
rect 10425 40137 10459 40171
rect 10793 40137 10827 40171
rect 13553 40137 13587 40171
rect 15117 40137 15151 40171
rect 15485 40137 15519 40171
rect 25605 40137 25639 40171
rect 29009 40137 29043 40171
rect 30481 40137 30515 40171
rect 31217 40137 31251 40171
rect 9965 40069 9999 40103
rect 12440 40069 12474 40103
rect 24492 40069 24526 40103
rect 27874 40069 27908 40103
rect 7205 40001 7239 40035
rect 8585 40001 8619 40035
rect 22937 40001 22971 40035
rect 23949 40001 23983 40035
rect 26525 40001 26559 40035
rect 29368 40001 29402 40035
rect 30573 40001 30607 40035
rect 31401 40001 31435 40035
rect 31493 40001 31527 40035
rect 6561 39933 6595 39967
rect 8677 39933 8711 39967
rect 8769 39933 8803 39967
rect 9321 39933 9355 39967
rect 10885 39933 10919 39967
rect 10977 39933 11011 39967
rect 12173 39933 12207 39967
rect 13645 39933 13679 39967
rect 14473 39933 14507 39967
rect 15577 39933 15611 39967
rect 15669 39933 15703 39967
rect 16865 39933 16899 39967
rect 17785 39933 17819 39967
rect 23765 39933 23799 39967
rect 24225 39933 24259 39967
rect 27629 39933 27663 39967
rect 29101 39933 29135 39967
rect 26709 39865 26743 39899
rect 32413 39865 32447 39899
rect 7113 39797 7147 39831
rect 7849 39797 7883 39831
rect 14289 39797 14323 39831
rect 15025 39797 15059 39831
rect 17509 39797 17543 39831
rect 18337 39797 18371 39831
rect 22569 39797 22603 39831
rect 23673 39797 23707 39831
rect 24133 39797 24167 39831
rect 25973 39797 26007 39831
rect 26341 39797 26375 39831
rect 27261 39797 27295 39831
rect 31677 39797 31711 39831
rect 32781 39797 32815 39831
rect 8953 39593 8987 39627
rect 11253 39593 11287 39627
rect 13553 39593 13587 39627
rect 21005 39593 21039 39627
rect 28181 39593 28215 39627
rect 8769 39525 8803 39559
rect 1869 39457 1903 39491
rect 6745 39457 6779 39491
rect 7389 39457 7423 39491
rect 9505 39457 9539 39491
rect 25145 39457 25179 39491
rect 1593 39389 1627 39423
rect 6009 39389 6043 39423
rect 9321 39389 9355 39423
rect 9873 39389 9907 39423
rect 10140 39389 10174 39423
rect 11529 39389 11563 39423
rect 12173 39389 12207 39423
rect 12440 39389 12474 39423
rect 14657 39389 14691 39423
rect 16589 39389 16623 39423
rect 18153 39389 18187 39423
rect 22661 39389 22695 39423
rect 24409 39389 24443 39423
rect 25329 39389 25363 39423
rect 26065 39389 26099 39423
rect 27537 39389 27571 39423
rect 28273 39389 28307 39423
rect 29561 39389 29595 39423
rect 31033 39389 31067 39423
rect 31300 39389 31334 39423
rect 43361 39389 43395 39423
rect 3157 39321 3191 39355
rect 7297 39321 7331 39355
rect 7634 39321 7668 39355
rect 14924 39321 14958 39355
rect 16856 39321 16890 39355
rect 18981 39321 19015 39355
rect 22109 39321 22143 39355
rect 22928 39321 22962 39355
rect 26332 39321 26366 39355
rect 29806 39321 29840 39355
rect 32689 39321 32723 39355
rect 6561 39253 6595 39287
rect 9413 39253 9447 39287
rect 12081 39253 12115 39287
rect 16037 39253 16071 39287
rect 16405 39253 16439 39287
rect 17969 39253 18003 39287
rect 18705 39253 18739 39287
rect 21465 39253 21499 39287
rect 22569 39253 22603 39287
rect 24041 39253 24075 39287
rect 25053 39253 25087 39287
rect 25513 39253 25547 39287
rect 25881 39253 25915 39287
rect 27445 39253 27479 39287
rect 28917 39253 28951 39287
rect 29193 39253 29227 39287
rect 30941 39253 30975 39287
rect 32413 39253 32447 39287
rect 43545 39253 43579 39287
rect 6377 39049 6411 39083
rect 6745 39049 6779 39083
rect 8953 39049 8987 39083
rect 9413 39049 9447 39083
rect 11253 39049 11287 39083
rect 11897 39049 11931 39083
rect 12725 39049 12759 39083
rect 13093 39049 13127 39083
rect 13921 39049 13955 39083
rect 16037 39049 16071 39083
rect 18153 39049 18187 39083
rect 18521 39049 18555 39083
rect 23213 39049 23247 39083
rect 26525 39049 26559 39083
rect 27353 39049 27387 39083
rect 28825 39049 28859 39083
rect 7840 38981 7874 39015
rect 9505 38981 9539 39015
rect 10140 38981 10174 39015
rect 12265 38981 12299 39015
rect 13185 38981 13219 39015
rect 14013 38981 14047 39015
rect 14924 38981 14958 39015
rect 16948 38981 16982 39015
rect 27690 38981 27724 39015
rect 14657 38913 14691 38947
rect 16681 38913 16715 38947
rect 18981 38913 19015 38947
rect 22089 38913 22123 38947
rect 23581 38913 23615 38947
rect 23673 38913 23707 38947
rect 23857 38913 23891 38947
rect 24593 38913 24627 38947
rect 24777 38913 24811 38947
rect 24869 38913 24903 38947
rect 25145 38913 25179 38947
rect 25412 38913 25446 38947
rect 26985 38913 27019 38947
rect 27169 38913 27203 38947
rect 27445 38913 27479 38947
rect 29285 38913 29319 38947
rect 29469 38913 29503 38947
rect 30021 38913 30055 38947
rect 31217 38913 31251 38947
rect 32137 38913 32171 38947
rect 5641 38845 5675 38879
rect 6837 38845 6871 38879
rect 7021 38845 7055 38879
rect 7573 38845 7607 38879
rect 9597 38845 9631 38879
rect 9873 38845 9907 38879
rect 12357 38845 12391 38879
rect 12449 38845 12483 38879
rect 13277 38845 13311 38879
rect 14197 38845 14231 38879
rect 18613 38845 18647 38879
rect 18797 38845 18831 38879
rect 21833 38845 21867 38879
rect 24317 38845 24351 38879
rect 29193 38845 29227 38879
rect 29929 38845 29963 38879
rect 31033 38845 31067 38879
rect 31493 38845 31527 38879
rect 6193 38709 6227 38743
rect 9045 38709 9079 38743
rect 13553 38709 13587 38743
rect 16405 38709 16439 38743
rect 18061 38709 18095 38743
rect 19625 38709 19659 38743
rect 20269 38709 20303 38743
rect 20545 38709 20579 38743
rect 21281 38709 21315 38743
rect 21649 38709 21683 38743
rect 24409 38709 24443 38743
rect 30665 38709 30699 38743
rect 32781 38709 32815 38743
rect 33149 38709 33183 38743
rect 6929 38505 6963 38539
rect 10517 38505 10551 38539
rect 13645 38505 13679 38539
rect 15209 38505 15243 38539
rect 16773 38505 16807 38539
rect 17601 38505 17635 38539
rect 20177 38505 20211 38539
rect 21281 38505 21315 38539
rect 20821 38437 20855 38471
rect 21833 38437 21867 38471
rect 33701 38437 33735 38471
rect 1869 38369 1903 38403
rect 10977 38369 11011 38403
rect 11161 38369 11195 38403
rect 12265 38369 12299 38403
rect 15853 38369 15887 38403
rect 16037 38369 16071 38403
rect 17417 38369 17451 38403
rect 18153 38369 18187 38403
rect 19257 38369 19291 38403
rect 20913 38369 20947 38403
rect 22017 38369 22051 38403
rect 22293 38369 22327 38403
rect 26893 38369 26927 38403
rect 27261 38369 27295 38403
rect 28917 38369 28951 38403
rect 29285 38369 29319 38403
rect 1593 38301 1627 38335
rect 3065 38301 3099 38335
rect 4169 38301 4203 38335
rect 4905 38301 4939 38335
rect 5549 38301 5583 38335
rect 7021 38301 7055 38335
rect 7288 38301 7322 38335
rect 9045 38301 9079 38335
rect 9873 38301 9907 38335
rect 10885 38301 10919 38335
rect 11621 38301 11655 38335
rect 12521 38301 12555 38335
rect 14473 38301 14507 38335
rect 17141 38301 17175 38335
rect 18429 38301 18463 38335
rect 21097 38301 21131 38335
rect 21373 38301 21407 38335
rect 21557 38301 21591 38335
rect 22109 38301 22143 38335
rect 22201 38301 22235 38335
rect 22477 38301 22511 38335
rect 23397 38301 23431 38335
rect 24409 38301 24443 38335
rect 26157 38301 26191 38335
rect 26249 38301 26283 38335
rect 26433 38301 26467 38335
rect 27353 38301 27387 38335
rect 27537 38301 27571 38335
rect 28089 38301 28123 38335
rect 29561 38301 29595 38335
rect 30849 38301 30883 38335
rect 30941 38301 30975 38335
rect 31033 38301 31067 38335
rect 31217 38301 31251 38335
rect 31585 38301 31619 38335
rect 32321 38301 32355 38335
rect 33057 38301 33091 38335
rect 5816 38233 5850 38267
rect 15577 38233 15611 38267
rect 16681 38233 16715 38267
rect 17969 38233 18003 38267
rect 19073 38233 19107 38267
rect 19993 38233 20027 38267
rect 21741 38233 21775 38267
rect 24654 38233 24688 38267
rect 27997 38233 28031 38267
rect 30297 38233 30331 38267
rect 32137 38233 32171 38267
rect 4721 38165 4755 38199
rect 5457 38165 5491 38199
rect 8401 38165 8435 38199
rect 8769 38165 8803 38199
rect 9689 38165 9723 38199
rect 10425 38165 10459 38199
rect 12173 38165 12207 38199
rect 15117 38165 15151 38199
rect 15669 38165 15703 38199
rect 17233 38165 17267 38199
rect 18061 38165 18095 38199
rect 19901 38165 19935 38199
rect 20193 38165 20227 38199
rect 20361 38165 20395 38199
rect 22707 38165 22741 38199
rect 24041 38165 24075 38199
rect 25789 38165 25823 38199
rect 30573 38165 30607 38199
rect 32965 38165 32999 38199
rect 4629 37961 4663 37995
rect 5825 37961 5859 37995
rect 6929 37961 6963 37995
rect 9045 37961 9079 37995
rect 9505 37961 9539 37995
rect 10793 37961 10827 37995
rect 11897 37961 11931 37995
rect 15669 37961 15703 37995
rect 26065 37961 26099 37995
rect 28825 37961 28859 37995
rect 29653 37961 29687 37995
rect 30021 37961 30055 37995
rect 31585 37961 31619 37995
rect 33517 37961 33551 37995
rect 6837 37893 6871 37927
rect 7932 37893 7966 37927
rect 16957 37893 16991 37927
rect 17592 37893 17626 37927
rect 22744 37893 22778 37927
rect 25237 37893 25271 37927
rect 34253 37893 34287 37927
rect 4537 37825 4571 37859
rect 4997 37825 5031 37859
rect 5089 37825 5123 37859
rect 7573 37825 7607 37859
rect 10885 37825 10919 37859
rect 12449 37825 12483 37859
rect 12633 37825 12667 37859
rect 12981 37825 13015 37859
rect 14565 37825 14599 37859
rect 15577 37825 15611 37859
rect 16129 37825 16163 37859
rect 16221 37825 16255 37859
rect 16681 37825 16715 37859
rect 16865 37825 16899 37859
rect 17049 37825 17083 37859
rect 17325 37825 17359 37859
rect 19717 37825 19751 37859
rect 19901 37825 19935 37859
rect 19993 37825 20027 37859
rect 20453 37825 20487 37859
rect 20821 37825 20855 37859
rect 20913 37825 20947 37859
rect 25053 37825 25087 37859
rect 25329 37825 25363 37859
rect 25513 37825 25547 37859
rect 27445 37825 27479 37859
rect 27712 37825 27746 37859
rect 29837 37825 29871 37859
rect 30113 37825 30147 37859
rect 30472 37825 30506 37859
rect 33333 37825 33367 37859
rect 33793 37825 33827 37859
rect 3985 37757 4019 37791
rect 5273 37757 5307 37791
rect 5917 37757 5951 37791
rect 6101 37757 6135 37791
rect 7021 37757 7055 37791
rect 7665 37757 7699 37791
rect 9597 37757 9631 37791
rect 9781 37757 9815 37791
rect 10977 37757 11011 37791
rect 11989 37757 12023 37791
rect 12173 37757 12207 37791
rect 12725 37757 12759 37791
rect 15761 37757 15795 37791
rect 18797 37757 18831 37791
rect 20269 37757 20303 37791
rect 22477 37757 22511 37791
rect 24133 37757 24167 37791
rect 26249 37757 26283 37791
rect 27261 37757 27295 37791
rect 28917 37757 28951 37791
rect 30205 37757 30239 37791
rect 32137 37757 32171 37791
rect 33609 37757 33643 37791
rect 9137 37689 9171 37723
rect 17233 37689 17267 37723
rect 19533 37689 19567 37723
rect 22385 37689 22419 37723
rect 23857 37689 23891 37723
rect 24869 37689 24903 37723
rect 32781 37689 32815 37723
rect 5457 37621 5491 37655
rect 6469 37621 6503 37655
rect 10241 37621 10275 37655
rect 10425 37621 10459 37655
rect 11529 37621 11563 37655
rect 12541 37621 12575 37655
rect 14105 37621 14139 37655
rect 15117 37621 15151 37655
rect 15209 37621 15243 37655
rect 16405 37621 16439 37655
rect 18705 37621 18739 37655
rect 19441 37621 19475 37655
rect 20637 37621 20671 37655
rect 21557 37621 21591 37655
rect 24777 37621 24811 37655
rect 26801 37621 26835 37655
rect 29561 37621 29595 37655
rect 31861 37621 31895 37655
rect 33149 37621 33183 37655
rect 33977 37621 34011 37655
rect 5549 37417 5583 37451
rect 7297 37417 7331 37451
rect 8769 37417 8803 37451
rect 11253 37417 11287 37451
rect 13829 37417 13863 37451
rect 14289 37417 14323 37451
rect 14473 37417 14507 37451
rect 33609 37417 33643 37451
rect 17509 37349 17543 37383
rect 19073 37349 19107 37383
rect 20361 37349 20395 37383
rect 27353 37349 27387 37383
rect 6745 37281 6779 37315
rect 9505 37281 9539 37315
rect 11989 37281 12023 37315
rect 12817 37281 12851 37315
rect 13553 37281 13587 37315
rect 13645 37281 13679 37315
rect 14657 37281 14691 37315
rect 16865 37281 16899 37315
rect 19349 37281 19383 37315
rect 19993 37281 20027 37315
rect 21281 37281 21315 37315
rect 21465 37281 21499 37315
rect 22937 37281 22971 37315
rect 23857 37281 23891 37315
rect 24777 37281 24811 37315
rect 24869 37281 24903 37315
rect 31769 37281 31803 37315
rect 1593 37213 1627 37247
rect 4169 37213 4203 37247
rect 7389 37213 7423 37247
rect 9873 37213 9907 37247
rect 11713 37213 11747 37247
rect 12633 37213 12667 37247
rect 13185 37213 13219 37247
rect 13277 37213 13311 37247
rect 13737 37213 13771 37247
rect 14924 37213 14958 37247
rect 16681 37213 16715 37247
rect 17693 37213 17727 37247
rect 17960 37213 17994 37247
rect 20177 37213 20211 37247
rect 22109 37213 22143 37247
rect 22201 37213 22235 37247
rect 22385 37213 22419 37247
rect 23950 37213 23984 37247
rect 24041 37213 24075 37247
rect 24133 37213 24167 37247
rect 24961 37213 24995 37247
rect 25053 37213 25087 37247
rect 25237 37213 25271 37247
rect 26801 37213 26835 37247
rect 27721 37213 27755 37247
rect 27988 37213 28022 37247
rect 29745 37213 29779 37247
rect 31033 37213 31067 37247
rect 31125 37213 31159 37247
rect 31309 37213 31343 37247
rect 31953 37213 31987 37247
rect 32220 37213 32254 37247
rect 2329 37145 2363 37179
rect 4436 37145 4470 37179
rect 6561 37145 6595 37179
rect 7656 37145 7690 37179
rect 9321 37145 9355 37179
rect 10140 37145 10174 37179
rect 14105 37145 14139 37179
rect 14321 37145 14355 37179
rect 16773 37145 16807 37179
rect 17141 37145 17175 37179
rect 22845 37145 22879 37179
rect 25504 37145 25538 37179
rect 3157 37077 3191 37111
rect 6101 37077 6135 37111
rect 6193 37077 6227 37111
rect 6653 37077 6687 37111
rect 8953 37077 8987 37111
rect 9413 37077 9447 37111
rect 11345 37077 11379 37111
rect 11805 37077 11839 37111
rect 12173 37077 12207 37111
rect 12541 37077 12575 37111
rect 13001 37077 13035 37111
rect 16037 37077 16071 37111
rect 19901 37077 19935 37111
rect 20821 37077 20855 37111
rect 21189 37077 21223 37111
rect 23581 37077 23615 37111
rect 23673 37077 23707 37111
rect 24593 37077 24627 37111
rect 26617 37077 26651 37111
rect 29101 37077 29135 37111
rect 30297 37077 30331 37111
rect 30573 37077 30607 37111
rect 33333 37077 33367 37111
rect 5549 36873 5583 36907
rect 6377 36873 6411 36907
rect 7941 36873 7975 36907
rect 8309 36873 8343 36907
rect 8769 36873 8803 36907
rect 11989 36873 12023 36907
rect 18153 36873 18187 36907
rect 18521 36873 18555 36907
rect 28733 36873 28767 36907
rect 31401 36873 31435 36907
rect 33149 36873 33183 36907
rect 33425 36873 33459 36907
rect 4436 36805 4470 36839
rect 6837 36805 6871 36839
rect 11897 36805 11931 36839
rect 14933 36805 14967 36839
rect 17233 36805 17267 36839
rect 20729 36805 20763 36839
rect 24777 36805 24811 36839
rect 3525 36737 3559 36771
rect 4169 36737 4203 36771
rect 6745 36737 6779 36771
rect 7205 36737 7239 36771
rect 7849 36737 7883 36771
rect 8677 36737 8711 36771
rect 9781 36737 9815 36771
rect 10048 36737 10082 36771
rect 12541 36737 12575 36771
rect 14105 36737 14139 36771
rect 14749 36737 14783 36771
rect 15025 36737 15059 36771
rect 15209 36737 15243 36771
rect 15485 36737 15519 36771
rect 15577 36737 15611 36771
rect 15945 36737 15979 36771
rect 17141 36737 17175 36771
rect 17601 36737 17635 36771
rect 18981 36737 19015 36771
rect 19165 36737 19199 36771
rect 20085 36737 20119 36771
rect 22201 36737 22235 36771
rect 22293 36737 22327 36771
rect 22477 36737 22511 36771
rect 23121 36737 23155 36771
rect 24133 36737 24167 36771
rect 24961 36737 24995 36771
rect 25228 36737 25262 36771
rect 26433 36737 26467 36771
rect 26617 36737 26651 36771
rect 27261 36737 27295 36771
rect 27353 36737 27387 36771
rect 27445 36737 27479 36771
rect 27629 36737 27663 36771
rect 27905 36737 27939 36771
rect 28089 36737 28123 36771
rect 28181 36737 28215 36771
rect 28641 36737 28675 36771
rect 29377 36737 29411 36771
rect 29469 36737 29503 36771
rect 29561 36737 29595 36771
rect 29745 36737 29779 36771
rect 30021 36737 30055 36771
rect 30288 36737 30322 36771
rect 32781 36737 32815 36771
rect 6929 36669 6963 36703
rect 8033 36669 8067 36703
rect 8953 36669 8987 36703
rect 12081 36669 12115 36703
rect 13277 36669 13311 36703
rect 17233 36669 17267 36703
rect 18613 36669 18647 36703
rect 18705 36669 18739 36703
rect 19257 36669 19291 36703
rect 21465 36669 21499 36703
rect 22937 36669 22971 36703
rect 23949 36669 23983 36703
rect 26985 36669 27019 36703
rect 27721 36669 27755 36703
rect 28825 36669 28859 36703
rect 32137 36669 32171 36703
rect 11161 36601 11195 36635
rect 14749 36601 14783 36635
rect 16405 36601 16439 36635
rect 17785 36601 17819 36635
rect 26341 36601 26375 36635
rect 26801 36601 26835 36635
rect 4077 36533 4111 36567
rect 6101 36533 6135 36567
rect 7297 36533 7331 36567
rect 7481 36533 7515 36567
rect 9597 36533 9631 36567
rect 11529 36533 11563 36567
rect 13185 36533 13219 36567
rect 13921 36533 13955 36567
rect 14657 36533 14691 36567
rect 19073 36533 19107 36567
rect 19901 36533 19935 36567
rect 20637 36533 20671 36567
rect 28273 36533 28307 36567
rect 29101 36533 29135 36567
rect 31769 36533 31803 36567
rect 5089 36329 5123 36363
rect 10977 36329 11011 36363
rect 11805 36329 11839 36363
rect 13369 36329 13403 36363
rect 19257 36329 19291 36363
rect 22477 36329 22511 36363
rect 24501 36329 24535 36363
rect 27537 36329 27571 36363
rect 8953 36261 8987 36295
rect 15117 36261 15151 36295
rect 24133 36261 24167 36295
rect 5641 36193 5675 36227
rect 10425 36193 10459 36227
rect 11253 36193 11287 36227
rect 11989 36193 12023 36227
rect 14749 36193 14783 36227
rect 15669 36193 15703 36227
rect 16681 36193 16715 36227
rect 19809 36193 19843 36227
rect 22753 36193 22787 36227
rect 25881 36193 25915 36227
rect 26709 36193 26743 36227
rect 26893 36193 26927 36227
rect 28457 36193 28491 36227
rect 28549 36193 28583 36227
rect 29009 36193 29043 36227
rect 29184 36193 29218 36227
rect 29285 36193 29319 36227
rect 29561 36193 29595 36227
rect 33149 36193 33183 36227
rect 1593 36125 1627 36159
rect 4445 36125 4479 36159
rect 5457 36125 5491 36159
rect 6009 36125 6043 36159
rect 6745 36125 6779 36159
rect 7481 36125 7515 36159
rect 8125 36125 8159 36159
rect 9229 36125 9263 36159
rect 9321 36125 9355 36159
rect 9413 36125 9447 36159
rect 9597 36125 9631 36159
rect 10241 36125 10275 36159
rect 12256 36125 12290 36159
rect 13645 36125 13679 36159
rect 13921 36125 13955 36159
rect 14565 36125 14599 36159
rect 15577 36125 15611 36159
rect 16037 36125 16071 36159
rect 17601 36125 17635 36159
rect 17693 36125 17727 36159
rect 17877 36125 17911 36159
rect 17969 36125 18003 36159
rect 18521 36125 18555 36159
rect 19717 36125 19751 36159
rect 20269 36125 20303 36159
rect 21833 36125 21867 36159
rect 24685 36125 24719 36159
rect 25053 36125 25087 36159
rect 26525 36125 26559 36159
rect 29101 36125 29135 36159
rect 31033 36125 31067 36159
rect 5549 36057 5583 36091
rect 8033 36057 8067 36091
rect 14473 36057 14507 36091
rect 15485 36057 15519 36091
rect 16589 36057 16623 36091
rect 20536 36057 20570 36091
rect 23020 36057 23054 36091
rect 25605 36057 25639 36091
rect 25697 36057 25731 36091
rect 29828 36057 29862 36091
rect 31677 36057 31711 36091
rect 32321 36057 32355 36091
rect 4997 35989 5031 36023
rect 6561 35989 6595 36023
rect 7297 35989 7331 36023
rect 8769 35989 8803 36023
rect 13461 35989 13495 36023
rect 13829 35989 13863 36023
rect 14105 35989 14139 36023
rect 17325 35989 17359 36023
rect 17417 35989 17451 36023
rect 18245 35989 18279 36023
rect 19073 35989 19107 36023
rect 19625 35989 19659 36023
rect 21649 35989 21683 36023
rect 25237 35989 25271 36023
rect 26065 35989 26099 36023
rect 26433 35989 26467 36023
rect 27813 35989 27847 36023
rect 27997 35989 28031 36023
rect 28365 35989 28399 36023
rect 28825 35989 28859 36023
rect 30941 35989 30975 36023
rect 31953 35989 31987 36023
rect 32689 35989 32723 36023
rect 4629 35785 4663 35819
rect 6377 35785 6411 35819
rect 6745 35785 6779 35819
rect 8033 35785 8067 35819
rect 8401 35785 8435 35819
rect 8861 35785 8895 35819
rect 12541 35785 12575 35819
rect 12633 35785 12667 35819
rect 13001 35785 13035 35819
rect 19901 35785 19935 35819
rect 21557 35785 21591 35819
rect 23213 35785 23247 35819
rect 23765 35785 23799 35819
rect 25329 35785 25363 35819
rect 25697 35785 25731 35819
rect 28641 35785 28675 35819
rect 29285 35785 29319 35819
rect 33057 35785 33091 35819
rect 5825 35717 5859 35751
rect 7573 35717 7607 35751
rect 7665 35717 7699 35751
rect 11805 35717 11839 35751
rect 13093 35717 13127 35751
rect 14565 35717 14599 35751
rect 15016 35717 15050 35751
rect 17693 35717 17727 35751
rect 18429 35717 18463 35751
rect 20444 35717 20478 35751
rect 22100 35717 22134 35751
rect 27445 35717 27479 35751
rect 29101 35717 29135 35751
rect 32781 35717 32815 35751
rect 3985 35649 4019 35683
rect 4537 35649 4571 35683
rect 4997 35649 5031 35683
rect 6837 35649 6871 35683
rect 9137 35649 9171 35683
rect 9229 35649 9263 35683
rect 9326 35649 9360 35683
rect 9505 35649 9539 35683
rect 9597 35649 9631 35683
rect 9781 35649 9815 35683
rect 11161 35649 11195 35683
rect 11897 35649 11931 35683
rect 13737 35649 13771 35683
rect 14749 35649 14783 35683
rect 17877 35649 17911 35683
rect 18153 35649 18187 35683
rect 18788 35649 18822 35683
rect 20177 35649 20211 35683
rect 21833 35649 21867 35683
rect 23673 35649 23707 35683
rect 24317 35649 24351 35683
rect 25145 35649 25179 35683
rect 25513 35649 25547 35683
rect 25789 35649 25823 35683
rect 26065 35649 26099 35683
rect 27261 35649 27295 35683
rect 28273 35649 28307 35683
rect 28457 35649 28491 35683
rect 29653 35649 29687 35683
rect 30481 35649 30515 35683
rect 30748 35649 30782 35683
rect 5089 35581 5123 35615
rect 5273 35581 5307 35615
rect 5917 35581 5951 35615
rect 6101 35581 6135 35615
rect 7021 35581 7055 35615
rect 7849 35581 7883 35615
rect 8493 35581 8527 35615
rect 8677 35581 8711 35615
rect 10977 35581 11011 35615
rect 13277 35581 13311 35615
rect 16957 35581 16991 35615
rect 17509 35581 17543 35615
rect 18521 35581 18555 35615
rect 23949 35581 23983 35615
rect 24961 35581 24995 35615
rect 25881 35581 25915 35615
rect 26617 35581 26651 35615
rect 27077 35581 27111 35615
rect 27537 35581 27571 35615
rect 29377 35581 29411 35615
rect 29561 35581 29595 35615
rect 32137 35581 32171 35615
rect 10885 35513 10919 35547
rect 17601 35513 17635 35547
rect 23305 35513 23339 35547
rect 25513 35513 25547 35547
rect 31861 35513 31895 35547
rect 5457 35445 5491 35479
rect 7205 35445 7239 35479
rect 9965 35445 9999 35479
rect 10517 35445 10551 35479
rect 11345 35445 11379 35479
rect 16129 35445 16163 35479
rect 16497 35445 16531 35479
rect 24869 35445 24903 35479
rect 26249 35445 26283 35479
rect 28181 35445 28215 35479
rect 28825 35445 28859 35479
rect 29837 35445 29871 35479
rect 3617 35241 3651 35275
rect 5641 35241 5675 35275
rect 7113 35241 7147 35275
rect 9597 35241 9631 35275
rect 10425 35241 10459 35275
rect 10609 35241 10643 35275
rect 11437 35241 11471 35275
rect 12725 35241 12759 35275
rect 12909 35241 12943 35275
rect 13921 35241 13955 35275
rect 16221 35241 16255 35275
rect 19073 35241 19107 35275
rect 23213 35241 23247 35275
rect 24869 35241 24903 35275
rect 25237 35241 25271 35275
rect 30389 35241 30423 35275
rect 32229 35241 32263 35275
rect 7481 35173 7515 35207
rect 7665 35173 7699 35207
rect 12633 35173 12667 35207
rect 17417 35173 17451 35207
rect 23581 35173 23615 35207
rect 24593 35173 24627 35207
rect 25973 35173 26007 35207
rect 27905 35173 27939 35207
rect 32505 35173 32539 35207
rect 8585 35105 8619 35139
rect 8953 35105 8987 35139
rect 9781 35105 9815 35139
rect 11253 35105 11287 35139
rect 13093 35105 13127 35139
rect 17141 35105 17175 35139
rect 28917 35105 28951 35139
rect 29009 35105 29043 35139
rect 29561 35105 29595 35139
rect 31033 35105 31067 35139
rect 31769 35105 31803 35139
rect 1593 35037 1627 35071
rect 4261 35037 4295 35071
rect 5733 35037 5767 35071
rect 7573 35037 7607 35071
rect 7757 35037 7791 35071
rect 9873 35037 9907 35071
rect 10333 35037 10367 35071
rect 10517 35037 10551 35071
rect 11713 35037 11747 35071
rect 11805 35037 11839 35071
rect 11897 35037 11931 35071
rect 12081 35037 12115 35071
rect 12817 35037 12851 35071
rect 13185 35037 13219 35071
rect 13369 35037 13403 35071
rect 13553 35037 13587 35071
rect 13645 35037 13679 35071
rect 13737 35037 13771 35071
rect 14105 35037 14139 35071
rect 15577 35037 15611 35071
rect 17785 35037 17819 35071
rect 18521 35037 18555 35071
rect 19257 35037 19291 35071
rect 20085 35037 20119 35071
rect 21005 35037 21039 35071
rect 21097 35037 21131 35071
rect 21189 35037 21223 35071
rect 21373 35037 21407 35071
rect 22477 35037 22511 35071
rect 22753 35037 22787 35071
rect 23121 35037 23155 35071
rect 23305 35037 23339 35071
rect 24133 35037 24167 35071
rect 24409 35037 24443 35071
rect 25421 35037 25455 35071
rect 25605 35037 25639 35071
rect 25881 35037 25915 35071
rect 26065 35037 26099 35071
rect 26617 35037 26651 35071
rect 27077 35037 27111 35071
rect 27905 35037 27939 35071
rect 28089 35037 28123 35071
rect 29745 35037 29779 35071
rect 30205 35037 30239 35071
rect 31125 35037 31159 35071
rect 31309 35037 31343 35071
rect 31953 35037 31987 35071
rect 32045 35037 32079 35071
rect 4528 34969 4562 35003
rect 6000 34969 6034 35003
rect 7849 34969 7883 35003
rect 11069 34969 11103 35003
rect 12265 34969 12299 35003
rect 14372 34969 14406 35003
rect 20637 34969 20671 35003
rect 21833 34969 21867 35003
rect 22201 34969 22235 35003
rect 25789 34969 25823 35003
rect 26801 34969 26835 35003
rect 27721 34969 27755 35003
rect 30021 34969 30055 35003
rect 3249 34901 3283 34935
rect 4169 34901 4203 34935
rect 10241 34901 10275 34935
rect 10977 34901 11011 34935
rect 13185 34901 13219 34935
rect 15485 34901 15519 34935
rect 16497 34901 16531 34935
rect 16865 34901 16899 34935
rect 16957 34901 16991 34935
rect 19901 34901 19935 34935
rect 20729 34901 20763 34935
rect 22293 34901 22327 34935
rect 22661 34901 22695 34935
rect 26985 34901 27019 34935
rect 28457 34901 28491 34935
rect 28825 34901 28859 34935
rect 29929 34901 29963 34935
rect 32873 34901 32907 34935
rect 4169 34697 4203 34731
rect 7757 34697 7791 34731
rect 8125 34697 8159 34731
rect 11805 34697 11839 34731
rect 12817 34697 12851 34731
rect 13185 34697 13219 34731
rect 14933 34697 14967 34731
rect 15301 34697 15335 34731
rect 16405 34697 16439 34731
rect 18245 34697 18279 34731
rect 21649 34697 21683 34731
rect 22201 34697 22235 34731
rect 22937 34697 22971 34731
rect 25881 34697 25915 34731
rect 28365 34697 28399 34731
rect 29285 34697 29319 34731
rect 31769 34697 31803 34731
rect 32321 34697 32355 34731
rect 9597 34629 9631 34663
rect 13001 34629 13035 34663
rect 14197 34629 14231 34663
rect 15025 34629 15059 34663
rect 20260 34629 20294 34663
rect 22017 34629 22051 34663
rect 24777 34629 24811 34663
rect 27252 34629 27286 34663
rect 29644 34629 29678 34663
rect 25007 34595 25041 34629
rect 4261 34561 4295 34595
rect 4528 34561 4562 34595
rect 6377 34561 6411 34595
rect 6644 34561 6678 34595
rect 8401 34561 8435 34595
rect 9505 34561 9539 34595
rect 9873 34561 9907 34595
rect 9965 34561 9999 34595
rect 10057 34561 10091 34595
rect 10241 34561 10275 34595
rect 11897 34561 11931 34595
rect 12081 34561 12115 34595
rect 12173 34561 12207 34595
rect 12265 34561 12299 34595
rect 12633 34561 12667 34595
rect 12909 34561 12943 34595
rect 13277 34561 13311 34595
rect 13645 34561 13679 34595
rect 13829 34561 13863 34595
rect 15209 34561 15243 34595
rect 16221 34561 16255 34595
rect 16497 34561 16531 34595
rect 16865 34561 16899 34595
rect 17132 34561 17166 34595
rect 19257 34561 19291 34595
rect 19625 34561 19659 34595
rect 19993 34561 20027 34595
rect 21465 34561 21499 34595
rect 21649 34561 21683 34595
rect 21833 34561 21867 34595
rect 23489 34561 23523 34595
rect 25329 34561 25363 34595
rect 25421 34561 25455 34595
rect 26341 34561 26375 34595
rect 26617 34561 26651 34595
rect 26801 34561 26835 34595
rect 26985 34561 27019 34595
rect 28641 34561 28675 34595
rect 30849 34561 30883 34595
rect 1777 34493 1811 34527
rect 2145 34493 2179 34527
rect 2697 34493 2731 34527
rect 2881 34493 2915 34527
rect 3525 34493 3559 34527
rect 8309 34493 8343 34527
rect 8861 34493 8895 34527
rect 9229 34493 9263 34527
rect 9321 34493 9355 34527
rect 13461 34493 13495 34527
rect 14289 34493 14323 34527
rect 16037 34493 16071 34527
rect 18613 34493 18647 34527
rect 19165 34493 19199 34527
rect 19717 34493 19751 34527
rect 22385 34493 22419 34527
rect 23213 34493 23247 34527
rect 23305 34493 23339 34527
rect 23397 34493 23431 34527
rect 23949 34493 23983 34527
rect 28457 34493 28491 34527
rect 29377 34493 29411 34527
rect 6193 34425 6227 34459
rect 8769 34425 8803 34459
rect 11989 34425 12023 34459
rect 13369 34425 13403 34459
rect 21373 34425 21407 34459
rect 25513 34425 25547 34459
rect 26433 34425 26467 34459
rect 26525 34425 26559 34459
rect 28825 34425 28859 34459
rect 30757 34425 30791 34459
rect 3433 34357 3467 34391
rect 5641 34357 5675 34391
rect 10517 34357 10551 34391
rect 10977 34357 11011 34391
rect 11345 34357 11379 34391
rect 12449 34357 12483 34391
rect 13001 34357 13035 34391
rect 15945 34357 15979 34391
rect 23029 34357 23063 34391
rect 24501 34357 24535 34391
rect 24961 34357 24995 34391
rect 25145 34357 25179 34391
rect 26157 34357 26191 34391
rect 31493 34357 31527 34391
rect 2697 34153 2731 34187
rect 4261 34153 4295 34187
rect 8401 34153 8435 34187
rect 8677 34153 8711 34187
rect 9413 34153 9447 34187
rect 9597 34153 9631 34187
rect 10149 34153 10183 34187
rect 11161 34153 11195 34187
rect 11805 34153 11839 34187
rect 25145 34153 25179 34187
rect 26709 34153 26743 34187
rect 29285 34153 29319 34187
rect 31401 34153 31435 34187
rect 4997 34085 5031 34119
rect 5089 34085 5123 34119
rect 9229 34085 9263 34119
rect 13645 34085 13679 34119
rect 17141 34085 17175 34119
rect 20637 34085 20671 34119
rect 3341 34017 3375 34051
rect 4445 34017 4479 34051
rect 5641 34017 5675 34051
rect 6469 34017 6503 34051
rect 6653 34017 6687 34051
rect 8125 34017 8159 34051
rect 10885 34017 10919 34051
rect 11253 34017 11287 34051
rect 11713 34017 11747 34051
rect 13277 34017 13311 34051
rect 15301 34017 15335 34051
rect 15853 34017 15887 34051
rect 18613 34017 18647 34051
rect 20821 34017 20855 34051
rect 24685 34017 24719 34051
rect 27997 34017 28031 34051
rect 29929 34017 29963 34051
rect 30665 34017 30699 34051
rect 30941 34017 30975 34051
rect 1593 33949 1627 33983
rect 2053 33949 2087 33983
rect 5549 33949 5583 33983
rect 6837 33949 6871 33983
rect 8033 33949 8067 33983
rect 8953 33949 8987 33983
rect 9505 33949 9539 33983
rect 9689 33949 9723 33983
rect 10977 33949 11011 33983
rect 11069 33949 11103 33983
rect 11989 33949 12023 33983
rect 12081 33949 12115 33983
rect 12173 33949 12207 33983
rect 12265 33949 12299 33983
rect 12449 33949 12483 33983
rect 12633 33949 12667 33983
rect 12909 33949 12943 33983
rect 13093 33949 13127 33983
rect 13185 33949 13219 33983
rect 13461 33949 13495 33983
rect 14105 33949 14139 33983
rect 14289 33949 14323 33983
rect 14565 33949 14599 33983
rect 14933 33949 14967 33983
rect 15485 33949 15519 33983
rect 15945 33949 15979 33983
rect 17417 33949 17451 33983
rect 17509 33949 17543 33983
rect 17601 33949 17635 33983
rect 17785 33949 17819 33983
rect 18521 33949 18555 33983
rect 18889 33949 18923 33983
rect 18981 33949 19015 33983
rect 19257 33949 19291 33983
rect 19625 33949 19659 33983
rect 20269 33949 20303 33983
rect 21465 33949 21499 33983
rect 22661 33949 22695 33983
rect 22845 33949 22879 33983
rect 23112 33949 23146 33983
rect 24409 33949 24443 33983
rect 24581 33949 24615 33983
rect 24777 33949 24811 33983
rect 24961 33949 24995 33983
rect 25329 33949 25363 33983
rect 26157 33949 26191 33983
rect 26249 33949 26283 33983
rect 26617 33949 26651 33983
rect 26985 33949 27019 33983
rect 27077 33949 27111 33983
rect 27169 33949 27203 33983
rect 27353 33949 27387 33983
rect 28089 33949 28123 33983
rect 28457 33949 28491 33983
rect 28733 33949 28767 33983
rect 28917 33949 28951 33983
rect 29101 33949 29135 33983
rect 30021 33949 30055 33983
rect 30205 33949 30239 33983
rect 3065 33881 3099 33915
rect 6377 33881 6411 33915
rect 7573 33881 7607 33915
rect 10517 33881 10551 33915
rect 12541 33881 12575 33915
rect 16681 33881 16715 33915
rect 17877 33881 17911 33915
rect 22201 33881 22235 33915
rect 26525 33881 26559 33915
rect 27445 33881 27479 33915
rect 2605 33813 2639 33847
rect 3157 33813 3191 33847
rect 5457 33813 5491 33847
rect 6009 33813 6043 33847
rect 14197 33813 14231 33847
rect 21373 33813 21407 33847
rect 24225 33813 24259 33847
rect 25881 33813 25915 33847
rect 25973 33813 26007 33847
rect 26341 33813 26375 33847
rect 27629 33813 27663 33847
rect 27721 33813 27755 33847
rect 27813 33813 27847 33847
rect 1961 33609 1995 33643
rect 3433 33609 3467 33643
rect 7021 33609 7055 33643
rect 8677 33609 8711 33643
rect 8769 33609 8803 33643
rect 9873 33609 9907 33643
rect 10609 33609 10643 33643
rect 11627 33609 11661 33643
rect 12449 33609 12483 33643
rect 13093 33609 13127 33643
rect 14013 33609 14047 33643
rect 23397 33609 23431 33643
rect 24409 33609 24443 33643
rect 25513 33609 25547 33643
rect 2320 33541 2354 33575
rect 9505 33541 9539 33575
rect 10977 33541 11011 33575
rect 11897 33541 11931 33575
rect 12817 33541 12851 33575
rect 14197 33541 14231 33575
rect 17509 33541 17543 33575
rect 24685 33541 24719 33575
rect 26157 33541 26191 33575
rect 26525 33541 26559 33575
rect 28917 33541 28951 33575
rect 29377 33541 29411 33575
rect 3893 33473 3927 33507
rect 5825 33473 5859 33507
rect 6377 33473 6411 33507
rect 8493 33473 8527 33507
rect 8677 33473 8711 33507
rect 8953 33473 8987 33507
rect 9229 33473 9263 33507
rect 9413 33473 9447 33507
rect 9689 33473 9723 33507
rect 10609 33473 10643 33507
rect 10701 33473 10735 33507
rect 11161 33473 11195 33507
rect 11529 33473 11563 33507
rect 11713 33473 11747 33507
rect 11805 33473 11839 33507
rect 12081 33473 12115 33507
rect 12265 33473 12299 33507
rect 12357 33473 12391 33507
rect 12633 33473 12667 33507
rect 12909 33473 12943 33507
rect 13001 33473 13035 33507
rect 13185 33473 13219 33507
rect 13277 33473 13311 33507
rect 13461 33473 13495 33507
rect 14105 33473 14139 33507
rect 14289 33473 14323 33507
rect 14565 33473 14599 33507
rect 14749 33473 14783 33507
rect 15485 33473 15519 33507
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 16313 33473 16347 33507
rect 16405 33473 16439 33507
rect 16865 33473 16899 33507
rect 17233 33473 17267 33507
rect 17693 33473 17727 33507
rect 18245 33473 18279 33507
rect 18889 33473 18923 33507
rect 19073 33473 19107 33507
rect 19625 33473 19659 33507
rect 19892 33473 19926 33507
rect 21281 33473 21315 33507
rect 21446 33473 21480 33507
rect 21557 33473 21591 33507
rect 21649 33473 21683 33507
rect 22284 33473 22318 33507
rect 23673 33473 23707 33507
rect 24041 33473 24075 33507
rect 24593 33473 24627 33507
rect 24777 33473 24811 33507
rect 24961 33473 24995 33507
rect 25053 33473 25087 33507
rect 25329 33473 25363 33507
rect 25789 33473 25823 33507
rect 26065 33473 26099 33507
rect 26249 33473 26283 33507
rect 28181 33473 28215 33507
rect 29653 33473 29687 33507
rect 29837 33473 29871 33507
rect 29929 33473 29963 33507
rect 2053 33405 2087 33439
rect 3985 33405 4019 33439
rect 4077 33405 4111 33439
rect 4905 33405 4939 33439
rect 5733 33405 5767 33439
rect 7389 33405 7423 33439
rect 10885 33405 10919 33439
rect 14841 33405 14875 33439
rect 15577 33405 15611 33439
rect 15761 33405 15795 33439
rect 16681 33405 16715 33439
rect 18521 33405 18555 33439
rect 22017 33405 22051 33439
rect 25145 33405 25179 33439
rect 25881 33405 25915 33439
rect 27537 33405 27571 33439
rect 28089 33405 28123 33439
rect 30021 33405 30055 33439
rect 3525 33337 3559 33371
rect 6193 33337 6227 33371
rect 27997 33337 28031 33371
rect 4537 33269 4571 33303
rect 5549 33269 5583 33303
rect 7941 33269 7975 33303
rect 8401 33269 8435 33303
rect 10517 33269 10551 33303
rect 11345 33269 11379 33303
rect 13369 33269 13403 33303
rect 14381 33269 14415 33303
rect 15117 33269 15151 33303
rect 16773 33269 16807 33303
rect 21005 33269 21039 33303
rect 21097 33269 21131 33303
rect 23581 33269 23615 33303
rect 27169 33269 27203 33303
rect 28365 33269 28399 33303
rect 29469 33269 29503 33303
rect 30665 33269 30699 33303
rect 3249 33065 3283 33099
rect 3525 33065 3559 33099
rect 6009 33065 6043 33099
rect 9137 33065 9171 33099
rect 9413 33065 9447 33099
rect 10425 33065 10459 33099
rect 10701 33065 10735 33099
rect 11621 33065 11655 33099
rect 12633 33065 12667 33099
rect 13829 33065 13863 33099
rect 16221 33065 16255 33099
rect 22293 33065 22327 33099
rect 25513 33065 25547 33099
rect 27905 33065 27939 33099
rect 28549 33065 28583 33099
rect 11253 32997 11287 33031
rect 12357 32997 12391 33031
rect 17693 32997 17727 33031
rect 18245 32997 18279 33031
rect 20821 32997 20855 33031
rect 25697 32997 25731 33031
rect 26249 32997 26283 33031
rect 10057 32929 10091 32963
rect 11897 32929 11931 32963
rect 13277 32929 13311 32963
rect 13461 32929 13495 32963
rect 17509 32929 17543 32963
rect 22385 32929 22419 32963
rect 29837 32929 29871 32963
rect 1409 32861 1443 32895
rect 1869 32861 1903 32895
rect 3433 32861 3467 32895
rect 4629 32861 4663 32895
rect 6377 32861 6411 32895
rect 8217 32861 8251 32895
rect 8953 32861 8987 32895
rect 9046 32861 9080 32895
rect 9781 32861 9815 32895
rect 10701 32861 10735 32895
rect 10885 32861 10919 32895
rect 11437 32861 11471 32895
rect 11713 32861 11747 32895
rect 11989 32861 12023 32895
rect 13553 32861 13587 32895
rect 14105 32861 14139 32895
rect 14841 32861 14875 32895
rect 16405 32861 16439 32895
rect 17969 32861 18003 32895
rect 18429 32861 18463 32895
rect 19717 32861 19751 32895
rect 19809 32861 19843 32895
rect 19901 32861 19935 32895
rect 20085 32861 20119 32895
rect 20269 32861 20303 32895
rect 20913 32861 20947 32895
rect 23305 32861 23339 32895
rect 23581 32861 23615 32895
rect 24501 32861 24535 32895
rect 25145 32861 25179 32895
rect 25421 32861 25455 32895
rect 26065 32861 26099 32895
rect 26341 32861 26375 32895
rect 26893 32861 26927 32895
rect 27077 32861 27111 32895
rect 27445 32861 27479 32895
rect 27537 32861 27571 32895
rect 27721 32861 27755 32895
rect 27813 32861 27847 32895
rect 28181 32861 28215 32895
rect 29101 32861 29135 32895
rect 29193 32861 29227 32895
rect 2136 32793 2170 32827
rect 4874 32793 4908 32827
rect 6644 32793 6678 32827
rect 10241 32793 10275 32827
rect 12449 32793 12483 32827
rect 12649 32793 12683 32827
rect 15108 32793 15142 32827
rect 18061 32793 18095 32827
rect 21180 32793 21214 32827
rect 23029 32793 23063 32827
rect 24133 32793 24167 32827
rect 25881 32793 25915 32827
rect 26617 32793 26651 32827
rect 27905 32793 27939 32827
rect 29377 32793 29411 32827
rect 30082 32793 30116 32827
rect 1593 32725 1627 32759
rect 3985 32725 4019 32759
rect 4537 32725 4571 32759
rect 7757 32725 7791 32759
rect 8769 32725 8803 32759
rect 9873 32725 9907 32759
rect 10441 32725 10475 32759
rect 10609 32725 10643 32759
rect 12817 32725 12851 32759
rect 14749 32725 14783 32759
rect 17049 32725 17083 32759
rect 17877 32725 17911 32759
rect 19073 32725 19107 32759
rect 19441 32725 19475 32759
rect 25053 32725 25087 32759
rect 26985 32725 27019 32759
rect 27261 32725 27295 32759
rect 28089 32725 28123 32759
rect 28825 32725 28859 32759
rect 31217 32725 31251 32759
rect 7941 32521 7975 32555
rect 8309 32521 8343 32555
rect 11345 32521 11379 32555
rect 13645 32521 13679 32555
rect 14105 32521 14139 32555
rect 15209 32521 15243 32555
rect 15577 32521 15611 32555
rect 15669 32521 15703 32555
rect 16497 32521 16531 32555
rect 20545 32521 20579 32555
rect 21005 32521 21039 32555
rect 22477 32521 22511 32555
rect 24777 32521 24811 32555
rect 24869 32521 24903 32555
rect 25697 32521 25731 32555
rect 27169 32521 27203 32555
rect 27721 32521 27755 32555
rect 28825 32521 28859 32555
rect 29653 32521 29687 32555
rect 8769 32453 8803 32487
rect 8985 32453 9019 32487
rect 13277 32453 13311 32487
rect 16129 32453 16163 32487
rect 22836 32453 22870 32487
rect 29285 32453 29319 32487
rect 30840 32453 30874 32487
rect 1593 32385 1627 32419
rect 3709 32385 3743 32419
rect 4629 32385 4663 32419
rect 4896 32385 4930 32419
rect 6644 32385 6678 32419
rect 11805 32385 11839 32419
rect 14013 32385 14047 32419
rect 14289 32385 14323 32419
rect 14381 32385 14415 32419
rect 14473 32385 14507 32419
rect 14591 32385 14625 32419
rect 14933 32385 14967 32419
rect 16313 32385 16347 32419
rect 16681 32385 16715 32419
rect 16865 32385 16899 32419
rect 17969 32385 18003 32419
rect 18236 32385 18270 32419
rect 19625 32385 19659 32419
rect 19993 32385 20027 32419
rect 20821 32385 20855 32419
rect 24041 32385 24075 32419
rect 24225 32385 24259 32419
rect 24593 32385 24627 32419
rect 25237 32385 25271 32419
rect 25513 32385 25547 32419
rect 25789 32385 25823 32419
rect 26065 32385 26099 32419
rect 26249 32385 26283 32419
rect 26341 32385 26375 32419
rect 26617 32385 26651 32419
rect 26801 32385 26835 32419
rect 27166 32385 27200 32419
rect 27629 32385 27663 32419
rect 27905 32385 27939 32419
rect 28181 32385 28215 32419
rect 28365 32385 28399 32419
rect 28641 32385 28675 32419
rect 28917 32385 28951 32419
rect 29101 32385 29135 32419
rect 29929 32385 29963 32419
rect 30021 32385 30055 32419
rect 30113 32385 30147 32419
rect 30297 32385 30331 32419
rect 30573 32385 30607 32419
rect 32137 32385 32171 32419
rect 32321 32385 32355 32419
rect 1869 32317 1903 32351
rect 2973 32317 3007 32351
rect 3985 32317 4019 32351
rect 6377 32317 6411 32351
rect 8401 32317 8435 32351
rect 8585 32317 8619 32351
rect 9229 32317 9263 32351
rect 9505 32317 9539 32351
rect 12541 32317 12575 32351
rect 14749 32317 14783 32351
rect 15853 32317 15887 32351
rect 17049 32317 17083 32351
rect 17233 32317 17267 32351
rect 19441 32317 19475 32351
rect 20637 32317 20671 32351
rect 22569 32317 22603 32351
rect 24317 32317 24351 32351
rect 24409 32317 24443 32351
rect 25053 32317 25087 32351
rect 25145 32317 25179 32351
rect 25329 32317 25363 32351
rect 27537 32317 27571 32351
rect 28549 32317 28583 32351
rect 6009 32249 6043 32283
rect 7757 32249 7791 32283
rect 9137 32249 9171 32283
rect 10977 32249 11011 32283
rect 15025 32249 15059 32283
rect 26525 32249 26559 32283
rect 26617 32249 26651 32283
rect 27997 32249 28031 32283
rect 28089 32249 28123 32283
rect 3525 32181 3559 32215
rect 8913 32181 8947 32215
rect 10333 32181 10367 32215
rect 12081 32181 12115 32215
rect 12909 32181 12943 32215
rect 17877 32181 17911 32215
rect 19349 32181 19383 32215
rect 19809 32181 19843 32215
rect 21281 32181 21315 32215
rect 22017 32181 22051 32215
rect 23949 32181 23983 32215
rect 25513 32181 25547 32215
rect 26341 32181 26375 32215
rect 26985 32181 27019 32215
rect 28641 32181 28675 32215
rect 31953 32181 31987 32215
rect 32137 32181 32171 32215
rect 32689 32181 32723 32215
rect 3801 31977 3835 32011
rect 4813 31977 4847 32011
rect 5917 31977 5951 32011
rect 7389 31977 7423 32011
rect 10333 31977 10367 32011
rect 15393 31977 15427 32011
rect 17877 31977 17911 32011
rect 18889 31977 18923 32011
rect 21557 31977 21591 32011
rect 25513 31977 25547 32011
rect 25697 31977 25731 32011
rect 31401 31977 31435 32011
rect 33057 31977 33091 32011
rect 6377 31909 6411 31943
rect 13093 31909 13127 31943
rect 19533 31909 19567 31943
rect 21005 31909 21039 31943
rect 23489 31909 23523 31943
rect 25145 31909 25179 31943
rect 28365 31909 28399 31943
rect 1685 31841 1719 31875
rect 4353 31841 4387 31875
rect 5273 31841 5307 31875
rect 5365 31841 5399 31875
rect 12817 31841 12851 31875
rect 14105 31841 14139 31875
rect 15669 31841 15703 31875
rect 18153 31841 18187 31875
rect 18245 31841 18279 31875
rect 19625 31841 19659 31875
rect 22109 31841 22143 31875
rect 24593 31841 24627 31875
rect 26525 31841 26559 31875
rect 26893 31841 26927 31875
rect 26985 31841 27019 31875
rect 30849 31841 30883 31875
rect 32229 31841 32263 31875
rect 32689 31841 32723 31875
rect 1952 31773 1986 31807
rect 6101 31773 6135 31807
rect 6377 31773 6411 31807
rect 6561 31773 6595 31807
rect 6837 31773 6871 31807
rect 8033 31773 8067 31807
rect 8125 31773 8159 31807
rect 8953 31773 8987 31807
rect 10701 31773 10735 31807
rect 11529 31773 11563 31807
rect 11897 31773 11931 31807
rect 12081 31773 12115 31807
rect 14381 31773 14415 31807
rect 15207 31773 15241 31807
rect 16405 31773 16439 31807
rect 18061 31773 18095 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 18705 31773 18739 31807
rect 19349 31773 19383 31807
rect 19892 31773 19926 31807
rect 21097 31773 21131 31807
rect 21189 31773 21223 31807
rect 21465 31773 21499 31807
rect 21649 31773 21683 31807
rect 22376 31773 22410 31807
rect 23581 31773 23615 31807
rect 24409 31773 24443 31807
rect 25145 31773 25179 31807
rect 25329 31773 25363 31807
rect 25421 31773 25455 31807
rect 26065 31773 26099 31807
rect 26341 31773 26375 31807
rect 26433 31773 26467 31807
rect 26709 31773 26743 31807
rect 26801 31773 26835 31807
rect 27169 31773 27203 31807
rect 28181 31773 28215 31807
rect 28825 31773 28859 31807
rect 28917 31773 28951 31807
rect 29745 31773 29779 31807
rect 30113 31773 30147 31807
rect 30297 31773 30331 31807
rect 30385 31773 30419 31807
rect 30481 31773 30515 31807
rect 31493 31773 31527 31807
rect 32413 31773 32447 31807
rect 32873 31773 32907 31807
rect 3433 31705 3467 31739
rect 4169 31705 4203 31739
rect 9198 31705 9232 31739
rect 15025 31705 15059 31739
rect 16672 31705 16706 31739
rect 21373 31705 21407 31739
rect 25979 31705 26013 31739
rect 27997 31705 28031 31739
rect 3065 31637 3099 31671
rect 3525 31637 3559 31671
rect 4261 31637 4295 31671
rect 5181 31637 5215 31671
rect 6285 31637 6319 31671
rect 8309 31637 8343 31671
rect 8769 31637 8803 31671
rect 11253 31637 11287 31671
rect 12265 31637 12299 31671
rect 13553 31637 13587 31671
rect 13921 31637 13955 31671
rect 16313 31637 16347 31671
rect 17785 31637 17819 31671
rect 21097 31637 21131 31671
rect 21925 31637 21959 31671
rect 24225 31637 24259 31671
rect 26157 31637 26191 31671
rect 28825 31637 28859 31671
rect 30665 31637 30699 31671
rect 32137 31637 32171 31671
rect 32597 31637 32631 31671
rect 3709 31433 3743 31467
rect 6837 31433 6871 31467
rect 8493 31433 8527 31467
rect 17049 31433 17083 31467
rect 17877 31433 17911 31467
rect 18429 31433 18463 31467
rect 19717 31433 19751 31467
rect 23673 31433 23707 31467
rect 24409 31433 24443 31467
rect 24501 31433 24535 31467
rect 26709 31433 26743 31467
rect 27629 31433 27663 31467
rect 29469 31433 29503 31467
rect 6193 31365 6227 31399
rect 6561 31365 6595 31399
rect 7389 31365 7423 31399
rect 8125 31365 8159 31399
rect 9045 31365 9079 31399
rect 18705 31365 18739 31399
rect 18797 31365 18831 31399
rect 18935 31365 18969 31399
rect 22017 31365 22051 31399
rect 22293 31365 22327 31399
rect 24777 31365 24811 31399
rect 24869 31365 24903 31399
rect 25421 31365 25455 31399
rect 1961 31297 1995 31331
rect 2228 31297 2262 31331
rect 4077 31297 4111 31331
rect 4905 31297 4939 31331
rect 4997 31297 5031 31331
rect 5089 31297 5123 31331
rect 5285 31297 5319 31331
rect 6377 31297 6411 31331
rect 7113 31297 7147 31331
rect 7665 31297 7699 31331
rect 7849 31297 7883 31331
rect 7941 31297 7975 31331
rect 8217 31297 8251 31331
rect 8309 31297 8343 31331
rect 8861 31297 8895 31331
rect 8953 31297 8987 31331
rect 9597 31297 9631 31331
rect 11529 31297 11563 31331
rect 11785 31297 11819 31331
rect 13185 31297 13219 31331
rect 13452 31297 13486 31331
rect 15025 31297 15059 31331
rect 15281 31297 15315 31331
rect 16773 31297 16807 31331
rect 16865 31297 16899 31331
rect 17693 31297 17727 31331
rect 17969 31297 18003 31331
rect 18153 31297 18187 31331
rect 18613 31297 18647 31331
rect 19165 31297 19199 31331
rect 19349 31297 19383 31331
rect 19901 31297 19935 31331
rect 20085 31297 20119 31331
rect 20177 31297 20211 31331
rect 20361 31297 20395 31331
rect 20545 31297 20579 31331
rect 21833 31297 21867 31331
rect 22523 31297 22557 31331
rect 22642 31297 22676 31331
rect 22753 31297 22787 31331
rect 22937 31297 22971 31331
rect 24685 31297 24719 31331
rect 25053 31297 25087 31331
rect 25145 31297 25179 31331
rect 25237 31297 25271 31331
rect 25697 31297 25731 31331
rect 25881 31297 25915 31331
rect 26341 31297 26375 31331
rect 26433 31297 26467 31331
rect 26617 31297 26651 31331
rect 26801 31297 26835 31331
rect 27997 31297 28031 31331
rect 28089 31297 28123 31331
rect 28457 31297 28491 31331
rect 28641 31297 28675 31331
rect 29101 31297 29135 31331
rect 29377 31297 29411 31331
rect 29561 31297 29595 31331
rect 29909 31297 29943 31331
rect 31585 31297 31619 31331
rect 4169 31229 4203 31263
rect 4353 31229 4387 31263
rect 5549 31229 5583 31263
rect 6745 31229 6779 31263
rect 7021 31229 7055 31263
rect 7481 31229 7515 31263
rect 7757 31229 7791 31263
rect 9321 31229 9355 31263
rect 9873 31229 9907 31263
rect 17601 31229 17635 31263
rect 19073 31229 19107 31263
rect 21005 31229 21039 31263
rect 23029 31229 23063 31263
rect 26157 31229 26191 31263
rect 26249 31229 26283 31263
rect 28181 31229 28215 31263
rect 29653 31229 29687 31263
rect 17509 31161 17543 31195
rect 19441 31161 19475 31195
rect 22201 31161 22235 31195
rect 25697 31161 25731 31195
rect 25973 31161 26007 31195
rect 28549 31161 28583 31195
rect 1869 31093 1903 31127
rect 3341 31093 3375 31127
rect 4629 31093 4663 31127
rect 8585 31093 8619 31127
rect 9229 31093 9263 31127
rect 10977 31093 11011 31127
rect 12909 31093 12943 31127
rect 14565 31093 14599 31127
rect 16405 31093 16439 31127
rect 17233 31093 17267 31127
rect 18337 31093 18371 31127
rect 20729 31093 20763 31127
rect 21649 31093 21683 31127
rect 25513 31093 25547 31127
rect 31033 31093 31067 31127
rect 31401 31093 31435 31127
rect 31769 31093 31803 31127
rect 2881 30889 2915 30923
rect 3985 30889 4019 30923
rect 4537 30889 4571 30923
rect 5733 30889 5767 30923
rect 6653 30889 6687 30923
rect 7113 30889 7147 30923
rect 8769 30889 8803 30923
rect 9689 30889 9723 30923
rect 10977 30889 11011 30923
rect 11161 30889 11195 30923
rect 14105 30889 14139 30923
rect 15209 30889 15243 30923
rect 16957 30889 16991 30923
rect 17509 30889 17543 30923
rect 18705 30889 18739 30923
rect 23305 30889 23339 30923
rect 27353 30889 27387 30923
rect 28181 30889 28215 30923
rect 28457 30889 28491 30923
rect 29561 30889 29595 30923
rect 30665 30889 30699 30923
rect 4445 30821 4479 30855
rect 5181 30821 5215 30855
rect 5549 30821 5583 30855
rect 7389 30821 7423 30855
rect 7665 30821 7699 30855
rect 8401 30821 8435 30855
rect 13921 30821 13955 30855
rect 15301 30821 15335 30855
rect 17049 30821 17083 30855
rect 17877 30821 17911 30855
rect 18889 30821 18923 30855
rect 26341 30821 26375 30855
rect 1869 30753 1903 30787
rect 3525 30753 3559 30787
rect 6837 30753 6871 30787
rect 9597 30753 9631 30787
rect 10333 30753 10367 30787
rect 11621 30753 11655 30787
rect 11805 30753 11839 30787
rect 12817 30753 12851 30787
rect 14749 30753 14783 30787
rect 15761 30753 15795 30787
rect 15945 30753 15979 30787
rect 18061 30753 18095 30787
rect 20913 30753 20947 30787
rect 23213 30753 23247 30787
rect 24501 30753 24535 30787
rect 24685 30753 24719 30787
rect 24777 30753 24811 30787
rect 24961 30753 24995 30787
rect 27537 30753 27571 30787
rect 28181 30753 28215 30787
rect 1593 30685 1627 30719
rect 3801 30685 3835 30719
rect 4721 30685 4755 30719
rect 4813 30685 4847 30719
rect 4997 30685 5031 30719
rect 5089 30685 5123 30719
rect 5365 30685 5399 30719
rect 5641 30685 5675 30719
rect 5733 30685 5767 30719
rect 5917 30685 5951 30719
rect 6745 30685 6779 30719
rect 6929 30685 6963 30719
rect 7113 30685 7147 30719
rect 7297 30685 7331 30719
rect 7573 30685 7607 30719
rect 7757 30685 7791 30719
rect 7849 30685 7883 30719
rect 9229 30685 9263 30719
rect 9413 30685 9447 30719
rect 10057 30685 10091 30719
rect 11529 30685 11563 30719
rect 12173 30685 12207 30719
rect 12449 30685 12483 30719
rect 12725 30685 12759 30719
rect 13461 30685 13495 30719
rect 16681 30685 16715 30719
rect 16773 30685 16807 30719
rect 17325 30685 17359 30719
rect 17785 30685 17819 30719
rect 17969 30685 18003 30719
rect 18245 30685 18279 30719
rect 18337 30685 18371 30719
rect 19257 30685 19291 30719
rect 19809 30685 19843 30719
rect 19993 30685 20027 30719
rect 20177 30685 20211 30719
rect 20453 30685 20487 30719
rect 22385 30685 22419 30719
rect 23121 30685 23155 30719
rect 23857 30685 23891 30719
rect 24869 30685 24903 30719
rect 25145 30685 25179 30719
rect 25329 30685 25363 30719
rect 25421 30685 25455 30719
rect 25605 30685 25639 30719
rect 27629 30685 27663 30719
rect 28089 30685 28123 30719
rect 28917 30685 28951 30719
rect 29745 30685 29779 30719
rect 29837 30685 29871 30719
rect 30113 30685 30147 30719
rect 30481 30685 30515 30719
rect 30849 30685 30883 30719
rect 31116 30685 31150 30719
rect 32413 30685 32447 30719
rect 3341 30617 3375 30651
rect 10149 30617 10183 30651
rect 11989 30617 12023 30651
rect 12357 30617 12391 30651
rect 14565 30617 14599 30651
rect 16313 30617 16347 30651
rect 17049 30617 17083 30651
rect 18705 30617 18739 30651
rect 19533 30617 19567 30651
rect 21180 30617 21214 30651
rect 23029 30617 23063 30651
rect 25513 30617 25547 30651
rect 25973 30617 26007 30651
rect 26157 30617 26191 30651
rect 27905 30617 27939 30651
rect 27997 30617 28031 30651
rect 28641 30617 28675 30651
rect 29193 30617 29227 30651
rect 29561 30617 29595 30651
rect 30297 30617 30331 30651
rect 30389 30617 30423 30651
rect 3249 30549 3283 30583
rect 6285 30549 6319 30583
rect 13093 30549 13127 30583
rect 14473 30549 14507 30583
rect 15669 30549 15703 30583
rect 17233 30549 17267 30583
rect 19901 30549 19935 30583
rect 20361 30549 20395 30583
rect 20545 30549 20579 30583
rect 22293 30549 22327 30583
rect 23489 30549 23523 30583
rect 25237 30549 25271 30583
rect 28825 30549 28859 30583
rect 29009 30549 29043 30583
rect 32229 30549 32263 30583
rect 32965 30549 32999 30583
rect 2053 30345 2087 30379
rect 2789 30345 2823 30379
rect 5457 30345 5491 30379
rect 6929 30345 6963 30379
rect 7849 30345 7883 30379
rect 8217 30345 8251 30379
rect 10241 30345 10275 30379
rect 10885 30345 10919 30379
rect 12265 30345 12299 30379
rect 13001 30345 13035 30379
rect 14289 30345 14323 30379
rect 15117 30345 15151 30379
rect 16497 30345 16531 30379
rect 21189 30345 21223 30379
rect 21833 30345 21867 30379
rect 29561 30345 29595 30379
rect 33517 30345 33551 30379
rect 2237 30277 2271 30311
rect 3801 30277 3835 30311
rect 3985 30277 4019 30311
rect 4077 30277 4111 30311
rect 4261 30277 4295 30311
rect 4353 30277 4387 30311
rect 4629 30277 4663 30311
rect 5825 30277 5859 30311
rect 7113 30277 7147 30311
rect 16957 30277 16991 30311
rect 21465 30277 21499 30311
rect 21649 30277 21683 30311
rect 23213 30277 23247 30311
rect 24225 30277 24259 30311
rect 24501 30277 24535 30311
rect 26985 30277 27019 30311
rect 30205 30277 30239 30311
rect 31677 30277 31711 30311
rect 2145 30209 2179 30243
rect 2329 30209 2363 30243
rect 2513 30209 2547 30243
rect 2605 30209 2639 30243
rect 3065 30209 3099 30243
rect 3341 30209 3375 30243
rect 3617 30209 3651 30243
rect 3709 30209 3743 30243
rect 4450 30209 4484 30243
rect 4813 30209 4847 30243
rect 5089 30209 5123 30243
rect 5549 30209 5583 30243
rect 6653 30209 6687 30243
rect 6745 30209 6779 30243
rect 7021 30209 7055 30243
rect 7205 30209 7239 30243
rect 7481 30209 7515 30243
rect 8401 30209 8435 30243
rect 8493 30209 8527 30243
rect 8677 30209 8711 30243
rect 8769 30209 8803 30243
rect 9045 30209 9079 30243
rect 10517 30209 10551 30243
rect 11345 30209 11379 30243
rect 11529 30209 11563 30243
rect 11622 30209 11656 30243
rect 12173 30209 12207 30243
rect 12357 30209 12391 30243
rect 12633 30209 12667 30243
rect 12726 30209 12760 30243
rect 13553 30209 13587 30243
rect 13737 30209 13771 30243
rect 14105 30209 14139 30243
rect 15025 30209 15059 30243
rect 15485 30209 15519 30243
rect 15945 30209 15979 30243
rect 16129 30209 16163 30243
rect 16681 30209 16715 30243
rect 16865 30209 16899 30243
rect 17049 30209 17083 30243
rect 17325 30209 17359 30243
rect 17601 30209 17635 30243
rect 17877 30209 17911 30243
rect 18061 30209 18095 30243
rect 19073 30209 19107 30243
rect 19349 30209 19383 30243
rect 19533 30209 19567 30243
rect 20076 30209 20110 30243
rect 21281 30209 21315 30243
rect 22109 30209 22143 30243
rect 22201 30209 22235 30243
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 22937 30209 22971 30243
rect 23121 30209 23155 30243
rect 23305 30209 23339 30243
rect 23581 30209 23615 30243
rect 23949 30209 23983 30243
rect 24041 30209 24075 30243
rect 24685 30209 24719 30243
rect 25329 30209 25363 30243
rect 25513 30209 25547 30243
rect 25605 30209 25639 30243
rect 25789 30209 25823 30243
rect 26065 30209 26099 30243
rect 26341 30209 26375 30243
rect 26525 30209 26559 30243
rect 26709 30209 26743 30243
rect 27353 30209 27387 30243
rect 27997 30209 28031 30243
rect 28457 30209 28491 30243
rect 28641 30209 28675 30243
rect 29009 30209 29043 30243
rect 29101 30209 29135 30243
rect 29193 30209 29227 30243
rect 29469 30209 29503 30243
rect 29653 30209 29687 30243
rect 29745 30209 29779 30243
rect 30021 30209 30055 30243
rect 30297 30209 30331 30243
rect 30389 30209 30423 30243
rect 30757 30209 30791 30243
rect 31401 30209 31435 30243
rect 31585 30209 31619 30243
rect 31769 30209 31803 30243
rect 32393 30209 32427 30243
rect 3249 30141 3283 30175
rect 4353 30141 4387 30175
rect 5181 30141 5215 30175
rect 7573 30141 7607 30175
rect 9137 30141 9171 30175
rect 9413 30141 9447 30175
rect 10609 30141 10643 30175
rect 11897 30141 11931 30175
rect 13921 30141 13955 30175
rect 14473 30141 14507 30175
rect 15577 30141 15611 30175
rect 15761 30141 15795 30175
rect 16037 30141 16071 30175
rect 17693 30141 17727 30175
rect 18337 30141 18371 30175
rect 19809 30141 19843 30175
rect 23857 30141 23891 30175
rect 24225 30141 24259 30175
rect 24961 30141 24995 30175
rect 26157 30141 26191 30175
rect 28273 30141 28307 30175
rect 29285 30141 29319 30175
rect 32137 30141 32171 30175
rect 3433 30073 3467 30107
rect 5641 30073 5675 30107
rect 13277 30073 13311 30107
rect 19441 30073 19475 30107
rect 25421 30073 25455 30107
rect 26249 30073 26283 30107
rect 27261 30073 27295 30107
rect 28825 30073 28859 30107
rect 2881 30005 2915 30039
rect 4997 30005 5031 30039
rect 5273 30005 5307 30039
rect 5733 30005 5767 30039
rect 7665 30005 7699 30039
rect 13553 30005 13587 30039
rect 17233 30005 17267 30039
rect 18889 30005 18923 30039
rect 19257 30005 19291 30039
rect 22753 30005 22787 30039
rect 23489 30005 23523 30039
rect 23673 30005 23707 30039
rect 23765 30005 23799 30039
rect 24869 30005 24903 30039
rect 25145 30005 25179 30039
rect 25881 30005 25915 30039
rect 26617 30005 26651 30039
rect 26985 30005 27019 30039
rect 27169 30005 27203 30039
rect 27813 30005 27847 30039
rect 28181 30005 28215 30039
rect 28549 30005 28583 30039
rect 29837 30005 29871 30039
rect 30573 30005 30607 30039
rect 31309 30005 31343 30039
rect 31953 30005 31987 30039
rect 3157 29801 3191 29835
rect 3525 29801 3559 29835
rect 4445 29801 4479 29835
rect 4721 29801 4755 29835
rect 6653 29801 6687 29835
rect 7665 29801 7699 29835
rect 8217 29801 8251 29835
rect 8585 29801 8619 29835
rect 9321 29801 9355 29835
rect 9965 29801 9999 29835
rect 11713 29801 11747 29835
rect 12449 29801 12483 29835
rect 20637 29801 20671 29835
rect 22109 29801 22143 29835
rect 24409 29801 24443 29835
rect 24777 29801 24811 29835
rect 26617 29801 26651 29835
rect 27721 29801 27755 29835
rect 27813 29801 27847 29835
rect 30941 29801 30975 29835
rect 32781 29801 32815 29835
rect 4261 29733 4295 29767
rect 12633 29733 12667 29767
rect 14565 29733 14599 29767
rect 16037 29733 16071 29767
rect 25053 29733 25087 29767
rect 25513 29733 25547 29767
rect 27261 29733 27295 29767
rect 1869 29665 1903 29699
rect 3065 29665 3099 29699
rect 3249 29635 3283 29669
rect 3617 29665 3651 29699
rect 3893 29665 3927 29699
rect 5365 29665 5399 29699
rect 5825 29665 5859 29699
rect 7297 29665 7331 29699
rect 8033 29665 8067 29699
rect 12173 29665 12207 29699
rect 13369 29665 13403 29699
rect 14749 29665 14783 29699
rect 16589 29665 16623 29699
rect 17693 29665 17727 29699
rect 20729 29665 20763 29699
rect 21465 29665 21499 29699
rect 23121 29665 23155 29699
rect 30573 29665 30607 29699
rect 31769 29665 31803 29699
rect 1593 29597 1627 29631
rect 2973 29597 3007 29631
rect 3341 29597 3375 29631
rect 3433 29597 3467 29631
rect 4077 29597 4111 29631
rect 4353 29597 4387 29631
rect 4537 29597 4571 29631
rect 4905 29597 4939 29631
rect 4997 29597 5031 29631
rect 5181 29597 5215 29631
rect 5273 29597 5307 29631
rect 5549 29597 5583 29631
rect 5733 29597 5767 29631
rect 6837 29597 6871 29631
rect 6929 29597 6963 29631
rect 7113 29597 7147 29631
rect 7205 29597 7239 29631
rect 7481 29597 7515 29631
rect 7757 29597 7791 29631
rect 7941 29597 7975 29631
rect 8125 29597 8159 29631
rect 8401 29597 8435 29631
rect 8677 29597 8711 29631
rect 9321 29597 9355 29631
rect 9505 29597 9539 29631
rect 10149 29597 10183 29631
rect 10425 29597 10459 29631
rect 11621 29597 11655 29631
rect 11805 29597 11839 29631
rect 11897 29597 11931 29631
rect 11989 29597 12023 29631
rect 13093 29597 13127 29631
rect 13185 29597 13219 29631
rect 13553 29597 13587 29631
rect 13737 29597 13771 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 14933 29597 14967 29631
rect 15393 29597 15427 29631
rect 15541 29597 15575 29631
rect 15858 29597 15892 29631
rect 19257 29597 19291 29631
rect 21005 29597 21039 29631
rect 21097 29597 21131 29631
rect 21189 29597 21223 29631
rect 21373 29597 21407 29631
rect 22201 29597 22235 29631
rect 22385 29597 22419 29631
rect 22753 29597 22787 29631
rect 22937 29597 22971 29631
rect 23029 29597 23063 29631
rect 23213 29597 23247 29631
rect 23397 29597 23431 29631
rect 23765 29597 23799 29631
rect 24593 29597 24627 29631
rect 24869 29597 24903 29631
rect 25053 29597 25087 29631
rect 25237 29597 25271 29631
rect 26249 29597 26283 29631
rect 27353 29597 27387 29631
rect 27813 29597 27847 29631
rect 27997 29597 28031 29631
rect 29193 29597 29227 29631
rect 29377 29597 29411 29631
rect 30297 29597 30331 29631
rect 30481 29597 30515 29631
rect 30757 29597 30791 29631
rect 31033 29597 31067 29631
rect 31401 29597 31435 29631
rect 32413 29597 32447 29631
rect 32965 29597 32999 29631
rect 35265 29597 35299 29631
rect 35449 29597 35483 29631
rect 12173 29529 12207 29563
rect 12311 29529 12345 29563
rect 12481 29529 12515 29563
rect 13645 29529 13679 29563
rect 15117 29529 15151 29563
rect 15669 29529 15703 29563
rect 15761 29529 15795 29563
rect 17509 29529 17543 29563
rect 17960 29529 17994 29563
rect 19524 29529 19558 29563
rect 23581 29529 23615 29563
rect 23673 29529 23707 29563
rect 26433 29529 26467 29563
rect 26893 29529 26927 29563
rect 27077 29529 27111 29563
rect 27537 29529 27571 29563
rect 31217 29529 31251 29563
rect 31309 29529 31343 29563
rect 33701 29529 33735 29563
rect 36277 29529 36311 29563
rect 10333 29461 10367 29495
rect 12725 29461 12759 29495
rect 17141 29461 17175 29495
rect 19073 29461 19107 29495
rect 22569 29461 22603 29495
rect 23949 29461 23983 29495
rect 29285 29461 29319 29495
rect 30389 29461 30423 29495
rect 31585 29461 31619 29495
rect 3449 29257 3483 29291
rect 3617 29257 3651 29291
rect 3801 29257 3835 29291
rect 4819 29257 4853 29291
rect 5181 29257 5215 29291
rect 7957 29257 7991 29291
rect 8125 29257 8159 29291
rect 9051 29257 9085 29291
rect 10701 29257 10735 29291
rect 12633 29257 12667 29291
rect 12817 29257 12851 29291
rect 14749 29257 14783 29291
rect 17877 29257 17911 29291
rect 18337 29257 18371 29291
rect 18521 29257 18555 29291
rect 19441 29257 19475 29291
rect 20821 29257 20855 29291
rect 25697 29257 25731 29291
rect 26985 29257 27019 29291
rect 30481 29257 30515 29291
rect 33609 29257 33643 29291
rect 34529 29257 34563 29291
rect 1869 29189 1903 29223
rect 2605 29189 2639 29223
rect 3249 29189 3283 29223
rect 4905 29189 4939 29223
rect 7757 29189 7791 29223
rect 8953 29189 8987 29223
rect 9689 29189 9723 29223
rect 10057 29189 10091 29223
rect 10425 29189 10459 29223
rect 14473 29189 14507 29223
rect 17049 29189 17083 29223
rect 24869 29189 24903 29223
rect 27997 29189 28031 29223
rect 29285 29189 29319 29223
rect 30849 29189 30883 29223
rect 30941 29189 30975 29223
rect 31953 29189 31987 29223
rect 32965 29189 32999 29223
rect 2053 29121 2087 29155
rect 2145 29121 2179 29155
rect 2421 29121 2455 29155
rect 2697 29121 2731 29155
rect 2881 29121 2915 29155
rect 3065 29121 3099 29155
rect 3709 29121 3743 29155
rect 3893 29121 3927 29155
rect 4537 29121 4571 29155
rect 4721 29121 4755 29155
rect 4997 29121 5031 29155
rect 5089 29121 5123 29155
rect 5285 29121 5319 29155
rect 6837 29121 6871 29155
rect 7021 29121 7055 29155
rect 7113 29121 7147 29155
rect 7389 29121 7423 29155
rect 7573 29121 7607 29155
rect 7665 29121 7699 29155
rect 9137 29121 9171 29155
rect 9229 29121 9263 29155
rect 9524 29121 9558 29155
rect 9781 29121 9815 29155
rect 10241 29121 10275 29155
rect 10527 29143 10561 29177
rect 10885 29121 10919 29155
rect 11069 29121 11103 29155
rect 11161 29121 11195 29155
rect 12265 29121 12299 29155
rect 12814 29121 12848 29155
rect 13645 29121 13679 29155
rect 14197 29121 14231 29155
rect 14381 29121 14415 29155
rect 14657 29121 14691 29155
rect 15485 29121 15519 29155
rect 16129 29121 16163 29155
rect 18797 29121 18831 29155
rect 18889 29121 18923 29155
rect 18981 29121 19015 29155
rect 19165 29121 19199 29155
rect 19717 29121 19751 29155
rect 19809 29121 19843 29155
rect 19901 29121 19935 29155
rect 20085 29121 20119 29155
rect 21097 29121 21131 29155
rect 21189 29121 21223 29155
rect 21373 29121 21407 29155
rect 21475 29121 21509 29155
rect 21925 29121 21959 29155
rect 23029 29121 23063 29155
rect 23213 29121 23247 29155
rect 23581 29121 23615 29155
rect 23673 29121 23707 29155
rect 23857 29121 23891 29155
rect 23949 29121 23983 29155
rect 24409 29121 24443 29155
rect 24501 29121 24535 29155
rect 24593 29121 24627 29155
rect 24685 29121 24719 29155
rect 25053 29121 25087 29155
rect 25329 29121 25363 29155
rect 25422 29121 25456 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 27629 29121 27663 29155
rect 27721 29121 27755 29155
rect 28181 29121 28215 29155
rect 28825 29121 28859 29155
rect 28917 29121 28951 29155
rect 29009 29121 29043 29155
rect 29193 29121 29227 29155
rect 29377 29121 29411 29155
rect 29469 29121 29503 29155
rect 29653 29121 29687 29155
rect 29745 29121 29779 29155
rect 29929 29121 29963 29155
rect 30297 29121 30331 29155
rect 30665 29121 30699 29155
rect 31033 29121 31067 29155
rect 31309 29121 31343 29155
rect 32137 29121 32171 29155
rect 33517 29121 33551 29155
rect 9321 29053 9355 29087
rect 12541 29053 12575 29087
rect 13277 29053 13311 29087
rect 13921 29053 13955 29087
rect 15669 29053 15703 29087
rect 15853 29053 15887 29087
rect 17325 29053 17359 29087
rect 20177 29053 20211 29087
rect 22937 29053 22971 29087
rect 24225 29053 24259 29087
rect 27261 29053 27295 29087
rect 27445 29053 27479 29087
rect 28733 29053 28767 29087
rect 30113 29053 30147 29087
rect 1685 28985 1719 29019
rect 1869 28985 1903 29019
rect 2881 28985 2915 29019
rect 6837 28985 6871 29019
rect 13185 28985 13219 29019
rect 13829 28985 13863 29019
rect 25237 28985 25271 29019
rect 27813 28985 27847 29019
rect 28365 28985 28399 29019
rect 28549 28985 28583 29019
rect 29745 28985 29779 29019
rect 31217 28985 31251 29019
rect 32781 28985 32815 29019
rect 34161 28985 34195 29019
rect 2237 28917 2271 28951
rect 3433 28917 3467 28951
rect 4261 28917 4295 28951
rect 7205 28917 7239 28951
rect 7941 28917 7975 28951
rect 12357 28917 12391 28951
rect 12449 28917 12483 28951
rect 13461 28917 13495 28951
rect 20913 28917 20947 28951
rect 23029 28917 23063 28951
rect 23397 28917 23431 28951
rect 25973 28917 26007 28951
rect 29469 28917 29503 28951
rect 33057 28917 33091 28951
rect 2881 28713 2915 28747
rect 3985 28713 4019 28747
rect 4997 28713 5031 28747
rect 6193 28713 6227 28747
rect 7113 28713 7147 28747
rect 7849 28713 7883 28747
rect 9781 28713 9815 28747
rect 9965 28713 9999 28747
rect 11069 28713 11103 28747
rect 11345 28713 11379 28747
rect 12817 28713 12851 28747
rect 13369 28713 13403 28747
rect 14381 28713 14415 28747
rect 17417 28713 17451 28747
rect 18153 28713 18187 28747
rect 19717 28713 19751 28747
rect 20269 28713 20303 28747
rect 23213 28713 23247 28747
rect 23949 28713 23983 28747
rect 26433 28713 26467 28747
rect 27077 28713 27111 28747
rect 27261 28713 27295 28747
rect 33425 28713 33459 28747
rect 11253 28645 11287 28679
rect 14749 28645 14783 28679
rect 15117 28645 15151 28679
rect 19625 28645 19659 28679
rect 19809 28645 19843 28679
rect 28365 28645 28399 28679
rect 29837 28645 29871 28679
rect 42165 28645 42199 28679
rect 1869 28577 1903 28611
rect 8309 28577 8343 28611
rect 8493 28577 8527 28611
rect 11989 28577 12023 28611
rect 12725 28577 12759 28611
rect 13461 28577 13495 28611
rect 18889 28577 18923 28611
rect 20637 28577 20671 28611
rect 24409 28577 24443 28611
rect 26893 28577 26927 28611
rect 29561 28577 29595 28611
rect 30021 28577 30055 28611
rect 32045 28577 32079 28611
rect 42901 28577 42935 28611
rect 43269 28577 43303 28611
rect 1593 28509 1627 28543
rect 3065 28509 3099 28543
rect 3341 28509 3375 28543
rect 5457 28509 5491 28543
rect 5549 28509 5583 28543
rect 5917 28509 5951 28543
rect 7113 28509 7147 28543
rect 7297 28509 7331 28543
rect 8217 28509 8251 28543
rect 12998 28509 13032 28543
rect 13737 28509 13771 28543
rect 16037 28509 16071 28543
rect 17601 28509 17635 28543
rect 17785 28509 17819 28543
rect 17969 28509 18003 28543
rect 18337 28509 18371 28543
rect 19533 28509 19567 28543
rect 19993 28509 20027 28543
rect 20085 28509 20119 28543
rect 20177 28509 20211 28543
rect 21281 28509 21315 28543
rect 23397 28509 23431 28543
rect 25973 28509 26007 28543
rect 26157 28509 26191 28543
rect 27077 28509 27111 28543
rect 27353 28509 27387 28543
rect 27537 28509 27571 28543
rect 27629 28509 27663 28543
rect 27813 28509 27847 28543
rect 28089 28509 28123 28543
rect 28365 28509 28399 28543
rect 28733 28509 28767 28543
rect 30481 28509 30515 28543
rect 30849 28509 30883 28543
rect 31125 28509 31159 28543
rect 31401 28509 31435 28543
rect 33517 28509 33551 28543
rect 33701 28509 33735 28543
rect 42073 28509 42107 28543
rect 42349 28509 42383 28543
rect 42625 28509 42659 28543
rect 43085 28509 43119 28543
rect 43177 28509 43211 28543
rect 5043 28475 5077 28509
rect 9827 28475 9861 28509
rect 3801 28441 3835 28475
rect 4445 28441 4479 28475
rect 4813 28441 4847 28475
rect 5273 28441 5307 28475
rect 9597 28441 9631 28475
rect 10885 28441 10919 28475
rect 13553 28441 13587 28475
rect 15485 28441 15519 28475
rect 16304 28441 16338 28475
rect 17877 28441 17911 28475
rect 21526 28441 21560 28475
rect 26249 28441 26283 28475
rect 26801 28441 26835 28475
rect 30665 28441 30699 28475
rect 30757 28441 30791 28475
rect 32312 28441 32346 28475
rect 3249 28373 3283 28407
rect 4001 28373 4035 28407
rect 4169 28373 4203 28407
rect 5181 28373 5215 28407
rect 5371 28373 5405 28407
rect 11085 28373 11119 28407
rect 11713 28373 11747 28407
rect 11805 28373 11839 28407
rect 13001 28373 13035 28407
rect 13921 28373 13955 28407
rect 15945 28373 15979 28407
rect 19257 28373 19291 28407
rect 20453 28373 20487 28407
rect 21189 28373 21223 28407
rect 22661 28373 22695 28407
rect 25053 28373 25087 28407
rect 26157 28373 26191 28407
rect 26449 28373 26483 28407
rect 26617 28373 26651 28407
rect 27445 28373 27479 28407
rect 27721 28373 27755 28407
rect 29285 28373 29319 28407
rect 31033 28373 31067 28407
rect 33885 28373 33919 28407
rect 41889 28373 41923 28407
rect 1685 28169 1719 28203
rect 1869 28169 1903 28203
rect 4353 28169 4387 28203
rect 4813 28169 4847 28203
rect 5917 28169 5951 28203
rect 7665 28169 7699 28203
rect 10149 28169 10183 28203
rect 10609 28169 10643 28203
rect 12081 28169 12115 28203
rect 12909 28169 12943 28203
rect 13277 28169 13311 28203
rect 15025 28169 15059 28203
rect 15485 28169 15519 28203
rect 24317 28169 24351 28203
rect 24593 28169 24627 28203
rect 28641 28169 28675 28203
rect 31953 28169 31987 28203
rect 33517 28169 33551 28203
rect 33977 28169 34011 28203
rect 1501 28101 1535 28135
rect 2237 28101 2271 28135
rect 3065 28101 3099 28135
rect 3157 28101 3191 28135
rect 5549 28101 5583 28135
rect 6469 28101 6503 28135
rect 9321 28101 9355 28135
rect 9689 28101 9723 28135
rect 10517 28101 10551 28135
rect 12449 28101 12483 28135
rect 14657 28101 14691 28135
rect 18981 28101 19015 28135
rect 19533 28101 19567 28135
rect 28978 28101 29012 28135
rect 42625 28101 42659 28135
rect 43002 28101 43036 28135
rect 1777 28033 1811 28067
rect 2329 28033 2363 28067
rect 3525 28033 3559 28067
rect 3709 28033 3743 28067
rect 4169 28033 4203 28067
rect 4445 28033 4479 28067
rect 4997 28033 5031 28067
rect 5089 28033 5123 28067
rect 5273 28033 5307 28067
rect 5461 28023 5495 28057
rect 5733 28033 5767 28067
rect 6009 28033 6043 28067
rect 6653 28033 6687 28067
rect 6745 28033 6779 28067
rect 7481 28033 7515 28067
rect 7757 28033 7791 28067
rect 8585 28033 8619 28067
rect 8861 28033 8895 28067
rect 9229 28033 9263 28067
rect 9413 28033 9447 28067
rect 9505 28033 9539 28067
rect 9781 28033 9815 28067
rect 9873 28033 9907 28067
rect 10977 28033 11011 28067
rect 11529 28033 11563 28067
rect 11713 28033 11747 28067
rect 13112 28033 13146 28067
rect 13369 28033 13403 28067
rect 13553 28033 13587 28067
rect 13645 28033 13679 28067
rect 13829 28033 13863 28067
rect 14565 28033 14599 28067
rect 14749 28033 14783 28067
rect 17601 28033 17635 28067
rect 17877 28033 17911 28067
rect 19073 28033 19107 28067
rect 19441 28033 19475 28067
rect 19717 28033 19751 28067
rect 19984 28033 20018 28067
rect 21925 28033 21959 28067
rect 22569 28033 22603 28067
rect 22937 28033 22971 28067
rect 23204 28033 23238 28067
rect 26065 28033 26099 28067
rect 26249 28033 26283 28067
rect 27169 28033 27203 28067
rect 27353 28033 27387 28067
rect 27629 28033 27663 28067
rect 27721 28033 27755 28067
rect 27905 28033 27939 28067
rect 28457 28033 28491 28067
rect 28733 28033 28767 28067
rect 32137 28033 32171 28067
rect 32404 28033 32438 28067
rect 33609 28033 33643 28067
rect 33793 28033 33827 28067
rect 43269 28033 43303 28067
rect 43361 28033 43395 28067
rect 2513 27965 2547 27999
rect 3341 27965 3375 27999
rect 5181 27965 5215 27999
rect 10793 27965 10827 27999
rect 11069 27965 11103 27999
rect 12541 27965 12575 27999
rect 12725 27965 12759 27999
rect 15577 27965 15611 27999
rect 16681 27965 16715 27999
rect 16865 27965 16899 27999
rect 17739 27965 17773 27999
rect 19165 27965 19199 27999
rect 27445 27965 27479 27999
rect 28273 27965 28307 27999
rect 30297 27965 30331 27999
rect 31309 27965 31343 27999
rect 1501 27897 1535 27931
rect 6469 27897 6503 27931
rect 10057 27897 10091 27931
rect 11621 27897 11655 27931
rect 17325 27897 17359 27931
rect 18521 27897 18555 27931
rect 21373 27897 21407 27931
rect 27261 27897 27295 27931
rect 28089 27897 28123 27931
rect 2697 27829 2731 27863
rect 3525 27829 3559 27863
rect 3985 27829 4019 27863
rect 7297 27829 7331 27863
rect 8401 27829 8435 27863
rect 8769 27829 8803 27863
rect 14381 27829 14415 27863
rect 16221 27829 16255 27863
rect 18613 27829 18647 27863
rect 21097 27829 21131 27863
rect 22477 27829 22511 27863
rect 22753 27829 22787 27863
rect 26433 27829 26467 27863
rect 26985 27829 27019 27863
rect 30113 27829 30147 27863
rect 30941 27829 30975 27863
rect 42993 27829 43027 27863
rect 43545 27829 43579 27863
rect 3617 27625 3651 27659
rect 4721 27625 4755 27659
rect 7113 27625 7147 27659
rect 8585 27625 8619 27659
rect 9781 27625 9815 27659
rect 10333 27625 10367 27659
rect 11253 27625 11287 27659
rect 11621 27625 11655 27659
rect 13829 27625 13863 27659
rect 16589 27625 16623 27659
rect 17141 27625 17175 27659
rect 18981 27625 19015 27659
rect 28733 27625 28767 27659
rect 34069 27625 34103 27659
rect 3985 27557 4019 27591
rect 5457 27557 5491 27591
rect 6377 27557 6411 27591
rect 6745 27557 6779 27591
rect 8401 27557 8435 27591
rect 13093 27557 13127 27591
rect 13737 27557 13771 27591
rect 15025 27557 15059 27591
rect 21465 27557 21499 27591
rect 22109 27557 22143 27591
rect 23489 27557 23523 27591
rect 24777 27557 24811 27591
rect 32689 27557 32723 27591
rect 33333 27557 33367 27591
rect 1869 27489 1903 27523
rect 8953 27489 8987 27523
rect 10241 27489 10275 27523
rect 11437 27489 11471 27523
rect 12265 27489 12299 27523
rect 13001 27489 13035 27523
rect 19809 27489 19843 27523
rect 21649 27489 21683 27523
rect 25053 27489 25087 27523
rect 29377 27489 29411 27523
rect 31401 27489 31435 27523
rect 1593 27421 1627 27455
rect 3065 27421 3099 27455
rect 3249 27421 3283 27455
rect 3433 27421 3467 27455
rect 4169 27421 4203 27455
rect 4261 27421 4295 27455
rect 4537 27421 4571 27455
rect 4629 27421 4663 27455
rect 4997 27421 5031 27455
rect 5089 27421 5123 27455
rect 5181 27421 5215 27455
rect 5365 27421 5399 27455
rect 5733 27421 5767 27455
rect 6745 27421 6779 27455
rect 7021 27421 7055 27455
rect 7389 27421 7423 27455
rect 7481 27421 7515 27455
rect 7573 27421 7607 27455
rect 7757 27421 7791 27455
rect 7849 27421 7883 27455
rect 8125 27421 8159 27455
rect 8217 27421 8251 27455
rect 8585 27421 8619 27455
rect 8769 27421 8803 27455
rect 9137 27421 9171 27455
rect 9229 27421 9263 27455
rect 9413 27421 9447 27455
rect 9505 27421 9539 27455
rect 9965 27421 9999 27455
rect 10149 27421 10183 27455
rect 10517 27421 10551 27455
rect 10609 27421 10643 27455
rect 10793 27421 10827 27455
rect 10885 27421 10919 27455
rect 11161 27421 11195 27455
rect 11345 27421 11379 27455
rect 12449 27421 12483 27455
rect 12541 27421 12575 27455
rect 12633 27421 12667 27455
rect 12909 27421 12943 27455
rect 13185 27421 13219 27455
rect 14197 27421 14231 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 15209 27421 15243 27455
rect 17233 27421 17267 27455
rect 17500 27421 17534 27455
rect 20085 27421 20119 27455
rect 20913 27421 20947 27455
rect 21741 27421 21775 27455
rect 24593 27421 24627 27455
rect 24869 27421 24903 27455
rect 25237 27421 25271 27455
rect 26709 27421 26743 27455
rect 26801 27421 26835 27455
rect 26893 27421 26927 27455
rect 27077 27421 27111 27455
rect 27353 27421 27387 27455
rect 27445 27421 27479 27455
rect 27629 27421 27663 27455
rect 27721 27421 27755 27455
rect 27997 27421 28031 27455
rect 28917 27421 28951 27455
rect 29009 27421 29043 27455
rect 29239 27421 29273 27455
rect 30113 27421 30147 27455
rect 30297 27421 30331 27455
rect 30389 27421 30423 27455
rect 30665 27421 30699 27455
rect 30849 27421 30883 27455
rect 30941 27421 30975 27455
rect 31033 27421 31067 27455
rect 31953 27421 31987 27455
rect 32137 27421 32171 27455
rect 32781 27421 32815 27455
rect 33057 27421 33091 27455
rect 33149 27421 33183 27455
rect 33517 27421 33551 27455
rect 33609 27421 33643 27455
rect 3341 27353 3375 27387
rect 4353 27353 4387 27387
rect 5457 27353 5491 27387
rect 8033 27353 8067 27387
rect 10977 27353 11011 27387
rect 11989 27353 12023 27387
rect 13369 27353 13403 27387
rect 14657 27353 14691 27387
rect 15476 27353 15510 27387
rect 19717 27353 19751 27387
rect 22201 27353 22235 27387
rect 26433 27353 26467 27387
rect 27813 27353 27847 27387
rect 29101 27353 29135 27387
rect 32965 27353 32999 27387
rect 5641 27285 5675 27319
rect 6009 27285 6043 27319
rect 6929 27285 6963 27319
rect 12081 27285 12115 27319
rect 12725 27285 12759 27319
rect 18613 27285 18647 27319
rect 19257 27285 19291 27319
rect 19625 27285 19659 27319
rect 20729 27285 20763 27319
rect 24409 27285 24443 27319
rect 25421 27285 25455 27319
rect 26065 27285 26099 27319
rect 27169 27285 27203 27319
rect 28181 27285 28215 27319
rect 29745 27285 29779 27319
rect 29929 27285 29963 27319
rect 31217 27285 31251 27319
rect 33793 27285 33827 27319
rect 3249 27081 3283 27115
rect 3433 27081 3467 27115
rect 5187 27081 5221 27115
rect 6193 27081 6227 27115
rect 8309 27081 8343 27115
rect 8585 27081 8619 27115
rect 8861 27081 8895 27115
rect 9321 27081 9355 27115
rect 9689 27081 9723 27115
rect 10609 27081 10643 27115
rect 10793 27081 10827 27115
rect 11161 27081 11195 27115
rect 12357 27081 12391 27115
rect 13461 27081 13495 27115
rect 13829 27081 13863 27115
rect 15301 27081 15335 27115
rect 18061 27081 18095 27115
rect 18521 27081 18555 27115
rect 23029 27081 23063 27115
rect 24317 27081 24351 27115
rect 26633 27081 26667 27115
rect 31953 27081 31987 27115
rect 33517 27081 33551 27115
rect 34253 27081 34287 27115
rect 3985 27013 4019 27047
rect 5825 27013 5859 27047
rect 6653 27013 6687 27047
rect 9229 27013 9263 27047
rect 12081 27013 12115 27047
rect 15669 27013 15703 27047
rect 16497 27013 16531 27047
rect 19432 27013 19466 27047
rect 25145 27013 25179 27047
rect 26249 27013 26283 27047
rect 26433 27013 26467 27047
rect 32404 27013 32438 27047
rect 1593 26945 1627 26979
rect 3617 26945 3651 26979
rect 3801 26945 3835 26979
rect 3893 26945 3927 26979
rect 4169 26945 4203 26979
rect 4261 26945 4295 26979
rect 4813 26945 4847 26979
rect 4905 26945 4939 26979
rect 5089 26945 5123 26979
rect 5273 26945 5307 26979
rect 5365 26945 5399 26979
rect 5549 26945 5583 26979
rect 5697 26945 5731 26979
rect 5917 26945 5951 26979
rect 6055 26945 6089 26979
rect 6377 26945 6411 26979
rect 6470 26945 6504 26979
rect 6745 26945 6779 26979
rect 6883 26945 6917 26979
rect 7757 26945 7791 26979
rect 7849 26945 7883 26979
rect 7941 26945 7975 26979
rect 8493 26945 8527 26979
rect 8769 26945 8803 26979
rect 9045 26945 9079 26979
rect 9505 26945 9539 26979
rect 9781 26945 9815 26979
rect 10517 26945 10551 26979
rect 10701 26945 10735 26979
rect 10977 26945 11011 26979
rect 11253 26945 11287 26979
rect 11713 26945 11747 26979
rect 11861 26945 11895 26979
rect 11989 26945 12023 26979
rect 12178 26945 12212 26979
rect 12909 26945 12943 26979
rect 14013 26945 14047 26979
rect 14565 26945 14599 26979
rect 15485 26945 15519 26979
rect 15761 26945 15795 26979
rect 16681 26945 16715 26979
rect 17417 26945 17451 26979
rect 18429 26945 18463 26979
rect 19165 26945 19199 26979
rect 22017 26945 22051 26979
rect 22109 26945 22143 26979
rect 22293 26945 22327 26979
rect 22753 26945 22787 26979
rect 23397 26945 23431 26979
rect 23489 26945 23523 26979
rect 24225 26945 24259 26979
rect 25053 26945 25087 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 26985 26945 27019 26979
rect 27169 26945 27203 26979
rect 27261 26945 27295 26979
rect 27445 26945 27479 26979
rect 27721 26945 27755 26979
rect 27905 26945 27939 26979
rect 28641 26945 28675 26979
rect 28819 26945 28853 26979
rect 29837 26945 29871 26979
rect 30317 26935 30351 26969
rect 30849 26945 30883 26979
rect 30941 26945 30975 26979
rect 31033 26945 31067 26979
rect 31217 26945 31251 26979
rect 31309 26945 31343 26979
rect 32137 26945 32171 26979
rect 33793 26945 33827 26979
rect 1869 26877 1903 26911
rect 4445 26877 4479 26911
rect 4629 26877 4663 26911
rect 4721 26877 4755 26911
rect 7665 26877 7699 26911
rect 9137 26877 9171 26911
rect 13185 26877 13219 26911
rect 14933 26877 14967 26911
rect 15853 26877 15887 26911
rect 16957 26877 16991 26911
rect 18613 26877 18647 26911
rect 20729 26877 20763 26911
rect 22201 26877 22235 26911
rect 23581 26877 23615 26911
rect 24409 26877 24443 26911
rect 25237 26877 25271 26911
rect 29929 26877 29963 26911
rect 30113 26877 30147 26911
rect 33609 26877 33643 26911
rect 3985 26809 4019 26843
rect 14013 26809 14047 26843
rect 16865 26809 16899 26843
rect 21833 26809 21867 26843
rect 24685 26809 24719 26843
rect 27629 26809 27663 26843
rect 29745 26809 29779 26843
rect 30481 26809 30515 26843
rect 33977 26809 34011 26843
rect 7021 26741 7055 26775
rect 7481 26741 7515 26775
rect 13001 26741 13035 26775
rect 16773 26741 16807 26775
rect 17969 26741 18003 26775
rect 20545 26741 20579 26775
rect 21373 26741 21407 26775
rect 22845 26741 22879 26775
rect 23857 26741 23891 26775
rect 25697 26741 25731 26775
rect 26617 26741 26651 26775
rect 26801 26741 26835 26775
rect 26985 26741 27019 26775
rect 27721 26741 27755 26775
rect 28089 26741 28123 26775
rect 28641 26741 28675 26775
rect 29377 26741 29411 26775
rect 30573 26741 30607 26775
rect 4169 26537 4203 26571
rect 6561 26537 6595 26571
rect 7941 26537 7975 26571
rect 8953 26537 8987 26571
rect 14841 26537 14875 26571
rect 16221 26537 16255 26571
rect 17233 26537 17267 26571
rect 18502 26537 18536 26571
rect 19625 26537 19659 26571
rect 21373 26537 21407 26571
rect 23489 26537 23523 26571
rect 24225 26537 24259 26571
rect 25145 26537 25179 26571
rect 25697 26537 25731 26571
rect 26249 26537 26283 26571
rect 28089 26537 28123 26571
rect 28825 26537 28859 26571
rect 29193 26537 29227 26571
rect 30757 26537 30791 26571
rect 33149 26537 33183 26571
rect 33885 26537 33919 26571
rect 4537 26469 4571 26503
rect 5549 26469 5583 26503
rect 9413 26469 9447 26503
rect 15025 26469 15059 26503
rect 15393 26469 15427 26503
rect 18613 26469 18647 26503
rect 30941 26469 30975 26503
rect 33425 26469 33459 26503
rect 8309 26401 8343 26435
rect 10609 26401 10643 26435
rect 11161 26401 11195 26435
rect 14657 26401 14691 26435
rect 15485 26401 15519 26435
rect 15577 26401 15611 26435
rect 15853 26401 15887 26435
rect 18705 26401 18739 26435
rect 18889 26401 18923 26435
rect 21005 26401 21039 26435
rect 21189 26401 21223 26435
rect 21649 26401 21683 26435
rect 21741 26401 21775 26435
rect 24593 26401 24627 26435
rect 26617 26401 26651 26435
rect 26893 26401 26927 26435
rect 27102 26401 27136 26435
rect 27353 26401 27387 26435
rect 27629 26401 27663 26435
rect 28181 26401 28215 26435
rect 29377 26401 29411 26435
rect 1593 26333 1627 26367
rect 4997 26333 5031 26367
rect 5181 26333 5215 26367
rect 5365 26333 5399 26367
rect 5917 26333 5951 26367
rect 6065 26333 6099 26367
rect 6193 26333 6227 26367
rect 6285 26333 6319 26367
rect 6423 26333 6457 26367
rect 7297 26333 7331 26367
rect 7390 26333 7424 26367
rect 7803 26333 7837 26367
rect 9137 26333 9171 26367
rect 9229 26333 9263 26367
rect 11621 26333 11655 26367
rect 13461 26333 13495 26367
rect 13615 26333 13649 26367
rect 13829 26333 13863 26367
rect 14841 26333 14875 26367
rect 15301 26333 15335 26367
rect 15761 26333 15795 26367
rect 17417 26333 17451 26367
rect 17601 26333 17635 26367
rect 17693 26333 17727 26367
rect 17785 26333 17819 26367
rect 19441 26333 19475 26367
rect 19881 26333 19915 26367
rect 19974 26333 20008 26367
rect 20085 26333 20119 26367
rect 20269 26333 20303 26367
rect 21557 26333 21591 26367
rect 21833 26333 21867 26367
rect 22017 26333 22051 26367
rect 23581 26333 23615 26367
rect 23729 26333 23763 26367
rect 24046 26333 24080 26367
rect 24777 26333 24811 26367
rect 25605 26333 25639 26367
rect 25789 26333 25823 26367
rect 26157 26333 26191 26367
rect 26249 26333 26283 26367
rect 27537 26333 27571 26367
rect 27721 26333 27755 26367
rect 27813 26333 27847 26367
rect 27997 26333 28031 26367
rect 28365 26333 28399 26367
rect 29101 26333 29135 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 30021 26333 30055 26367
rect 30205 26333 30239 26367
rect 30665 26333 30699 26367
rect 30757 26333 30791 26367
rect 31125 26333 31159 26367
rect 31769 26333 31803 26367
rect 2605 26265 2639 26299
rect 3249 26265 3283 26299
rect 5273 26265 5307 26299
rect 7573 26265 7607 26299
rect 7665 26265 7699 26299
rect 8677 26265 8711 26299
rect 8953 26265 8987 26299
rect 13369 26265 13403 26299
rect 14565 26265 14599 26299
rect 16957 26265 16991 26299
rect 17141 26265 17175 26299
rect 18337 26265 18371 26299
rect 23857 26265 23891 26299
rect 23949 26265 23983 26299
rect 24685 26265 24719 26299
rect 25421 26265 25455 26299
rect 28089 26265 28123 26299
rect 28641 26265 28675 26299
rect 28841 26265 28875 26299
rect 29377 26265 29411 26299
rect 30297 26265 30331 26299
rect 32036 26265 32070 26299
rect 3617 26197 3651 26231
rect 4905 26197 4939 26231
rect 6929 26197 6963 26231
rect 14381 26197 14415 26231
rect 15117 26197 15151 26231
rect 16221 26197 16255 26231
rect 16405 26197 16439 26231
rect 16681 26197 16715 26231
rect 17969 26197 18003 26231
rect 20545 26197 20579 26231
rect 20913 26197 20947 26231
rect 22385 26197 22419 26231
rect 26525 26197 26559 26231
rect 26985 26197 27019 26231
rect 27261 26197 27295 26231
rect 28549 26197 28583 26231
rect 29009 26197 29043 26231
rect 29561 26197 29595 26231
rect 31401 26197 31435 26231
rect 4997 25993 5031 26027
rect 5641 25993 5675 26027
rect 9045 25993 9079 26027
rect 9505 25993 9539 26027
rect 10333 25993 10367 26027
rect 11345 25993 11379 26027
rect 11713 25993 11747 26027
rect 13461 25993 13495 26027
rect 13829 25993 13863 26027
rect 15393 25993 15427 26027
rect 20177 25993 20211 26027
rect 20269 25993 20303 26027
rect 20637 25993 20671 26027
rect 21649 25993 21683 26027
rect 26709 25993 26743 26027
rect 33517 25993 33551 26027
rect 3709 25925 3743 25959
rect 3985 25925 4019 25959
rect 4629 25925 4663 25959
rect 8033 25925 8067 25959
rect 8401 25925 8435 25959
rect 10977 25925 11011 25959
rect 11069 25925 11103 25959
rect 11529 25925 11563 25959
rect 12173 25925 12207 25959
rect 15945 25925 15979 25959
rect 17693 25925 17727 25959
rect 24409 25925 24443 25959
rect 25697 25925 25731 25959
rect 26065 25925 26099 25959
rect 26985 25925 27019 25959
rect 27721 25925 27755 25959
rect 29806 25925 29840 25959
rect 32382 25925 32416 25959
rect 1676 25857 1710 25891
rect 3801 25857 3835 25891
rect 4073 25857 4107 25891
rect 4169 25857 4203 25891
rect 4445 25857 4479 25891
rect 4721 25857 4755 25891
rect 4813 25857 4847 25891
rect 5089 25857 5123 25891
rect 5273 25857 5307 25891
rect 5365 25857 5399 25891
rect 5503 25857 5537 25891
rect 6745 25857 6779 25891
rect 6929 25857 6963 25891
rect 7021 25857 7055 25891
rect 7113 25857 7147 25891
rect 8861 25857 8895 25891
rect 9137 25857 9171 25891
rect 10609 25857 10643 25891
rect 10793 25857 10827 25891
rect 11161 25857 11195 25891
rect 11805 25857 11839 25891
rect 13645 25857 13679 25891
rect 13921 25857 13955 25891
rect 14565 25857 14599 25891
rect 15577 25857 15611 25891
rect 15853 25857 15887 25891
rect 16129 25857 16163 25891
rect 16221 25857 16255 25891
rect 16681 25857 16715 25891
rect 17509 25857 17543 25891
rect 17877 25857 17911 25891
rect 19625 25857 19659 25891
rect 19993 25857 20027 25891
rect 20729 25857 20763 25891
rect 21097 25857 21131 25891
rect 22109 25857 22143 25891
rect 22477 25857 22511 25891
rect 22937 25857 22971 25891
rect 23305 25857 23339 25891
rect 23397 25857 23431 25891
rect 23673 25857 23707 25891
rect 24225 25857 24259 25891
rect 25881 25857 25915 25891
rect 26157 25857 26191 25891
rect 26249 25857 26283 25891
rect 28365 25857 28399 25891
rect 28549 25857 28583 25891
rect 28641 25857 28675 25891
rect 29561 25857 29595 25891
rect 32137 25857 32171 25891
rect 1409 25789 1443 25823
rect 18061 25789 18095 25823
rect 20821 25789 20855 25823
rect 23949 25789 23983 25823
rect 24593 25789 24627 25823
rect 25237 25789 25271 25823
rect 28917 25789 28951 25823
rect 31125 25789 31159 25823
rect 31401 25789 31435 25823
rect 2789 25721 2823 25755
rect 3341 25721 3375 25755
rect 4353 25721 4387 25755
rect 8861 25721 8895 25755
rect 11529 25721 11563 25755
rect 13277 25721 13311 25755
rect 15761 25721 15795 25755
rect 15945 25721 15979 25755
rect 17141 25721 17175 25755
rect 30941 25721 30975 25755
rect 6009 25653 6043 25687
rect 6653 25653 6687 25687
rect 7297 25653 7331 25687
rect 7573 25653 7607 25687
rect 8677 25653 8711 25687
rect 9873 25653 9907 25687
rect 14841 25653 14875 25687
rect 15301 25653 15335 25687
rect 16773 25653 16807 25687
rect 18337 25653 18371 25687
rect 18705 25653 18739 25687
rect 19165 25653 19199 25687
rect 19533 25653 19567 25687
rect 19993 25653 20027 25687
rect 21189 25653 21223 25687
rect 24869 25653 24903 25687
rect 26433 25653 26467 25687
rect 28365 25653 28399 25687
rect 2789 25449 2823 25483
rect 3249 25449 3283 25483
rect 3617 25449 3651 25483
rect 5641 25449 5675 25483
rect 8677 25449 8711 25483
rect 9505 25449 9539 25483
rect 10425 25449 10459 25483
rect 11989 25449 12023 25483
rect 14657 25449 14691 25483
rect 15485 25449 15519 25483
rect 15945 25449 15979 25483
rect 16313 25449 16347 25483
rect 16589 25449 16623 25483
rect 17509 25449 17543 25483
rect 17969 25449 18003 25483
rect 19625 25449 19659 25483
rect 20177 25449 20211 25483
rect 21281 25449 21315 25483
rect 21649 25449 21683 25483
rect 22937 25449 22971 25483
rect 28641 25449 28675 25483
rect 29653 25449 29687 25483
rect 32321 25449 32355 25483
rect 32505 25449 32539 25483
rect 33517 25449 33551 25483
rect 7205 25381 7239 25415
rect 7941 25381 7975 25415
rect 11069 25381 11103 25415
rect 17693 25381 17727 25415
rect 20453 25381 20487 25415
rect 21925 25381 21959 25415
rect 23305 25381 23339 25415
rect 24409 25381 24443 25415
rect 27629 25381 27663 25415
rect 31585 25381 31619 25415
rect 12909 25313 12943 25347
rect 16037 25313 16071 25347
rect 16681 25313 16715 25347
rect 26985 25313 27019 25347
rect 27997 25313 28031 25347
rect 30205 25313 30239 25347
rect 31677 25313 31711 25347
rect 32689 25313 32723 25347
rect 1409 25245 1443 25279
rect 2881 25245 2915 25279
rect 3065 25245 3099 25279
rect 3893 25245 3927 25279
rect 5089 25245 5123 25279
rect 5273 25245 5307 25279
rect 5365 25245 5399 25279
rect 5457 25245 5491 25279
rect 5733 25245 5767 25279
rect 5826 25245 5860 25279
rect 6009 25245 6043 25279
rect 6239 25245 6273 25279
rect 6469 25245 6503 25279
rect 6562 25245 6596 25279
rect 6745 25245 6779 25279
rect 6934 25245 6968 25279
rect 7389 25245 7423 25279
rect 7573 25245 7607 25279
rect 7665 25245 7699 25279
rect 8125 25245 8159 25279
rect 8309 25245 8343 25279
rect 8493 25245 8527 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9229 25245 9263 25279
rect 9321 25245 9355 25279
rect 9873 25245 9907 25279
rect 10241 25245 10275 25279
rect 10517 25245 10551 25279
rect 10701 25245 10735 25279
rect 10885 25245 10919 25279
rect 11161 25245 11195 25279
rect 11345 25245 11379 25279
rect 11437 25245 11471 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 12541 25245 12575 25279
rect 13185 25245 13219 25279
rect 13461 25245 13495 25279
rect 13829 25245 13863 25279
rect 14105 25245 14139 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 14473 25245 14507 25279
rect 14841 25245 14875 25279
rect 15025 25245 15059 25279
rect 15761 25245 15795 25279
rect 16221 25245 16255 25279
rect 16405 25245 16439 25279
rect 16497 25245 16531 25279
rect 16773 25245 16807 25279
rect 17877 25245 17911 25279
rect 18429 25245 18463 25279
rect 20085 25245 20119 25279
rect 20361 25245 20395 25279
rect 20545 25245 20579 25279
rect 20637 25245 20671 25279
rect 21097 25245 21131 25279
rect 21557 25245 21591 25279
rect 21741 25245 21775 25279
rect 22109 25245 22143 25279
rect 22201 25245 22235 25279
rect 22385 25245 22419 25279
rect 22477 25245 22511 25279
rect 23121 25245 23155 25279
rect 23213 25245 23247 25279
rect 23386 25245 23420 25279
rect 23765 25245 23799 25279
rect 23857 25245 23891 25279
rect 24041 25245 24075 25279
rect 24133 25245 24167 25279
rect 24685 25245 24719 25279
rect 24777 25245 24811 25279
rect 24961 25245 24995 25279
rect 25077 25245 25111 25279
rect 26709 25245 26743 25279
rect 26893 25245 26927 25279
rect 29009 25245 29043 25279
rect 29101 25242 29135 25276
rect 29193 25245 29227 25279
rect 29389 25245 29423 25279
rect 29561 25245 29595 25279
rect 30021 25245 30055 25279
rect 32413 25245 32447 25279
rect 32965 25245 32999 25279
rect 1676 25177 1710 25211
rect 4997 25177 5031 25211
rect 6101 25177 6135 25211
rect 6837 25177 6871 25211
rect 8401 25177 8435 25211
rect 10057 25177 10091 25211
rect 10149 25177 10183 25211
rect 10793 25177 10827 25211
rect 17141 25177 17175 25211
rect 20913 25177 20947 25211
rect 24409 25177 24443 25211
rect 24869 25177 24903 25211
rect 28733 25177 28767 25211
rect 30472 25177 30506 25211
rect 4445 25109 4479 25143
rect 6377 25109 6411 25143
rect 7113 25109 7147 25143
rect 14841 25109 14875 25143
rect 15577 25109 15611 25143
rect 16957 25109 16991 25143
rect 17518 25109 17552 25143
rect 22845 25109 22879 25143
rect 23581 25109 23615 25143
rect 24593 25109 24627 25143
rect 25145 25109 25179 25143
rect 26801 25109 26835 25143
rect 32689 25109 32723 25143
rect 1777 24905 1811 24939
rect 5365 24905 5399 24939
rect 8401 24905 8435 24939
rect 9045 24905 9079 24939
rect 10701 24905 10735 24939
rect 13461 24905 13495 24939
rect 21097 24905 21131 24939
rect 27721 24905 27755 24939
rect 30481 24905 30515 24939
rect 32781 24905 32815 24939
rect 34069 24905 34103 24939
rect 5089 24837 5123 24871
rect 5917 24837 5951 24871
rect 7297 24837 7331 24871
rect 9413 24837 9447 24871
rect 10333 24837 10367 24871
rect 13093 24837 13127 24871
rect 16037 24837 16071 24871
rect 20637 24837 20671 24871
rect 21833 24837 21867 24871
rect 23213 24837 23247 24871
rect 23949 24837 23983 24871
rect 24041 24837 24075 24871
rect 24159 24837 24193 24871
rect 24685 24837 24719 24871
rect 24777 24837 24811 24871
rect 33149 24837 33183 24871
rect 1593 24769 1627 24803
rect 2513 24769 2547 24803
rect 2605 24769 2639 24803
rect 2872 24769 2906 24803
rect 4813 24769 4847 24803
rect 4997 24769 5031 24803
rect 5181 24769 5215 24803
rect 5549 24769 5583 24803
rect 5697 24769 5731 24803
rect 5825 24769 5859 24803
rect 6055 24769 6089 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 6745 24769 6779 24803
rect 7021 24769 7055 24803
rect 7169 24769 7203 24803
rect 7389 24769 7423 24803
rect 7527 24769 7561 24803
rect 8493 24769 8527 24803
rect 8677 24769 8711 24803
rect 8769 24769 8803 24803
rect 8861 24769 8895 24803
rect 9137 24769 9171 24803
rect 9275 24769 9309 24803
rect 9505 24769 9539 24803
rect 9602 24769 9636 24803
rect 10149 24769 10183 24803
rect 10425 24769 10459 24803
rect 10517 24769 10551 24803
rect 10977 24769 11011 24803
rect 11069 24769 11103 24803
rect 11253 24769 11287 24803
rect 11345 24769 11379 24803
rect 11621 24769 11655 24803
rect 11805 24769 11839 24803
rect 11897 24769 11931 24803
rect 11989 24769 12023 24803
rect 12909 24769 12943 24803
rect 13185 24769 13219 24803
rect 13277 24769 13311 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 15301 24769 15335 24803
rect 15577 24769 15611 24803
rect 15945 24769 15979 24803
rect 16129 24769 16163 24803
rect 16267 24769 16301 24803
rect 16681 24769 16715 24803
rect 16957 24769 16991 24803
rect 17693 24769 17727 24803
rect 17877 24769 17911 24803
rect 17969 24769 18003 24803
rect 18245 24769 18279 24803
rect 18797 24769 18831 24803
rect 19533 24737 19567 24771
rect 19901 24769 19935 24803
rect 20177 24769 20211 24803
rect 20269 24769 20303 24803
rect 20821 24769 20855 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 21465 24769 21499 24803
rect 21649 24769 21683 24803
rect 22017 24769 22051 24803
rect 22201 24769 22235 24803
rect 23029 24769 23063 24803
rect 23305 24769 23339 24803
rect 23397 24769 23431 24803
rect 23857 24769 23891 24803
rect 24593 24769 24627 24803
rect 24895 24769 24929 24803
rect 26985 24769 27019 24803
rect 27077 24769 27111 24803
rect 27445 24769 27479 24803
rect 27537 24769 27571 24803
rect 27997 24769 28031 24803
rect 28181 24769 28215 24803
rect 28365 24769 28399 24803
rect 28825 24769 28859 24803
rect 29368 24769 29402 24803
rect 31217 24769 31251 24803
rect 31401 24769 31435 24803
rect 32873 24769 32907 24803
rect 33517 24769 33551 24803
rect 33609 24769 33643 24803
rect 34529 24769 34563 24803
rect 1409 24701 1443 24735
rect 1961 24701 1995 24735
rect 4077 24701 4111 24735
rect 14013 24701 14047 24735
rect 14381 24701 14415 24735
rect 16405 24701 16439 24735
rect 17141 24701 17175 24735
rect 19349 24701 19383 24735
rect 19691 24701 19725 24735
rect 24317 24701 24351 24735
rect 25053 24701 25087 24735
rect 27261 24701 27295 24735
rect 27905 24701 27939 24735
rect 28089 24701 28123 24735
rect 28457 24701 28491 24735
rect 29101 24701 29135 24735
rect 30573 24701 30607 24735
rect 32137 24701 32171 24735
rect 3985 24633 4019 24667
rect 8033 24633 8067 24667
rect 12173 24633 12207 24667
rect 14657 24633 14691 24667
rect 16773 24633 16807 24667
rect 20269 24633 20303 24667
rect 20453 24633 20487 24667
rect 20545 24633 20579 24667
rect 28917 24633 28951 24667
rect 4721 24565 4755 24599
rect 6193 24565 6227 24599
rect 6929 24565 6963 24599
rect 7665 24565 7699 24599
rect 9781 24565 9815 24599
rect 10793 24565 10827 24599
rect 12817 24565 12851 24599
rect 15761 24565 15795 24599
rect 17509 24565 17543 24599
rect 19901 24565 19935 24599
rect 22845 24565 22879 24599
rect 23581 24565 23615 24599
rect 23673 24565 23707 24599
rect 24409 24565 24443 24599
rect 27169 24565 27203 24599
rect 28365 24565 28399 24599
rect 28733 24565 28767 24599
rect 31953 24565 31987 24599
rect 33793 24565 33827 24599
rect 2881 24361 2915 24395
rect 8769 24361 8803 24395
rect 9597 24361 9631 24395
rect 11253 24361 11287 24395
rect 11897 24361 11931 24395
rect 14473 24361 14507 24395
rect 15301 24361 15335 24395
rect 15761 24361 15795 24395
rect 17877 24361 17911 24395
rect 21373 24361 21407 24395
rect 21557 24361 21591 24395
rect 22109 24361 22143 24395
rect 23397 24361 23431 24395
rect 23857 24361 23891 24395
rect 29745 24361 29779 24395
rect 30297 24361 30331 24395
rect 4445 24293 4479 24327
rect 5089 24293 5123 24327
rect 9965 24293 9999 24327
rect 10517 24293 10551 24327
rect 13921 24293 13955 24327
rect 1869 24225 1903 24259
rect 3525 24225 3559 24259
rect 12725 24225 12759 24259
rect 20913 24225 20947 24259
rect 23489 24225 23523 24259
rect 30481 24225 30515 24259
rect 32413 24225 32447 24259
rect 1593 24157 1627 24191
rect 3341 24157 3375 24191
rect 3801 24157 3835 24191
rect 4537 24157 4571 24191
rect 4813 24157 4847 24191
rect 4905 24157 4939 24191
rect 5181 24157 5215 24191
rect 5457 24157 5491 24191
rect 5549 24157 5583 24191
rect 6009 24157 6043 24191
rect 6102 24157 6136 24191
rect 6377 24157 6411 24191
rect 6493 24157 6527 24191
rect 7021 24157 7055 24191
rect 7169 24157 7203 24191
rect 7297 24157 7331 24191
rect 7527 24157 7561 24191
rect 7941 24157 7975 24191
rect 8125 24157 8159 24191
rect 8218 24157 8252 24191
rect 8631 24157 8665 24191
rect 8953 24157 8987 24191
rect 9046 24157 9080 24191
rect 9229 24157 9263 24191
rect 9459 24157 9493 24191
rect 10701 24157 10735 24191
rect 10977 24157 11011 24191
rect 11069 24157 11103 24191
rect 11345 24157 11379 24191
rect 11529 24157 11563 24191
rect 11621 24157 11655 24191
rect 11713 24157 11747 24191
rect 12909 24157 12943 24191
rect 13001 24157 13035 24191
rect 13185 24157 13219 24191
rect 13277 24157 13311 24191
rect 13369 24157 13403 24191
rect 13737 24157 13771 24191
rect 14657 24157 14691 24191
rect 14933 24157 14967 24191
rect 15577 24157 15611 24191
rect 16129 24157 16163 24191
rect 16497 24157 16531 24191
rect 16865 24157 16899 24191
rect 17233 24157 17267 24191
rect 17417 24157 17451 24191
rect 18245 24157 18279 24191
rect 18613 24157 18647 24191
rect 19073 24157 19107 24191
rect 19441 24157 19475 24191
rect 20545 24157 20579 24191
rect 21005 24157 21039 24191
rect 21373 24157 21407 24191
rect 21741 24157 21775 24191
rect 22109 24157 22143 24191
rect 22385 24157 22419 24191
rect 23673 24157 23707 24191
rect 24685 24157 24719 24191
rect 24777 24157 24811 24191
rect 24869 24157 24903 24191
rect 25053 24157 25087 24191
rect 25697 24157 25731 24191
rect 25973 24157 26007 24191
rect 26065 24157 26099 24191
rect 26341 24157 26375 24191
rect 26525 24157 26559 24191
rect 26617 24157 26651 24191
rect 26709 24157 26743 24191
rect 27445 24157 27479 24191
rect 27629 24157 27663 24191
rect 27813 24157 27847 24191
rect 30665 24157 30699 24191
rect 30941 24157 30975 24191
rect 32680 24157 32714 24191
rect 3249 24089 3283 24123
rect 4721 24089 4755 24123
rect 5365 24089 5399 24123
rect 6285 24089 6319 24123
rect 7389 24089 7423 24123
rect 8401 24089 8435 24123
rect 8493 24089 8527 24123
rect 9321 24089 9355 24123
rect 10885 24089 10919 24123
rect 12265 24089 12299 24123
rect 13553 24089 13587 24123
rect 13645 24089 13679 24123
rect 14841 24089 14875 24123
rect 15393 24089 15427 24123
rect 23397 24089 23431 24123
rect 25881 24089 25915 24123
rect 27721 24089 27755 24123
rect 28089 24089 28123 24123
rect 28917 24089 28951 24123
rect 31186 24089 31220 24123
rect 5733 24021 5767 24055
rect 6653 24021 6687 24055
rect 7665 24021 7699 24055
rect 15945 24021 15979 24055
rect 19625 24021 19659 24055
rect 21925 24021 21959 24055
rect 24409 24021 24443 24055
rect 26249 24021 26283 24055
rect 26893 24021 26927 24055
rect 27261 24021 27295 24055
rect 27997 24021 28031 24055
rect 30849 24021 30883 24055
rect 32321 24021 32355 24055
rect 33793 24021 33827 24055
rect 1961 23817 1995 23851
rect 5549 23817 5583 23851
rect 6745 23817 6779 23851
rect 7481 23817 7515 23851
rect 9137 23817 9171 23851
rect 9781 23817 9815 23851
rect 13645 23817 13679 23851
rect 14197 23817 14231 23851
rect 15209 23817 15243 23851
rect 21189 23817 21223 23851
rect 21465 23817 21499 23851
rect 23673 23817 23707 23851
rect 25513 23817 25547 23851
rect 28457 23817 28491 23851
rect 28917 23817 28951 23851
rect 30849 23817 30883 23851
rect 4813 23749 4847 23783
rect 14657 23749 14691 23783
rect 17601 23749 17635 23783
rect 20177 23749 20211 23783
rect 22293 23749 22327 23783
rect 23305 23749 23339 23783
rect 23397 23749 23431 23783
rect 24041 23749 24075 23783
rect 24961 23749 24995 23783
rect 25973 23749 26007 23783
rect 27261 23749 27295 23783
rect 27813 23749 27847 23783
rect 31677 23749 31711 23783
rect 1593 23681 1627 23715
rect 2320 23681 2354 23715
rect 3525 23681 3559 23715
rect 4445 23681 4479 23715
rect 4538 23681 4572 23715
rect 4721 23681 4755 23715
rect 4951 23681 4985 23715
rect 5641 23681 5675 23715
rect 6377 23681 6411 23715
rect 6561 23681 6595 23715
rect 8953 23681 8987 23715
rect 10793 23681 10827 23715
rect 11805 23681 11839 23715
rect 12633 23681 12667 23715
rect 13093 23681 13127 23715
rect 13277 23681 13311 23715
rect 13369 23681 13403 23715
rect 13461 23681 13495 23715
rect 14473 23681 14507 23715
rect 14933 23681 14967 23715
rect 15301 23681 15335 23715
rect 15945 23681 15979 23715
rect 16037 23681 16071 23715
rect 16405 23681 16439 23715
rect 16681 23681 16715 23715
rect 16865 23671 16899 23705
rect 16957 23681 16991 23715
rect 17141 23681 17175 23715
rect 18061 23681 18095 23715
rect 18429 23681 18463 23715
rect 18521 23671 18555 23705
rect 18955 23681 18989 23715
rect 19349 23681 19383 23715
rect 19441 23681 19475 23715
rect 19717 23681 19751 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 20913 23681 20947 23715
rect 21097 23681 21131 23715
rect 21373 23681 21407 23715
rect 21557 23681 21591 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 22385 23681 22419 23715
rect 23121 23681 23155 23715
rect 23489 23681 23523 23715
rect 23765 23681 23799 23715
rect 23949 23681 23983 23715
rect 24133 23681 24167 23715
rect 25145 23681 25179 23715
rect 25421 23681 25455 23715
rect 25697 23681 25731 23715
rect 25881 23681 25915 23715
rect 26065 23681 26099 23715
rect 26985 23681 27019 23715
rect 27169 23681 27203 23715
rect 27353 23681 27387 23715
rect 27629 23681 27663 23715
rect 27905 23681 27939 23715
rect 27997 23681 28031 23715
rect 29009 23681 29043 23715
rect 29193 23681 29227 23715
rect 29377 23681 29411 23715
rect 29745 23681 29779 23715
rect 31585 23681 31619 23715
rect 32597 23681 32631 23715
rect 1685 23613 1719 23647
rect 2053 23613 2087 23647
rect 4169 23613 4203 23647
rect 8769 23613 8803 23647
rect 10977 23613 11011 23647
rect 14841 23613 14875 23647
rect 15393 23613 15427 23647
rect 17877 23613 17911 23647
rect 29469 23613 29503 23647
rect 3433 23545 3467 23579
rect 8677 23545 8711 23579
rect 12173 23545 12207 23579
rect 18245 23545 18279 23579
rect 19533 23545 19567 23579
rect 20545 23545 20579 23579
rect 22569 23545 22603 23579
rect 25237 23545 25271 23579
rect 26709 23545 26743 23579
rect 5089 23477 5123 23511
rect 5825 23477 5859 23511
rect 6193 23477 6227 23511
rect 7021 23477 7055 23511
rect 7849 23477 7883 23511
rect 8217 23477 8251 23511
rect 10057 23477 10091 23511
rect 10609 23477 10643 23511
rect 13001 23477 13035 23511
rect 16773 23477 16807 23511
rect 17233 23477 17267 23511
rect 18061 23477 18095 23511
rect 18889 23477 18923 23511
rect 24317 23477 24351 23511
rect 25329 23477 25363 23511
rect 26249 23477 26283 23511
rect 27537 23477 27571 23511
rect 28181 23477 28215 23511
rect 33149 23477 33183 23511
rect 2881 23273 2915 23307
rect 4905 23273 4939 23307
rect 5641 23273 5675 23307
rect 8769 23273 8803 23307
rect 9137 23273 9171 23307
rect 15669 23273 15703 23307
rect 16221 23273 16255 23307
rect 17049 23273 17083 23307
rect 17141 23273 17175 23307
rect 17601 23273 17635 23307
rect 18521 23273 18555 23307
rect 19901 23273 19935 23307
rect 22109 23273 22143 23307
rect 22293 23273 22327 23307
rect 25145 23273 25179 23307
rect 32505 23273 32539 23307
rect 6377 23205 6411 23239
rect 8033 23205 8067 23239
rect 32689 23205 32723 23239
rect 33057 23205 33091 23239
rect 1869 23137 1903 23171
rect 3341 23137 3375 23171
rect 3525 23137 3559 23171
rect 4169 23137 4203 23171
rect 11529 23137 11563 23171
rect 17233 23137 17267 23171
rect 25053 23137 25087 23171
rect 27629 23137 27663 23171
rect 28365 23137 28399 23171
rect 28825 23137 28859 23171
rect 32413 23137 32447 23171
rect 1593 23069 1627 23103
rect 3249 23069 3283 23103
rect 4261 23069 4295 23103
rect 4409 23069 4443 23103
rect 4537 23069 4571 23103
rect 4726 23069 4760 23103
rect 4997 23069 5031 23103
rect 5090 23069 5124 23103
rect 5273 23069 5307 23103
rect 5365 23069 5399 23103
rect 5462 23069 5496 23103
rect 5733 23069 5767 23103
rect 5826 23069 5860 23103
rect 6101 23069 6135 23103
rect 6198 23069 6232 23103
rect 6929 23069 6963 23103
rect 7022 23069 7056 23103
rect 7205 23069 7239 23103
rect 7394 23069 7428 23103
rect 9321 23069 9355 23103
rect 10793 23069 10827 23103
rect 11069 23069 11103 23103
rect 11253 23069 11287 23103
rect 11621 23069 11655 23103
rect 11897 23069 11931 23103
rect 11990 23069 12024 23103
rect 12173 23069 12207 23103
rect 12403 23069 12437 23103
rect 12633 23069 12667 23103
rect 13001 23069 13035 23103
rect 13277 23069 13311 23103
rect 14565 23069 14599 23103
rect 17417 23069 17451 23103
rect 17785 23069 17819 23103
rect 18061 23069 18095 23103
rect 18245 23069 18279 23103
rect 18441 23069 18475 23103
rect 18705 23069 18739 23103
rect 18797 23069 18831 23103
rect 18889 23069 18923 23103
rect 19073 23069 19107 23103
rect 19349 23069 19383 23103
rect 19993 23069 20027 23103
rect 20177 23069 20211 23103
rect 20361 23069 20395 23103
rect 20499 23069 20533 23103
rect 20637 23069 20671 23103
rect 20729 23069 20763 23103
rect 20821 23069 20855 23103
rect 21005 23069 21039 23103
rect 21557 23069 21591 23103
rect 21649 23069 21683 23103
rect 21741 23069 21775 23103
rect 21833 23069 21867 23103
rect 22017 23069 22051 23103
rect 22109 23069 22143 23103
rect 22661 23069 22695 23103
rect 23213 23069 23247 23103
rect 23673 23069 23707 23103
rect 25145 23069 25179 23103
rect 25789 23069 25823 23103
rect 25882 23069 25916 23103
rect 26157 23069 26191 23103
rect 26295 23069 26329 23103
rect 26525 23069 26559 23103
rect 26709 23069 26743 23103
rect 26801 23069 26835 23103
rect 26893 23069 26927 23103
rect 27997 23069 28031 23103
rect 28089 23069 28123 23103
rect 28733 23069 28767 23103
rect 32137 23069 32171 23103
rect 3801 23001 3835 23035
rect 3985 23001 4019 23035
rect 4629 23001 4663 23035
rect 6009 23001 6043 23035
rect 7297 23001 7331 23035
rect 9588 23001 9622 23035
rect 12262 23001 12296 23035
rect 12817 23001 12851 23035
rect 12909 23001 12943 23035
rect 13553 23001 13587 23035
rect 14381 23001 14415 23035
rect 16589 23001 16623 23035
rect 17141 23001 17175 23035
rect 18337 23001 18371 23035
rect 18521 23001 18555 23035
rect 23949 23001 23983 23035
rect 24869 23001 24903 23035
rect 26065 23001 26099 23035
rect 6653 22933 6687 22967
rect 7573 22933 7607 22967
rect 8309 22933 8343 22967
rect 10701 22933 10735 22967
rect 10885 22933 10919 22967
rect 12541 22933 12575 22967
rect 13185 22933 13219 22967
rect 14657 22933 14691 22967
rect 15393 22933 15427 22967
rect 17877 22933 17911 22967
rect 18981 22933 19015 22967
rect 20085 22933 20119 22967
rect 21189 22933 21223 22967
rect 22937 22933 22971 22967
rect 23305 22933 23339 22967
rect 25329 22933 25363 22967
rect 26433 22933 26467 22967
rect 27077 22933 27111 22967
rect 28273 22933 28307 22967
rect 29009 22933 29043 22967
rect 3525 22729 3559 22763
rect 8953 22729 8987 22763
rect 10333 22729 10367 22763
rect 13185 22729 13219 22763
rect 15577 22729 15611 22763
rect 17325 22729 17359 22763
rect 19901 22729 19935 22763
rect 21557 22729 21591 22763
rect 23489 22729 23523 22763
rect 25973 22729 26007 22763
rect 28181 22729 28215 22763
rect 28549 22729 28583 22763
rect 7205 22661 7239 22695
rect 7297 22661 7331 22695
rect 7941 22661 7975 22695
rect 8033 22661 8067 22695
rect 9321 22661 9355 22695
rect 12173 22661 12207 22695
rect 18705 22661 18739 22695
rect 21833 22661 21867 22695
rect 24685 22661 24719 22695
rect 25513 22661 25547 22695
rect 27169 22661 27203 22695
rect 27353 22661 27387 22695
rect 27905 22661 27939 22695
rect 29101 22661 29135 22695
rect 1676 22593 1710 22627
rect 4537 22593 4571 22627
rect 4630 22593 4664 22627
rect 4813 22593 4847 22627
rect 4905 22593 4939 22627
rect 5043 22593 5077 22627
rect 5549 22593 5583 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 5917 22593 5951 22627
rect 6009 22593 6043 22627
rect 6929 22593 6963 22627
rect 7022 22593 7056 22627
rect 7435 22593 7469 22627
rect 7665 22593 7699 22627
rect 7813 22593 7847 22627
rect 8171 22593 8205 22627
rect 8769 22593 8803 22627
rect 8953 22593 8987 22627
rect 9045 22593 9079 22627
rect 9229 22593 9263 22627
rect 9413 22593 9447 22627
rect 10425 22593 10459 22627
rect 10573 22593 10607 22627
rect 10701 22593 10735 22627
rect 10793 22593 10827 22627
rect 10890 22593 10924 22627
rect 12633 22593 12667 22627
rect 13369 22593 13403 22627
rect 13737 22593 13771 22627
rect 13921 22593 13955 22627
rect 14473 22593 14507 22627
rect 14657 22593 14691 22627
rect 14749 22593 14783 22627
rect 14933 22593 14967 22627
rect 15485 22593 15519 22627
rect 15669 22593 15703 22627
rect 16037 22593 16071 22627
rect 16681 22593 16715 22627
rect 18061 22593 18095 22627
rect 18245 22593 18279 22627
rect 18981 22593 19015 22627
rect 19257 22593 19291 22627
rect 19441 22593 19475 22627
rect 19809 22593 19843 22627
rect 19993 22593 20027 22627
rect 20085 22593 20119 22627
rect 20269 22593 20303 22627
rect 20361 22593 20395 22627
rect 20545 22593 20579 22627
rect 20821 22593 20855 22627
rect 21005 22593 21039 22627
rect 21097 22593 21131 22627
rect 21281 22593 21315 22627
rect 22109 22593 22143 22627
rect 22477 22593 22511 22627
rect 22661 22593 22695 22627
rect 22753 22593 22787 22627
rect 22845 22593 22879 22627
rect 23213 22593 23247 22627
rect 23857 22593 23891 22627
rect 23949 22593 23983 22627
rect 24133 22593 24167 22627
rect 24225 22593 24259 22627
rect 24409 22593 24443 22627
rect 24593 22593 24627 22627
rect 24777 22593 24811 22627
rect 25789 22593 25823 22627
rect 27629 22593 27663 22627
rect 27813 22593 27847 22627
rect 27997 22593 28031 22627
rect 28273 22593 28307 22627
rect 28457 22593 28491 22627
rect 28917 22593 28951 22627
rect 1409 22525 1443 22559
rect 2973 22525 3007 22559
rect 3709 22525 3743 22559
rect 8677 22525 8711 22559
rect 9781 22525 9815 22559
rect 11529 22525 11563 22559
rect 12449 22525 12483 22559
rect 12541 22525 12575 22559
rect 12725 22525 12759 22559
rect 15117 22525 15151 22559
rect 17049 22525 17083 22559
rect 18797 22525 18831 22559
rect 21925 22525 21959 22559
rect 25605 22525 25639 22559
rect 2789 22457 2823 22491
rect 6837 22457 6871 22491
rect 9597 22457 9631 22491
rect 16957 22457 16991 22491
rect 20085 22457 20119 22491
rect 21097 22457 21131 22491
rect 23029 22457 23063 22491
rect 4261 22389 4295 22423
rect 5181 22389 5215 22423
rect 6193 22389 6227 22423
rect 7573 22389 7607 22423
rect 8309 22389 8343 22423
rect 11069 22389 11103 22423
rect 12265 22389 12299 22423
rect 16405 22389 16439 22423
rect 16846 22389 16880 22423
rect 17877 22389 17911 22423
rect 18337 22389 18371 22423
rect 18705 22389 18739 22423
rect 19165 22389 19199 22423
rect 19625 22389 19659 22423
rect 20361 22389 20395 22423
rect 20821 22389 20855 22423
rect 21833 22389 21867 22423
rect 22293 22389 22327 22423
rect 23673 22389 23707 22423
rect 24961 22389 24995 22423
rect 25789 22389 25823 22423
rect 27537 22389 27571 22423
rect 29285 22389 29319 22423
rect 3617 22185 3651 22219
rect 5365 22185 5399 22219
rect 8401 22185 8435 22219
rect 9229 22185 9263 22219
rect 10241 22185 10275 22219
rect 11069 22185 11103 22219
rect 16865 22185 16899 22219
rect 18613 22185 18647 22219
rect 19441 22185 19475 22219
rect 19809 22185 19843 22219
rect 20269 22185 20303 22219
rect 21097 22185 21131 22219
rect 24225 22185 24259 22219
rect 25789 22185 25823 22219
rect 26709 22185 26743 22219
rect 27445 22185 27479 22219
rect 27997 22185 28031 22219
rect 28733 22185 28767 22219
rect 6009 22117 6043 22151
rect 6745 22117 6779 22151
rect 9965 22117 9999 22151
rect 11897 22117 11931 22151
rect 17325 22117 17359 22151
rect 18521 22117 18555 22151
rect 19073 22117 19107 22151
rect 1869 22049 1903 22083
rect 4169 22049 4203 22083
rect 10885 22049 10919 22083
rect 15577 22049 15611 22083
rect 16957 22049 16991 22083
rect 17693 22049 17727 22083
rect 17877 22049 17911 22083
rect 18797 22049 18831 22083
rect 19533 22049 19567 22083
rect 20177 22049 20211 22083
rect 21005 22049 21039 22083
rect 21465 22049 21499 22083
rect 26709 22049 26743 22083
rect 27353 22049 27387 22083
rect 27813 22049 27847 22083
rect 1593 21981 1627 22015
rect 3065 21981 3099 22015
rect 3801 21981 3835 22015
rect 3985 21981 4019 22015
rect 4813 21981 4847 22015
rect 5089 21981 5123 22015
rect 5181 21981 5215 22015
rect 5457 21981 5491 22015
rect 5641 21981 5675 22015
rect 5825 21981 5859 22015
rect 6101 21981 6135 22015
rect 6194 21981 6228 22015
rect 6585 21981 6619 22015
rect 7849 21981 7883 22015
rect 8217 21981 8251 22015
rect 8585 21981 8619 22015
rect 8769 21981 8803 22015
rect 9321 21981 9355 22015
rect 9414 21981 9448 22015
rect 9597 21981 9631 22015
rect 9689 21981 9723 22015
rect 9827 21981 9861 22015
rect 10425 21981 10459 22015
rect 10517 21981 10551 22015
rect 10727 21981 10761 22015
rect 10977 21981 11011 22015
rect 11161 21981 11195 22015
rect 11345 21981 11379 22015
rect 11713 21981 11747 22015
rect 11989 21981 12023 22015
rect 12137 21981 12171 22015
rect 12265 21981 12299 22015
rect 12495 21981 12529 22015
rect 13277 21981 13311 22015
rect 13370 21981 13404 22015
rect 13553 21981 13587 22015
rect 13645 21981 13679 22015
rect 13742 21981 13776 22015
rect 14105 21981 14139 22015
rect 14933 21981 14967 22015
rect 15117 21981 15151 22015
rect 15209 21981 15243 22015
rect 15393 21981 15427 22015
rect 16037 21981 16071 22015
rect 17141 21981 17175 22015
rect 17601 21981 17635 22015
rect 17785 21981 17819 22015
rect 18889 21981 18923 22015
rect 19257 21981 19291 22015
rect 20269 21981 20303 22015
rect 20637 21981 20671 22015
rect 20815 21981 20849 22015
rect 20913 21981 20947 22015
rect 21373 21981 21407 22015
rect 21557 21981 21591 22015
rect 22661 21981 22695 22015
rect 23213 21981 23247 22015
rect 23581 21981 23615 22015
rect 24409 21981 24443 22015
rect 24502 21981 24536 22015
rect 24774 21981 24808 22015
rect 24874 21981 24908 22015
rect 25145 21981 25179 22015
rect 25238 21981 25272 22015
rect 25513 21981 25547 22015
rect 25610 21981 25644 22015
rect 25881 21981 25915 22015
rect 25974 21981 26008 22015
rect 26249 21981 26283 22015
rect 26346 21981 26380 22015
rect 26617 21981 26651 22015
rect 26893 21981 26927 22015
rect 27261 21981 27295 22015
rect 27721 21981 27755 22015
rect 27997 21981 28031 22015
rect 28273 21981 28307 22015
rect 28457 21981 28491 22015
rect 28733 21981 28767 22015
rect 28825 21981 28859 22015
rect 4721 21913 4755 21947
rect 4997 21913 5031 21947
rect 5733 21913 5767 21947
rect 6377 21913 6411 21947
rect 6469 21913 6503 21947
rect 6837 21913 6871 21947
rect 7573 21913 7607 21947
rect 8033 21913 8067 21947
rect 8125 21913 8159 21947
rect 10609 21913 10643 21947
rect 11529 21913 11563 21947
rect 11621 21913 11655 21947
rect 12357 21913 12391 21947
rect 16497 21913 16531 21947
rect 16865 21913 16899 21947
rect 18613 21913 18647 21947
rect 19993 21913 20027 21947
rect 20729 21913 20763 21947
rect 22937 21913 22971 21947
rect 23397 21913 23431 21947
rect 23489 21913 23523 21947
rect 24685 21913 24719 21947
rect 25421 21913 25455 21947
rect 26157 21913 26191 21947
rect 3985 21845 4019 21879
rect 8769 21845 8803 21879
rect 12633 21845 12667 21879
rect 13185 21845 13219 21879
rect 13921 21845 13955 21879
rect 16221 21845 16255 21879
rect 20453 21845 20487 21879
rect 21281 21845 21315 21879
rect 21833 21845 21867 21879
rect 22569 21845 22603 21879
rect 23765 21845 23799 21879
rect 25053 21845 25087 21879
rect 26525 21845 26559 21879
rect 27077 21845 27111 21879
rect 27629 21845 27663 21879
rect 28181 21845 28215 21879
rect 28641 21845 28675 21879
rect 29101 21845 29135 21879
rect 1501 21641 1535 21675
rect 3801 21641 3835 21675
rect 5641 21641 5675 21675
rect 5825 21641 5859 21675
rect 5917 21641 5951 21675
rect 9505 21641 9539 21675
rect 10885 21641 10919 21675
rect 11161 21641 11195 21675
rect 11345 21641 11379 21675
rect 13277 21641 13311 21675
rect 14565 21641 14599 21675
rect 16313 21641 16347 21675
rect 17141 21641 17175 21675
rect 17693 21641 17727 21675
rect 18889 21641 18923 21675
rect 21281 21641 21315 21675
rect 25973 21641 26007 21675
rect 26617 21641 26651 21675
rect 1961 21573 1995 21607
rect 2596 21573 2630 21607
rect 5273 21573 5307 21607
rect 7205 21573 7239 21607
rect 7757 21573 7791 21607
rect 8309 21573 8343 21607
rect 8401 21573 8435 21607
rect 10149 21573 10183 21607
rect 10517 21573 10551 21607
rect 11713 21573 11747 21607
rect 12909 21573 12943 21607
rect 13645 21573 13679 21607
rect 15853 21573 15887 21607
rect 22477 21573 22511 21607
rect 24501 21573 24535 21607
rect 24593 21573 24627 21607
rect 25513 21573 25547 21607
rect 26157 21573 26191 21607
rect 1869 21505 1903 21539
rect 3985 21505 4019 21539
rect 4077 21505 4111 21539
rect 4169 21505 4203 21539
rect 4287 21505 4321 21539
rect 4445 21505 4479 21539
rect 4629 21505 4663 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 5090 21505 5124 21539
rect 5365 21505 5399 21539
rect 5462 21505 5496 21539
rect 5733 21505 5767 21539
rect 6469 21505 6503 21539
rect 7481 21505 7515 21539
rect 7665 21505 7699 21539
rect 7849 21505 7883 21539
rect 8125 21505 8159 21539
rect 8493 21505 8527 21539
rect 8953 21505 8987 21539
rect 9137 21505 9171 21539
rect 9229 21505 9263 21539
rect 9367 21505 9401 21539
rect 10977 21505 11011 21539
rect 11069 21505 11103 21539
rect 12081 21505 12115 21539
rect 12633 21505 12667 21539
rect 12725 21505 12759 21539
rect 13001 21505 13035 21539
rect 13093 21505 13127 21539
rect 13369 21505 13403 21539
rect 13517 21505 13551 21539
rect 13737 21505 13771 21539
rect 13834 21505 13868 21539
rect 14105 21505 14139 21539
rect 14381 21505 14415 21539
rect 15117 21505 15151 21539
rect 15209 21505 15243 21539
rect 15393 21505 15427 21539
rect 15485 21505 15519 21539
rect 16129 21505 16163 21539
rect 16681 21505 16715 21539
rect 16957 21505 16991 21539
rect 17233 21505 17267 21539
rect 17509 21505 17543 21539
rect 17969 21505 18003 21539
rect 18153 21505 18187 21539
rect 18429 21505 18463 21539
rect 18705 21505 18739 21539
rect 18981 21505 19015 21539
rect 19165 21505 19199 21539
rect 19257 21505 19291 21539
rect 19717 21505 19751 21539
rect 19901 21505 19935 21539
rect 20018 21505 20052 21539
rect 20269 21505 20303 21539
rect 20637 21505 20671 21539
rect 21189 21505 21223 21539
rect 21373 21505 21407 21539
rect 21925 21505 21959 21539
rect 22201 21505 22235 21539
rect 22385 21505 22419 21539
rect 22569 21505 22603 21539
rect 22865 21505 22899 21539
rect 23029 21505 23063 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 23673 21505 23707 21539
rect 23949 21505 23983 21539
rect 24317 21505 24351 21539
rect 24685 21505 24719 21539
rect 25789 21505 25823 21539
rect 26433 21505 26467 21539
rect 26985 21505 27019 21539
rect 27261 21505 27295 21539
rect 27721 21505 27755 21539
rect 27905 21505 27939 21539
rect 27997 21505 28031 21539
rect 28278 21505 28312 21539
rect 28457 21505 28491 21539
rect 2145 21437 2179 21471
rect 2329 21437 2363 21471
rect 6101 21437 6135 21471
rect 11345 21437 11379 21471
rect 14197 21437 14231 21471
rect 16037 21437 16071 21471
rect 16865 21437 16899 21471
rect 17325 21437 17359 21471
rect 18521 21437 18555 21471
rect 20177 21437 20211 21471
rect 20821 21437 20855 21471
rect 23765 21437 23799 21471
rect 25605 21437 25639 21471
rect 26341 21437 26375 21471
rect 27077 21437 27111 21471
rect 3709 21369 3743 21403
rect 5825 21369 5859 21403
rect 19441 21369 19475 21403
rect 20453 21369 20487 21403
rect 23397 21369 23431 21403
rect 24133 21369 24167 21403
rect 28641 21369 28675 21403
rect 4905 21301 4939 21335
rect 8033 21301 8067 21335
rect 8677 21301 8711 21335
rect 14013 21301 14047 21335
rect 14933 21301 14967 21335
rect 15853 21301 15887 21335
rect 16681 21301 16715 21335
rect 17509 21301 17543 21335
rect 17969 21301 18003 21335
rect 18337 21301 18371 21335
rect 18521 21301 18555 21335
rect 19073 21301 19107 21335
rect 19717 21301 19751 21335
rect 20269 21301 20303 21335
rect 22017 21301 22051 21335
rect 22753 21301 22787 21335
rect 23949 21301 23983 21335
rect 24869 21301 24903 21335
rect 25789 21301 25823 21335
rect 26433 21301 26467 21335
rect 27169 21301 27203 21335
rect 27445 21301 27479 21335
rect 27997 21301 28031 21335
rect 28181 21301 28215 21335
rect 28457 21301 28491 21335
rect 3617 21097 3651 21131
rect 5365 21097 5399 21131
rect 8769 21097 8803 21131
rect 11897 21097 11931 21131
rect 12357 21097 12391 21131
rect 16957 21097 16991 21131
rect 17325 21097 17359 21131
rect 19625 21097 19659 21131
rect 20545 21097 20579 21131
rect 21833 21097 21867 21131
rect 23121 21097 23155 21131
rect 24041 21097 24075 21131
rect 25329 21097 25363 21131
rect 26525 21097 26559 21131
rect 27261 21097 27295 21131
rect 28089 21097 28123 21131
rect 28273 21097 28307 21131
rect 28457 21097 28491 21131
rect 30941 21097 30975 21131
rect 7389 21029 7423 21063
rect 14749 21029 14783 21063
rect 17969 21029 18003 21063
rect 18245 21029 18279 21063
rect 18337 21029 18371 21063
rect 20729 21029 20763 21063
rect 21465 21029 21499 21063
rect 1869 20961 1903 20995
rect 4353 20961 4387 20995
rect 4813 20961 4847 20995
rect 5181 20961 5215 20995
rect 6377 20961 6411 20995
rect 7573 20961 7607 20995
rect 12909 20961 12943 20995
rect 13093 20961 13127 20995
rect 16589 20961 16623 20995
rect 20085 20961 20119 20995
rect 26617 20961 26651 20995
rect 27353 20961 27387 20995
rect 1593 20893 1627 20927
rect 3065 20893 3099 20927
rect 3249 20893 3283 20927
rect 3341 20893 3375 20927
rect 3433 20893 3467 20927
rect 4077 20893 4111 20927
rect 4537 20893 4571 20927
rect 4905 20893 4939 20927
rect 5641 20893 5675 20927
rect 5825 20893 5859 20927
rect 6469 20893 6503 20927
rect 6653 20893 6687 20927
rect 6745 20893 6779 20927
rect 6838 20893 6872 20927
rect 7021 20893 7055 20927
rect 7113 20893 7147 20927
rect 7210 20893 7244 20927
rect 8217 20893 8251 20927
rect 8493 20893 8527 20927
rect 8585 20893 8619 20927
rect 8953 20893 8987 20927
rect 9046 20893 9080 20927
rect 9229 20893 9263 20927
rect 9321 20893 9355 20927
rect 9418 20893 9452 20927
rect 9781 20893 9815 20927
rect 10057 20893 10091 20927
rect 10149 20893 10183 20927
rect 10425 20893 10459 20927
rect 10573 20893 10607 20927
rect 10701 20893 10735 20927
rect 10890 20893 10924 20927
rect 11253 20893 11287 20927
rect 11437 20893 11471 20927
rect 12449 20893 12483 20927
rect 12633 20893 12667 20927
rect 13001 20893 13035 20927
rect 13185 20893 13219 20927
rect 13553 20893 13587 20927
rect 13829 20893 13863 20927
rect 14105 20893 14139 20927
rect 14657 20893 14691 20927
rect 14841 20893 14875 20927
rect 15209 20893 15243 20927
rect 15485 20893 15519 20927
rect 15669 20893 15703 20927
rect 16037 20893 16071 20927
rect 16865 20893 16899 20927
rect 17325 20893 17359 20927
rect 17509 20893 17543 20927
rect 17785 20893 17819 20927
rect 17877 20893 17911 20927
rect 18245 20893 18279 20927
rect 18705 20893 18739 20927
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 19533 20893 19567 20927
rect 19725 20887 19759 20921
rect 20177 20893 20211 20927
rect 20361 20893 20395 20927
rect 20637 20893 20671 20927
rect 20913 20893 20947 20927
rect 21465 20893 21499 20927
rect 21649 20893 21683 20927
rect 22017 20893 22051 20927
rect 22109 20893 22143 20927
rect 22293 20893 22327 20927
rect 22385 20893 22419 20927
rect 22569 20893 22603 20927
rect 22845 20893 22879 20927
rect 22937 20893 22971 20927
rect 23213 20893 23247 20927
rect 23397 20893 23431 20927
rect 23489 20893 23523 20927
rect 23581 20893 23615 20927
rect 24409 20893 24443 20927
rect 24502 20893 24536 20927
rect 24777 20893 24811 20927
rect 24913 20893 24947 20927
rect 25145 20893 25179 20927
rect 25329 20893 25363 20927
rect 25421 20893 25455 20927
rect 26065 20893 26099 20927
rect 26157 20893 26191 20927
rect 26341 20893 26375 20927
rect 26433 20893 26467 20927
rect 26525 20893 26559 20927
rect 27537 20893 27571 20927
rect 27813 20893 27847 20927
rect 27997 20893 28031 20927
rect 28089 20893 28123 20927
rect 28365 20893 28399 20927
rect 28733 20893 28767 20927
rect 29561 20893 29595 20927
rect 4169 20825 4203 20859
rect 5549 20825 5583 20859
rect 8401 20825 8435 20859
rect 9965 20825 9999 20859
rect 10793 20825 10827 20859
rect 14381 20825 14415 20859
rect 16681 20825 16715 20859
rect 18521 20825 18555 20859
rect 22753 20825 22787 20859
rect 23857 20825 23891 20859
rect 24057 20825 24091 20859
rect 24685 20825 24719 20859
rect 25881 20825 25915 20859
rect 27261 20825 27295 20859
rect 29806 20825 29840 20859
rect 6653 20757 6687 20791
rect 8125 20757 8159 20791
rect 9597 20757 9631 20791
rect 10333 20757 10367 20791
rect 11069 20757 11103 20791
rect 11437 20757 11471 20791
rect 12541 20757 12575 20791
rect 12725 20757 12759 20791
rect 13369 20757 13403 20791
rect 13737 20757 13771 20791
rect 15025 20757 15059 20791
rect 15393 20757 15427 20791
rect 15853 20757 15887 20791
rect 21097 20757 21131 20791
rect 23765 20757 23799 20791
rect 24225 20757 24259 20791
rect 25053 20757 25087 20791
rect 25605 20757 25639 20791
rect 26893 20757 26927 20791
rect 27721 20757 27755 20791
rect 28917 20757 28951 20791
rect 1685 20553 1719 20587
rect 6377 20553 6411 20587
rect 10609 20553 10643 20587
rect 11989 20553 12023 20587
rect 12081 20553 12115 20587
rect 13737 20553 13771 20587
rect 14565 20553 14599 20587
rect 16037 20553 16071 20587
rect 17049 20553 17083 20587
rect 18429 20553 18463 20587
rect 19165 20553 19199 20587
rect 19533 20553 19567 20587
rect 22201 20553 22235 20587
rect 24501 20553 24535 20587
rect 26709 20553 26743 20587
rect 28641 20553 28675 20587
rect 3709 20485 3743 20519
rect 5080 20485 5114 20519
rect 6863 20485 6897 20519
rect 8401 20485 8435 20519
rect 10057 20485 10091 20519
rect 10517 20485 10551 20519
rect 14924 20485 14958 20519
rect 19901 20485 19935 20519
rect 20177 20485 20211 20519
rect 25145 20485 25179 20519
rect 27169 20485 27203 20519
rect 1501 20417 1535 20451
rect 1685 20417 1719 20451
rect 2044 20417 2078 20451
rect 3617 20417 3651 20451
rect 4169 20417 4203 20451
rect 4813 20417 4847 20451
rect 6561 20417 6595 20451
rect 6653 20417 6687 20451
rect 6746 20417 6780 20451
rect 7021 20417 7055 20451
rect 7297 20417 7331 20451
rect 7750 20407 7784 20441
rect 7849 20417 7883 20451
rect 7960 20417 7994 20451
rect 8125 20417 8159 20451
rect 8493 20417 8527 20451
rect 8677 20417 8711 20451
rect 9045 20417 9079 20451
rect 9137 20417 9171 20451
rect 9597 20417 9631 20451
rect 9689 20417 9723 20451
rect 9781 20417 9815 20451
rect 9965 20417 9999 20451
rect 10149 20417 10183 20451
rect 10425 20417 10459 20451
rect 10793 20417 10827 20451
rect 10891 20417 10925 20451
rect 11069 20417 11103 20451
rect 11897 20417 11931 20451
rect 12357 20417 12391 20451
rect 12624 20417 12658 20451
rect 13829 20417 13863 20451
rect 14657 20417 14691 20451
rect 16313 20417 16347 20451
rect 16497 20417 16531 20451
rect 16681 20417 16715 20451
rect 17509 20417 17543 20451
rect 17877 20417 17911 20451
rect 18245 20417 18279 20451
rect 18797 20417 18831 20451
rect 19349 20417 19383 20451
rect 19533 20417 19567 20451
rect 20085 20417 20119 20451
rect 20269 20417 20303 20451
rect 20637 20417 20671 20451
rect 22569 20417 22603 20451
rect 22661 20417 22695 20451
rect 22845 20417 22879 20451
rect 22937 20417 22971 20451
rect 23305 20417 23339 20451
rect 23581 20417 23615 20451
rect 24777 20417 24811 20451
rect 24925 20417 24959 20451
rect 25053 20417 25087 20451
rect 25242 20417 25276 20451
rect 25789 20417 25823 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 27445 20417 27479 20451
rect 27721 20417 27755 20451
rect 27997 20417 28031 20451
rect 28273 20417 28307 20451
rect 28457 20417 28491 20451
rect 1777 20349 1811 20383
rect 3801 20349 3835 20383
rect 7389 20349 7423 20383
rect 7481 20349 7515 20383
rect 7573 20349 7607 20383
rect 8217 20349 8251 20383
rect 9505 20349 9539 20383
rect 12265 20349 12299 20383
rect 16773 20349 16807 20383
rect 23397 20349 23431 20383
rect 24041 20349 24075 20383
rect 25881 20349 25915 20383
rect 26433 20349 26467 20383
rect 27261 20349 27295 20383
rect 27813 20349 27847 20383
rect 3157 20281 3191 20315
rect 7113 20281 7147 20315
rect 9321 20281 9355 20315
rect 26249 20281 26283 20315
rect 27629 20281 27663 20315
rect 3249 20213 3283 20247
rect 4721 20213 4755 20247
rect 6193 20213 6227 20247
rect 8033 20213 8067 20247
rect 10517 20213 10551 20247
rect 10977 20213 11011 20247
rect 11805 20213 11839 20247
rect 12173 20213 12207 20247
rect 14013 20213 14047 20247
rect 16313 20213 16347 20247
rect 16865 20213 16899 20247
rect 21189 20213 21223 20247
rect 21557 20213 21591 20247
rect 22385 20213 22419 20247
rect 23581 20213 23615 20247
rect 23765 20213 23799 20247
rect 25421 20213 25455 20247
rect 25789 20213 25823 20247
rect 26525 20213 26559 20247
rect 27169 20213 27203 20247
rect 27997 20213 28031 20247
rect 28181 20213 28215 20247
rect 28365 20213 28399 20247
rect 3617 20009 3651 20043
rect 5365 20009 5399 20043
rect 9597 20009 9631 20043
rect 11897 20009 11931 20043
rect 13277 20009 13311 20043
rect 13921 20009 13955 20043
rect 18705 20009 18739 20043
rect 21465 20009 21499 20043
rect 22109 20009 22143 20043
rect 25421 20009 25455 20043
rect 25789 20009 25823 20043
rect 26893 20009 26927 20043
rect 27537 20009 27571 20043
rect 27905 20009 27939 20043
rect 28181 20009 28215 20043
rect 5825 19941 5859 19975
rect 6377 19941 6411 19975
rect 8769 19941 8803 19975
rect 11161 19941 11195 19975
rect 14197 19941 14231 19975
rect 16221 19941 16255 19975
rect 17601 19941 17635 19975
rect 20177 19941 20211 19975
rect 27353 19941 27387 19975
rect 1869 19873 1903 19907
rect 3065 19873 3099 19907
rect 4077 19873 4111 19907
rect 4721 19873 4755 19907
rect 9045 19873 9079 19907
rect 9781 19873 9815 19907
rect 11253 19873 11287 19907
rect 12357 19873 12391 19907
rect 14381 19873 14415 19907
rect 16037 19873 16071 19907
rect 18153 19873 18187 19907
rect 19717 19873 19751 19907
rect 20729 19873 20763 19907
rect 25421 19873 25455 19907
rect 26985 19873 27019 19907
rect 27537 19873 27571 19907
rect 1593 19805 1627 19839
rect 4813 19805 4847 19839
rect 4997 19805 5031 19839
rect 5089 19805 5123 19839
rect 5181 19805 5215 19839
rect 5457 19805 5491 19839
rect 5641 19805 5675 19839
rect 6285 19805 6319 19839
rect 6561 19805 6595 19839
rect 6745 19805 6779 19839
rect 7085 19805 7119 19839
rect 7297 19805 7331 19839
rect 7389 19805 7423 19839
rect 12173 19805 12207 19839
rect 12265 19805 12299 19839
rect 12449 19805 12483 19839
rect 12633 19805 12667 19839
rect 14105 19805 14139 19839
rect 14565 19805 14599 19839
rect 14933 19805 14967 19839
rect 15117 19805 15151 19839
rect 16313 19805 16347 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 17049 19805 17083 19839
rect 17785 19805 17819 19839
rect 17877 19805 17911 19839
rect 18245 19805 18279 19839
rect 18705 19805 18739 19839
rect 18889 19805 18923 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19809 19805 19843 19839
rect 19947 19805 19981 19839
rect 20453 19805 20487 19839
rect 21465 19805 21499 19839
rect 21649 19805 21683 19839
rect 24593 19805 24627 19839
rect 24961 19805 24995 19839
rect 25329 19805 25363 19839
rect 25605 19805 25639 19839
rect 26249 19805 26283 19839
rect 26525 19805 26559 19839
rect 26617 19805 26651 19839
rect 27169 19805 27203 19839
rect 27721 19805 27755 19839
rect 27985 19805 28019 19839
rect 28089 19805 28123 19839
rect 28457 19805 28491 19839
rect 28641 19805 28675 19839
rect 6193 19737 6227 19771
rect 7656 19737 7690 19771
rect 10048 19737 10082 19771
rect 15209 19737 15243 19771
rect 22293 19737 22327 19771
rect 23029 19737 23063 19771
rect 24777 19737 24811 19771
rect 24869 19737 24903 19771
rect 26433 19737 26467 19771
rect 26893 19737 26927 19771
rect 27445 19737 27479 19771
rect 11989 19669 12023 19703
rect 21833 19669 21867 19703
rect 23489 19669 23523 19703
rect 25145 19669 25179 19703
rect 26801 19669 26835 19703
rect 28365 19669 28399 19703
rect 28825 19669 28859 19703
rect 3249 19465 3283 19499
rect 3709 19465 3743 19499
rect 4261 19465 4295 19499
rect 6929 19465 6963 19499
rect 7297 19465 7331 19499
rect 8493 19465 8527 19499
rect 9413 19465 9447 19499
rect 9505 19465 9539 19499
rect 9597 19465 9631 19499
rect 10701 19465 10735 19499
rect 11345 19465 11379 19499
rect 12633 19465 12667 19499
rect 16773 19465 16807 19499
rect 23121 19465 23155 19499
rect 24501 19465 24535 19499
rect 25421 19465 25455 19499
rect 28641 19465 28675 19499
rect 1777 19397 1811 19431
rect 2114 19397 2148 19431
rect 8861 19397 8895 19431
rect 11621 19397 11655 19431
rect 12909 19397 12943 19431
rect 13001 19397 13035 19431
rect 14105 19397 14139 19431
rect 15577 19397 15611 19431
rect 20821 19397 20855 19431
rect 21281 19397 21315 19431
rect 23397 19397 23431 19431
rect 24133 19397 24167 19431
rect 24225 19397 24259 19431
rect 25053 19397 25087 19431
rect 27261 19397 27295 19431
rect 27353 19397 27387 19431
rect 27721 19397 27755 19431
rect 1593 19329 1627 19363
rect 3801 19329 3835 19363
rect 4445 19329 4479 19363
rect 4629 19329 4663 19363
rect 4997 19329 5031 19363
rect 5457 19329 5491 19363
rect 5733 19329 5767 19363
rect 5917 19329 5951 19363
rect 6101 19329 6135 19363
rect 6193 19329 6227 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 7113 19329 7147 19363
rect 7297 19329 7331 19363
rect 8585 19329 8619 19363
rect 8769 19329 8803 19363
rect 8953 19329 8987 19363
rect 9091 19329 9125 19363
rect 9321 19329 9355 19363
rect 9689 19329 9723 19363
rect 11989 19329 12023 19363
rect 12357 19329 12391 19363
rect 12541 19329 12575 19363
rect 12817 19329 12851 19363
rect 13119 19329 13153 19363
rect 13277 19329 13311 19363
rect 13645 19329 13679 19363
rect 13829 19329 13863 19363
rect 14841 19329 14875 19363
rect 15301 19329 15335 19363
rect 15485 19329 15519 19363
rect 16681 19329 16715 19363
rect 17325 19329 17359 19363
rect 17417 19329 17451 19363
rect 17693 19329 17727 19363
rect 18337 19329 18371 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19717 19329 19751 19363
rect 19993 19329 20027 19363
rect 20177 19329 20211 19363
rect 20545 19329 20579 19363
rect 20729 19329 20763 19363
rect 21097 19329 21131 19363
rect 21833 19329 21867 19363
rect 22569 19329 22603 19363
rect 23305 19329 23339 19363
rect 23489 19329 23523 19363
rect 23673 19329 23707 19363
rect 23765 19329 23799 19363
rect 23857 19329 23891 19363
rect 23950 19329 23984 19363
rect 24361 19329 24395 19363
rect 24869 19329 24903 19363
rect 25145 19329 25179 19363
rect 25237 19329 25271 19363
rect 26525 19329 26559 19363
rect 26974 19329 27008 19363
rect 27078 19329 27112 19363
rect 27450 19329 27484 19363
rect 27997 19329 28031 19363
rect 28273 19329 28307 19363
rect 28457 19329 28491 19363
rect 1409 19261 1443 19295
rect 1869 19261 1903 19295
rect 3893 19261 3927 19295
rect 4169 19261 4203 19295
rect 4905 19261 4939 19295
rect 5549 19261 5583 19295
rect 5641 19261 5675 19295
rect 7941 19261 7975 19295
rect 9229 19261 9263 19295
rect 10057 19261 10091 19295
rect 11529 19261 11563 19295
rect 11897 19261 11931 19295
rect 15393 19261 15427 19295
rect 16313 19261 16347 19295
rect 17601 19261 17635 19295
rect 18429 19261 18463 19295
rect 19257 19261 19291 19295
rect 19625 19261 19659 19295
rect 20269 19261 20303 19295
rect 25973 19261 26007 19295
rect 27813 19261 27847 19295
rect 13921 19193 13955 19227
rect 18153 19193 18187 19227
rect 21465 19193 21499 19227
rect 27629 19193 27663 19227
rect 3341 19125 3375 19159
rect 5273 19125 5307 19159
rect 5917 19125 5951 19159
rect 6469 19125 6503 19159
rect 7757 19125 7791 19159
rect 17141 19125 17175 19159
rect 19901 19125 19935 19159
rect 27721 19125 27755 19159
rect 28181 19125 28215 19159
rect 3525 18921 3559 18955
rect 5365 18921 5399 18955
rect 6745 18921 6779 18955
rect 8401 18921 8435 18955
rect 9505 18921 9539 18955
rect 10057 18921 10091 18955
rect 11621 18921 11655 18955
rect 15485 18921 15519 18955
rect 15945 18921 15979 18955
rect 21005 18921 21039 18955
rect 21097 18921 21131 18955
rect 21833 18921 21867 18955
rect 22201 18921 22235 18955
rect 23121 18921 23155 18955
rect 24041 18921 24075 18955
rect 24225 18921 24259 18955
rect 24593 18921 24627 18955
rect 25145 18921 25179 18955
rect 26525 18921 26559 18955
rect 29101 18921 29135 18955
rect 12725 18853 12759 18887
rect 13185 18853 13219 18887
rect 14381 18853 14415 18887
rect 17509 18853 17543 18887
rect 19717 18853 19751 18887
rect 22293 18853 22327 18887
rect 23029 18853 23063 18887
rect 3801 18785 3835 18819
rect 5917 18785 5951 18819
rect 10701 18785 10735 18819
rect 11253 18785 11287 18819
rect 18981 18785 19015 18819
rect 20269 18785 20303 18819
rect 22661 18785 22695 18819
rect 1593 18717 1627 18751
rect 2973 18717 3007 18751
rect 5641 18717 5675 18751
rect 6101 18717 6135 18751
rect 6194 18717 6228 18751
rect 6469 18717 6503 18751
rect 6566 18717 6600 18751
rect 6837 18717 6871 18751
rect 7021 18717 7055 18751
rect 10241 18717 10275 18751
rect 10333 18717 10367 18751
rect 11529 18717 11563 18751
rect 12173 18717 12207 18751
rect 12357 18717 12391 18751
rect 12817 18717 12851 18751
rect 13369 18717 13403 18751
rect 13737 18717 13771 18751
rect 13921 18717 13955 18751
rect 14197 18717 14231 18751
rect 15025 18717 15059 18751
rect 15761 18717 15795 18751
rect 16037 18717 16071 18751
rect 16405 18717 16439 18751
rect 16865 18717 16899 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 17877 18717 17911 18751
rect 18153 18717 18187 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 19441 18717 19475 18751
rect 19717 18717 19751 18751
rect 20361 18717 20395 18751
rect 21281 18717 21315 18751
rect 21373 18717 21407 18751
rect 21465 18717 21499 18751
rect 21741 18717 21775 18751
rect 22109 18717 22143 18751
rect 22569 18717 22603 18751
rect 22845 18717 22879 18751
rect 23305 18717 23339 18751
rect 23489 18717 23523 18751
rect 23627 18717 23661 18751
rect 23765 18717 23799 18751
rect 24409 18717 24443 18751
rect 25329 18717 25363 18751
rect 25513 18717 25547 18751
rect 25631 18717 25665 18751
rect 25789 18717 25823 18751
rect 25881 18717 25915 18751
rect 25974 18717 26008 18751
rect 26249 18717 26283 18751
rect 26346 18717 26380 18751
rect 26617 18717 26651 18751
rect 26710 18717 26744 18751
rect 27082 18717 27116 18751
rect 27721 18717 27755 18751
rect 27988 18717 28022 18751
rect 2329 18649 2363 18683
rect 4068 18649 4102 18683
rect 6377 18649 6411 18683
rect 7941 18649 7975 18683
rect 8769 18649 8803 18683
rect 10425 18649 10459 18683
rect 10543 18649 10577 18683
rect 11345 18649 11379 18683
rect 13645 18649 13679 18683
rect 18429 18649 18463 18683
rect 19901 18649 19935 18683
rect 20085 18649 20119 18683
rect 21603 18649 21637 18683
rect 23397 18649 23431 18683
rect 23857 18649 23891 18683
rect 25421 18649 25455 18683
rect 26157 18649 26191 18683
rect 26893 18649 26927 18683
rect 26985 18649 27019 18683
rect 5181 18581 5215 18615
rect 5825 18581 5859 18615
rect 6929 18581 6963 18615
rect 7665 18581 7699 18615
rect 9137 18581 9171 18615
rect 9965 18581 9999 18615
rect 12357 18581 12391 18615
rect 12909 18581 12943 18615
rect 13553 18581 13587 18615
rect 13829 18581 13863 18615
rect 15577 18581 15611 18615
rect 22477 18581 22511 18615
rect 24057 18581 24091 18615
rect 24869 18581 24903 18615
rect 27261 18581 27295 18615
rect 3065 18377 3099 18411
rect 3525 18377 3559 18411
rect 3617 18377 3651 18411
rect 4905 18377 4939 18411
rect 5733 18377 5767 18411
rect 7119 18377 7153 18411
rect 7849 18377 7883 18411
rect 7941 18377 7975 18411
rect 8585 18377 8619 18411
rect 10977 18377 11011 18411
rect 11345 18377 11379 18411
rect 13185 18377 13219 18411
rect 13737 18377 13771 18411
rect 16497 18377 16531 18411
rect 16957 18377 16991 18411
rect 18705 18377 18739 18411
rect 20913 18377 20947 18411
rect 21097 18377 21131 18411
rect 23857 18377 23891 18411
rect 24685 18377 24719 18411
rect 25329 18377 25363 18411
rect 26341 18377 26375 18411
rect 7021 18309 7055 18343
rect 7205 18309 7239 18343
rect 8861 18309 8895 18343
rect 9781 18309 9815 18343
rect 11989 18309 12023 18343
rect 12127 18309 12161 18343
rect 22109 18309 22143 18343
rect 22661 18309 22695 18343
rect 23397 18309 23431 18343
rect 24317 18309 24351 18343
rect 27252 18309 27286 18343
rect 1685 18241 1719 18275
rect 1952 18241 1986 18275
rect 5089 18241 5123 18275
rect 5825 18241 5859 18275
rect 6009 18241 6043 18275
rect 6745 18241 6779 18275
rect 7297 18241 7331 18275
rect 7389 18241 7423 18275
rect 7573 18241 7607 18275
rect 7757 18241 7791 18275
rect 8405 18241 8439 18275
rect 8493 18241 8527 18275
rect 9045 18241 9079 18275
rect 9137 18241 9171 18275
rect 9229 18241 9263 18275
rect 9413 18241 9447 18275
rect 9965 18241 9999 18275
rect 10057 18241 10091 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 11805 18241 11839 18275
rect 11897 18241 11931 18275
rect 12541 18241 12575 18275
rect 13001 18241 13035 18275
rect 13277 18241 13311 18275
rect 13553 18241 13587 18275
rect 13829 18241 13863 18275
rect 13921 18241 13955 18275
rect 14105 18241 14139 18275
rect 14197 18241 14231 18275
rect 14381 18241 14415 18275
rect 14473 18241 14507 18275
rect 14565 18241 14599 18275
rect 14749 18241 14783 18275
rect 14841 18241 14875 18275
rect 14933 18241 14967 18275
rect 15301 18241 15335 18275
rect 15577 18241 15611 18275
rect 16129 18241 16163 18275
rect 16313 18241 16347 18275
rect 16957 18241 16991 18275
rect 17141 18241 17175 18275
rect 17325 18241 17359 18275
rect 17601 18241 17635 18275
rect 17877 18241 17911 18275
rect 17969 18241 18003 18275
rect 18889 18241 18923 18275
rect 19165 18241 19199 18275
rect 19901 18241 19935 18275
rect 20821 18241 20855 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 21373 18241 21407 18275
rect 21557 18241 21591 18275
rect 21649 18241 21683 18275
rect 22201 18241 22235 18275
rect 22845 18241 22879 18275
rect 24133 18241 24167 18275
rect 24409 18241 24443 18275
rect 24501 18241 24535 18275
rect 24777 18241 24811 18275
rect 24961 18241 24995 18275
rect 25053 18241 25087 18275
rect 25145 18241 25179 18275
rect 25513 18241 25547 18275
rect 26525 18241 26559 18275
rect 3801 18173 3835 18207
rect 4353 18173 4387 18207
rect 6377 18173 6411 18207
rect 6561 18173 6595 18207
rect 6653 18173 6687 18207
rect 6837 18173 6871 18207
rect 8125 18173 8159 18207
rect 8769 18173 8803 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 12633 18173 12667 18207
rect 12725 18173 12759 18207
rect 12817 18173 12851 18207
rect 15761 18173 15795 18207
rect 18429 18173 18463 18207
rect 19349 18173 19383 18207
rect 20453 18173 20487 18207
rect 22753 18173 22787 18207
rect 23305 18173 23339 18207
rect 26801 18173 26835 18207
rect 26985 18173 27019 18207
rect 8677 18105 8711 18139
rect 8861 18105 8895 18139
rect 9781 18105 9815 18139
rect 15393 18105 15427 18139
rect 17601 18105 17635 18139
rect 18981 18105 19015 18139
rect 23765 18105 23799 18139
rect 26709 18105 26743 18139
rect 3157 18037 3191 18071
rect 6193 18037 6227 18071
rect 7481 18037 7515 18071
rect 7849 18037 7883 18071
rect 9321 18037 9355 18071
rect 10241 18037 10275 18071
rect 11621 18037 11655 18071
rect 13001 18037 13035 18071
rect 13369 18037 13403 18071
rect 15117 18037 15151 18071
rect 18337 18037 18371 18071
rect 21925 18037 21959 18071
rect 26065 18037 26099 18071
rect 28365 18037 28399 18071
rect 3617 17833 3651 17867
rect 4353 17833 4387 17867
rect 7113 17833 7147 17867
rect 8677 17833 8711 17867
rect 11069 17833 11103 17867
rect 13921 17833 13955 17867
rect 14197 17833 14231 17867
rect 17233 17833 17267 17867
rect 18521 17833 18555 17867
rect 20637 17833 20671 17867
rect 21189 17833 21223 17867
rect 22569 17833 22603 17867
rect 23121 17833 23155 17867
rect 25421 17833 25455 17867
rect 25881 17833 25915 17867
rect 26801 17833 26835 17867
rect 8953 17765 8987 17799
rect 17601 17765 17635 17799
rect 18705 17765 18739 17799
rect 21649 17765 21683 17799
rect 21925 17765 21959 17799
rect 22109 17765 22143 17799
rect 23489 17765 23523 17799
rect 24041 17765 24075 17799
rect 1869 17697 1903 17731
rect 2973 17697 3007 17731
rect 5089 17697 5123 17731
rect 6193 17697 6227 17731
rect 7297 17697 7331 17731
rect 7389 17697 7423 17731
rect 7481 17697 7515 17731
rect 7573 17697 7607 17731
rect 9229 17697 9263 17731
rect 9321 17697 9355 17731
rect 9413 17697 9447 17731
rect 10517 17697 10551 17731
rect 11345 17697 11379 17731
rect 11713 17697 11747 17731
rect 16037 17697 16071 17731
rect 16405 17697 16439 17731
rect 18061 17697 18095 17731
rect 18613 17697 18647 17731
rect 19257 17697 19291 17731
rect 21373 17697 21407 17731
rect 25053 17697 25087 17731
rect 1593 17629 1627 17663
rect 4077 17629 4111 17663
rect 4261 17629 4295 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 4997 17629 5031 17663
rect 5825 17629 5859 17663
rect 5917 17629 5951 17663
rect 6377 17629 6411 17663
rect 7849 17629 7883 17663
rect 8585 17629 8619 17663
rect 8769 17629 8803 17663
rect 9137 17629 9171 17663
rect 9781 17629 9815 17663
rect 9965 17629 9999 17663
rect 10241 17629 10275 17663
rect 10609 17629 10643 17663
rect 10701 17629 10735 17663
rect 10793 17629 10827 17663
rect 10977 17629 11011 17663
rect 12725 17629 12759 17663
rect 13553 17629 13587 17663
rect 14105 17629 14139 17663
rect 14565 17629 14599 17663
rect 14887 17629 14921 17663
rect 15025 17629 15059 17663
rect 15117 17629 15151 17663
rect 15393 17629 15427 17663
rect 15577 17629 15611 17663
rect 16129 17629 16163 17663
rect 16773 17629 16807 17663
rect 16865 17629 16899 17663
rect 16957 17629 16991 17663
rect 17049 17629 17083 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 18153 17629 18187 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 19717 17629 19751 17663
rect 19901 17629 19935 17663
rect 20085 17629 20119 17663
rect 20545 17629 20579 17663
rect 20821 17629 20855 17663
rect 21097 17629 21131 17663
rect 21189 17629 21223 17663
rect 21465 17629 21499 17663
rect 21833 17629 21867 17663
rect 22293 17629 22327 17663
rect 22385 17629 22419 17663
rect 23305 17629 23339 17663
rect 23581 17629 23615 17663
rect 24593 17629 24627 17663
rect 26157 17629 26191 17663
rect 26433 17629 26467 17663
rect 4169 17561 4203 17595
rect 4629 17561 4663 17595
rect 4839 17561 4873 17595
rect 5733 17561 5767 17595
rect 9873 17561 9907 17595
rect 10103 17561 10137 17595
rect 13369 17561 13403 17595
rect 13645 17561 13679 17595
rect 13737 17561 13771 17595
rect 14381 17561 14415 17595
rect 14657 17561 14691 17595
rect 14749 17561 14783 17595
rect 16497 17561 16531 17595
rect 20269 17561 20303 17595
rect 23673 17561 23707 17595
rect 24685 17561 24719 17595
rect 24777 17561 24811 17595
rect 24895 17561 24929 17595
rect 25513 17561 25547 17595
rect 25697 17561 25731 17595
rect 25973 17561 26007 17595
rect 26341 17561 26375 17595
rect 26617 17561 26651 17595
rect 6009 17493 6043 17527
rect 6101 17493 6135 17527
rect 6929 17493 6963 17527
rect 8493 17493 8527 17527
rect 9597 17493 9631 17527
rect 10333 17493 10367 17527
rect 11069 17493 11103 17527
rect 11161 17493 11195 17527
rect 12357 17493 12391 17527
rect 13277 17493 13311 17527
rect 15209 17493 15243 17527
rect 15853 17493 15887 17527
rect 16589 17493 16623 17527
rect 21005 17493 21039 17527
rect 24133 17493 24167 17527
rect 24409 17493 24443 17527
rect 1685 17289 1719 17323
rect 3617 17289 3651 17323
rect 5089 17289 5123 17323
rect 6377 17289 6411 17323
rect 7757 17289 7791 17323
rect 7849 17289 7883 17323
rect 10885 17289 10919 17323
rect 12909 17289 12943 17323
rect 13093 17289 13127 17323
rect 13185 17289 13219 17323
rect 13461 17289 13495 17323
rect 20637 17289 20671 17323
rect 21281 17289 21315 17323
rect 21649 17289 21683 17323
rect 22477 17289 22511 17323
rect 22845 17289 22879 17323
rect 24501 17289 24535 17323
rect 43269 17289 43303 17323
rect 5457 17221 5491 17255
rect 5549 17221 5583 17255
rect 5667 17221 5701 17255
rect 5917 17221 5951 17255
rect 6653 17221 6687 17255
rect 8125 17221 8159 17255
rect 9965 17221 9999 17255
rect 11796 17221 11830 17255
rect 19717 17221 19751 17255
rect 21373 17221 21407 17255
rect 22017 17221 22051 17255
rect 24041 17221 24075 17255
rect 2044 17153 2078 17187
rect 3433 17153 3467 17187
rect 3709 17153 3743 17187
rect 3976 17153 4010 17187
rect 5365 17153 5399 17187
rect 6101 17153 6135 17187
rect 6193 17153 6227 17187
rect 6561 17153 6595 17187
rect 6745 17153 6779 17187
rect 6863 17153 6897 17187
rect 7205 17153 7239 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 8335 17153 8369 17187
rect 8677 17153 8711 17187
rect 9413 17153 9447 17187
rect 10057 17153 10091 17187
rect 10793 17153 10827 17187
rect 10977 17153 11011 17187
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 13369 17153 13403 17187
rect 13645 17153 13679 17187
rect 13921 17153 13955 17187
rect 14197 17153 14231 17187
rect 15577 17153 15611 17187
rect 15761 17153 15795 17187
rect 16037 17153 16071 17187
rect 17049 17153 17083 17187
rect 17141 17153 17175 17187
rect 17509 17153 17543 17187
rect 17785 17153 17819 17187
rect 17877 17153 17911 17187
rect 18429 17153 18463 17187
rect 19073 17153 19107 17187
rect 19257 17153 19291 17187
rect 19625 17153 19659 17187
rect 19809 17153 19843 17187
rect 19993 17153 20027 17187
rect 20085 17153 20119 17187
rect 20453 17153 20487 17187
rect 21005 17153 21039 17187
rect 22753 17153 22787 17187
rect 23029 17153 23063 17187
rect 23121 17153 23155 17187
rect 23397 17153 23431 17187
rect 23581 17153 23615 17187
rect 43177 17153 43211 17187
rect 1777 17085 1811 17119
rect 3249 17085 3283 17119
rect 5825 17085 5859 17119
rect 7021 17085 7055 17119
rect 8493 17085 8527 17119
rect 9229 17085 9263 17119
rect 11529 17085 11563 17119
rect 14933 17085 14967 17119
rect 17233 17085 17267 17119
rect 21490 17085 21524 17119
rect 22569 17085 22603 17119
rect 23857 17085 23891 17119
rect 16221 17017 16255 17051
rect 22017 17017 22051 17051
rect 24409 17017 24443 17051
rect 3157 16949 3191 16983
rect 5181 16949 5215 16983
rect 5917 16949 5951 16983
rect 10701 16949 10735 16983
rect 13093 16949 13127 16983
rect 13829 16949 13863 16983
rect 14749 16949 14783 16983
rect 15485 16949 15519 16983
rect 15669 16949 15703 16983
rect 19441 16949 19475 16983
rect 20453 16949 20487 16983
rect 23305 16949 23339 16983
rect 4169 16745 4203 16779
rect 4905 16745 4939 16779
rect 8769 16745 8803 16779
rect 9045 16745 9079 16779
rect 13093 16745 13127 16779
rect 14197 16745 14231 16779
rect 16313 16745 16347 16779
rect 17417 16745 17451 16779
rect 17509 16745 17543 16779
rect 18521 16745 18555 16779
rect 18889 16745 18923 16779
rect 19625 16745 19659 16779
rect 19993 16745 20027 16779
rect 2881 16677 2915 16711
rect 7297 16677 7331 16711
rect 10977 16677 11011 16711
rect 15761 16677 15795 16711
rect 17141 16677 17175 16711
rect 3525 16609 3559 16643
rect 3801 16609 3835 16643
rect 4353 16609 4387 16643
rect 5917 16609 5951 16643
rect 9321 16609 9355 16643
rect 12357 16609 12391 16643
rect 13277 16609 13311 16643
rect 16681 16609 16715 16643
rect 17601 16609 17635 16643
rect 18613 16609 18647 16643
rect 20545 16609 20579 16643
rect 21557 16609 21591 16643
rect 21925 16609 21959 16643
rect 22661 16609 22695 16643
rect 1593 16541 1627 16575
rect 3249 16541 3283 16575
rect 3341 16541 3375 16575
rect 3985 16541 4019 16575
rect 4997 16541 5031 16575
rect 6184 16541 6218 16575
rect 7389 16541 7423 16575
rect 7656 16541 7690 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9588 16541 9622 16575
rect 11345 16541 11379 16575
rect 11529 16541 11563 16575
rect 11621 16541 11655 16575
rect 11897 16541 11931 16575
rect 12173 16541 12207 16575
rect 13020 16519 13054 16553
rect 13645 16541 13679 16575
rect 13829 16541 13863 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 14648 16541 14682 16575
rect 15853 16541 15887 16575
rect 17325 16541 17359 16575
rect 18061 16541 18095 16575
rect 18153 16541 18187 16575
rect 19257 16541 19291 16575
rect 19625 16541 19659 16575
rect 19901 16541 19935 16575
rect 19993 16541 20027 16575
rect 20177 16541 20211 16575
rect 20453 16541 20487 16575
rect 20637 16541 20671 16575
rect 20729 16541 20763 16575
rect 22109 16541 22143 16575
rect 22477 16541 22511 16575
rect 23029 16541 23063 16575
rect 2329 16473 2363 16507
rect 13277 16473 13311 16507
rect 13461 16473 13495 16507
rect 13921 16473 13955 16507
rect 21649 16473 21683 16507
rect 23305 16473 23339 16507
rect 5641 16405 5675 16439
rect 10701 16405 10735 16439
rect 11161 16405 11195 16439
rect 11713 16405 11747 16439
rect 12081 16405 12115 16439
rect 12909 16405 12943 16439
rect 16037 16405 16071 16439
rect 19441 16405 19475 16439
rect 20821 16405 20855 16439
rect 22017 16405 22051 16439
rect 22293 16405 22327 16439
rect 3433 16201 3467 16235
rect 4629 16201 4663 16235
rect 6101 16201 6135 16235
rect 7481 16201 7515 16235
rect 8217 16201 8251 16235
rect 9781 16201 9815 16235
rect 10149 16201 10183 16235
rect 10793 16201 10827 16235
rect 11897 16201 11931 16235
rect 15853 16201 15887 16235
rect 16129 16201 16163 16235
rect 16865 16201 16899 16235
rect 19533 16201 19567 16235
rect 23213 16201 23247 16235
rect 1961 16133 1995 16167
rect 2298 16133 2332 16167
rect 3893 16133 3927 16167
rect 7021 16133 7055 16167
rect 12633 16133 12667 16167
rect 13829 16133 13863 16167
rect 14740 16133 14774 16167
rect 1685 16065 1719 16099
rect 1777 16065 1811 16099
rect 2053 16065 2087 16099
rect 4997 16065 5031 16099
rect 5549 16065 5583 16099
rect 6469 16065 6503 16099
rect 7297 16065 7331 16099
rect 7573 16065 7607 16099
rect 8033 16065 8067 16099
rect 8309 16065 8343 16099
rect 9597 16065 9631 16099
rect 9873 16065 9907 16099
rect 13645 16065 13679 16099
rect 14473 16065 14507 16099
rect 17417 16065 17451 16099
rect 18981 16065 19015 16099
rect 19257 16065 19291 16099
rect 20536 16065 20570 16099
rect 22100 16065 22134 16099
rect 3985 15997 4019 16031
rect 4077 15997 4111 16031
rect 5089 15997 5123 16031
rect 5181 15997 5215 16031
rect 8769 15997 8803 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 13001 15997 13035 16031
rect 17233 15997 17267 16031
rect 20269 15997 20303 16031
rect 21833 15997 21867 16031
rect 11253 15929 11287 15963
rect 21649 15929 21683 15963
rect 3525 15861 3559 15895
rect 7113 15861 7147 15895
rect 7849 15861 7883 15895
rect 9321 15861 9355 15895
rect 9413 15861 9447 15895
rect 11529 15861 11563 15895
rect 13921 15861 13955 15895
rect 17601 15861 17635 15895
rect 17969 15861 18003 15895
rect 19257 15861 19291 15895
rect 3617 15657 3651 15691
rect 7481 15657 7515 15691
rect 8585 15657 8619 15691
rect 8953 15657 8987 15691
rect 12449 15657 12483 15691
rect 22753 15657 22787 15691
rect 16037 15589 16071 15623
rect 16313 15589 16347 15623
rect 18521 15589 18555 15623
rect 1869 15521 1903 15555
rect 3065 15521 3099 15555
rect 6285 15521 6319 15555
rect 8033 15521 8067 15555
rect 9505 15521 9539 15555
rect 9873 15521 9907 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14657 15521 14691 15555
rect 14933 15521 14967 15555
rect 17141 15521 17175 15555
rect 21373 15521 21407 15555
rect 1593 15453 1627 15487
rect 3893 15453 3927 15487
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 6101 15453 6135 15487
rect 6561 15453 6595 15487
rect 10609 15453 10643 15487
rect 10793 15453 10827 15487
rect 11069 15453 11103 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 14473 15453 14507 15487
rect 15577 15453 15611 15487
rect 17408 15453 17442 15487
rect 21640 15453 21674 15487
rect 4169 15385 4203 15419
rect 4506 15385 4540 15419
rect 7205 15385 7239 15419
rect 9321 15385 9355 15419
rect 10425 15385 10459 15419
rect 10977 15385 11011 15419
rect 11314 15385 11348 15419
rect 13001 15385 13035 15419
rect 5641 15317 5675 15351
rect 5733 15317 5767 15351
rect 6193 15317 6227 15351
rect 9413 15317 9447 15351
rect 12541 15317 12575 15351
rect 13737 15317 13771 15351
rect 14105 15317 14139 15351
rect 14565 15317 14599 15351
rect 1685 15113 1719 15147
rect 2881 15113 2915 15147
rect 3617 15113 3651 15147
rect 3985 15113 4019 15147
rect 5457 15113 5491 15147
rect 7665 15113 7699 15147
rect 8493 15113 8527 15147
rect 9965 15113 9999 15147
rect 10425 15113 10459 15147
rect 12909 15113 12943 15147
rect 14565 15113 14599 15147
rect 15025 15113 15059 15147
rect 5917 15045 5951 15079
rect 6745 15045 6779 15079
rect 8830 15045 8864 15079
rect 3065 14977 3099 15011
rect 4077 14977 4111 15011
rect 4344 14977 4378 15011
rect 5733 14977 5767 15011
rect 6009 14977 6043 15011
rect 7021 14977 7055 15011
rect 8125 14977 8159 15011
rect 8309 14977 8343 15011
rect 8585 14977 8619 15011
rect 11161 14977 11195 15011
rect 11529 14977 11563 15011
rect 11796 14977 11830 15011
rect 13185 14977 13219 15011
rect 13452 14977 13486 15011
rect 2329 14909 2363 14943
rect 6837 14909 6871 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 10977 14909 11011 14943
rect 7297 14841 7331 14875
rect 2145 14773 2179 14807
rect 5549 14773 5583 14807
rect 7205 14773 7239 14807
rect 10885 14773 10919 14807
rect 11345 14773 11379 14807
rect 3249 14569 3283 14603
rect 3525 14569 3559 14603
rect 4169 14569 4203 14603
rect 6653 14569 6687 14603
rect 8125 14569 8159 14603
rect 8493 14569 8527 14603
rect 9229 14569 9263 14603
rect 11529 14569 11563 14603
rect 13921 14569 13955 14603
rect 14289 14569 14323 14603
rect 4537 14501 4571 14535
rect 9873 14501 9907 14535
rect 13369 14501 13403 14535
rect 1869 14433 1903 14467
rect 3801 14433 3835 14467
rect 4997 14433 5031 14467
rect 6745 14433 6779 14467
rect 1593 14365 1627 14399
rect 3985 14365 4019 14399
rect 5273 14365 5307 14399
rect 7012 14365 7046 14399
rect 5540 14297 5574 14331
rect 2053 14025 2087 14059
rect 5181 14025 5215 14059
rect 6193 14025 6227 14059
rect 6377 14025 6411 14059
rect 6837 14025 6871 14059
rect 7849 14025 7883 14059
rect 8125 14025 8159 14059
rect 8953 14025 8987 14059
rect 3341 13957 3375 13991
rect 4077 13957 4111 13991
rect 4445 13957 4479 13991
rect 4905 13957 4939 13991
rect 3801 13889 3835 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 6009 13889 6043 13923
rect 6745 13889 6779 13923
rect 7205 13889 7239 13923
rect 6929 13821 6963 13855
rect 8585 13753 8619 13787
rect 3617 13481 3651 13515
rect 4261 13481 4295 13515
rect 4629 13481 4663 13515
rect 5181 13481 5215 13515
rect 6009 13481 6043 13515
rect 6377 13481 6411 13515
rect 6929 13481 6963 13515
rect 7481 13481 7515 13515
rect 5549 13413 5583 13447
rect 8125 13413 8159 13447
rect 1869 13345 1903 13379
rect 7849 13345 7883 13379
rect 1593 13277 1627 13311
rect 4261 12937 4295 12971
rect 5917 12937 5951 12971
rect 6653 12937 6687 12971
rect 7665 12869 7699 12903
rect 6929 12801 6963 12835
rect 7297 12801 7331 12835
rect 1869 12257 1903 12291
rect 1593 12189 1627 12223
rect 1869 11169 1903 11203
rect 1593 11101 1627 11135
rect 1869 10081 1903 10115
rect 1593 10013 1627 10047
rect 1869 8993 1903 9027
rect 1593 8925 1627 8959
rect 1869 7905 1903 7939
rect 1593 7837 1627 7871
rect 1869 6817 1903 6851
rect 1593 6749 1627 6783
rect 1869 5729 1903 5763
rect 1593 5661 1627 5695
rect 3157 5525 3191 5559
rect 3157 4777 3191 4811
rect 1869 4641 1903 4675
rect 1593 4573 1627 4607
rect 3157 3689 3191 3723
rect 1869 3553 1903 3587
rect 1593 3485 1627 3519
rect 24685 2601 24719 2635
rect 23029 2465 23063 2499
rect 22753 2397 22787 2431
<< metal1 >>
rect 1104 42458 43884 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 43884 42458
rect 1104 42384 43884 42406
rect 24210 42304 24216 42356
rect 24268 42304 24274 42356
rect 25406 42304 25412 42356
rect 25464 42304 25470 42356
rect 26602 42304 26608 42356
rect 26660 42304 26666 42356
rect 27798 42304 27804 42356
rect 27856 42304 27862 42356
rect 28994 42304 29000 42356
rect 29052 42304 29058 42356
rect 30190 42304 30196 42356
rect 30248 42344 30254 42356
rect 30248 42316 30512 42344
rect 30248 42304 30254 42316
rect 24228 42208 24256 42304
rect 24581 42211 24639 42217
rect 24581 42208 24593 42211
rect 24228 42180 24593 42208
rect 24581 42177 24593 42180
rect 24627 42177 24639 42211
rect 25424 42208 25452 42304
rect 25685 42211 25743 42217
rect 25685 42208 25697 42211
rect 25424 42180 25697 42208
rect 24581 42171 24639 42177
rect 25685 42177 25697 42180
rect 25731 42177 25743 42211
rect 26620 42208 26648 42304
rect 27157 42211 27215 42217
rect 27157 42208 27169 42211
rect 26620 42180 27169 42208
rect 25685 42171 25743 42177
rect 27157 42177 27169 42180
rect 27203 42177 27215 42211
rect 27816 42208 27844 42304
rect 28077 42211 28135 42217
rect 28077 42208 28089 42211
rect 27816 42180 28089 42208
rect 27157 42171 27215 42177
rect 28077 42177 28089 42180
rect 28123 42177 28135 42211
rect 29012 42208 29040 42304
rect 30484 42217 30512 42316
rect 31386 42304 31392 42356
rect 31444 42304 31450 42356
rect 32582 42304 32588 42356
rect 32640 42304 32646 42356
rect 36170 42304 36176 42356
rect 36228 42304 36234 42356
rect 37366 42304 37372 42356
rect 37424 42304 37430 42356
rect 29273 42211 29331 42217
rect 29273 42208 29285 42211
rect 29012 42180 29285 42208
rect 28077 42171 28135 42177
rect 29273 42177 29285 42180
rect 29319 42177 29331 42211
rect 29273 42171 29331 42177
rect 30469 42211 30527 42217
rect 30469 42177 30481 42211
rect 30515 42177 30527 42211
rect 31404 42208 31432 42304
rect 31665 42211 31723 42217
rect 31665 42208 31677 42211
rect 31404 42180 31677 42208
rect 30469 42171 30527 42177
rect 31665 42177 31677 42180
rect 31711 42177 31723 42211
rect 32600 42208 32628 42304
rect 34974 42236 34980 42288
rect 35032 42276 35038 42288
rect 35161 42279 35219 42285
rect 35161 42276 35173 42279
rect 35032 42248 35173 42276
rect 35032 42236 35038 42248
rect 35161 42245 35173 42248
rect 35207 42245 35219 42279
rect 35161 42239 35219 42245
rect 32861 42211 32919 42217
rect 32861 42208 32873 42211
rect 32600 42180 32873 42208
rect 31665 42171 31723 42177
rect 32861 42177 32873 42180
rect 32907 42177 32919 42211
rect 36188 42208 36216 42304
rect 36265 42211 36323 42217
rect 36265 42208 36277 42211
rect 36188 42180 36277 42208
rect 32861 42171 32919 42177
rect 36265 42177 36277 42180
rect 36311 42177 36323 42211
rect 37384 42208 37412 42304
rect 37461 42211 37519 42217
rect 37461 42208 37473 42211
rect 37384 42180 37473 42208
rect 36265 42171 36323 42177
rect 37461 42177 37473 42180
rect 37507 42177 37519 42211
rect 37461 42171 37519 42177
rect 23934 42032 23940 42084
rect 23992 42072 23998 42084
rect 25501 42075 25559 42081
rect 25501 42072 25513 42075
rect 23992 42044 25513 42072
rect 23992 42032 23998 42044
rect 25501 42041 25513 42044
rect 25547 42041 25559 42075
rect 25501 42035 25559 42041
rect 24397 42007 24455 42013
rect 24397 41973 24409 42007
rect 24443 42004 24455 42007
rect 24486 42004 24492 42016
rect 24443 41976 24492 42004
rect 24443 41973 24455 41976
rect 24397 41967 24455 41973
rect 24486 41964 24492 41976
rect 24544 41964 24550 42016
rect 26973 42007 27031 42013
rect 26973 41973 26985 42007
rect 27019 42004 27031 42007
rect 27338 42004 27344 42016
rect 27019 41976 27344 42004
rect 27019 41973 27031 41976
rect 26973 41967 27031 41973
rect 27338 41964 27344 41976
rect 27396 41964 27402 42016
rect 27890 41964 27896 42016
rect 27948 41964 27954 42016
rect 29086 41964 29092 42016
rect 29144 41964 29150 42016
rect 30285 42007 30343 42013
rect 30285 41973 30297 42007
rect 30331 42004 30343 42007
rect 31018 42004 31024 42016
rect 30331 41976 31024 42004
rect 30331 41973 30343 41976
rect 30285 41967 30343 41973
rect 31018 41964 31024 41976
rect 31076 41964 31082 42016
rect 31478 41964 31484 42016
rect 31536 41964 31542 42016
rect 32674 41964 32680 42016
rect 32732 41964 32738 42016
rect 32766 41964 32772 42016
rect 32824 42004 32830 42016
rect 35253 42007 35311 42013
rect 35253 42004 35265 42007
rect 32824 41976 35265 42004
rect 32824 41964 32830 41976
rect 35253 41973 35265 41976
rect 35299 41973 35311 42007
rect 35253 41967 35311 41973
rect 36446 41964 36452 42016
rect 36504 41964 36510 42016
rect 37642 41964 37648 42016
rect 37700 41964 37706 42016
rect 1104 41914 43884 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 43884 41914
rect 1104 41840 43884 41862
rect 17678 41760 17684 41812
rect 17736 41800 17742 41812
rect 32766 41800 32772 41812
rect 17736 41772 32772 41800
rect 17736 41760 17742 41772
rect 32766 41760 32772 41772
rect 32824 41760 32830 41812
rect 934 41556 940 41608
rect 992 41596 998 41608
rect 1581 41599 1639 41605
rect 1581 41596 1593 41599
rect 992 41568 1593 41596
rect 992 41556 998 41568
rect 1581 41565 1593 41568
rect 1627 41565 1639 41599
rect 1581 41559 1639 41565
rect 28718 41488 28724 41540
rect 28776 41528 28782 41540
rect 29273 41531 29331 41537
rect 29273 41528 29285 41531
rect 28776 41500 29285 41528
rect 28776 41488 28782 41500
rect 29273 41497 29285 41500
rect 29319 41497 29331 41531
rect 29273 41491 29331 41497
rect 28997 41463 29055 41469
rect 28997 41429 29009 41463
rect 29043 41460 29055 41463
rect 29178 41460 29184 41472
rect 29043 41432 29184 41460
rect 29043 41429 29055 41432
rect 28997 41423 29055 41429
rect 29178 41420 29184 41432
rect 29236 41420 29242 41472
rect 1104 41370 43884 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 43884 41370
rect 1104 41296 43884 41318
rect 28810 41216 28816 41268
rect 28868 41256 28874 41268
rect 29638 41256 29644 41268
rect 28868 41228 29644 41256
rect 28868 41216 28874 41228
rect 29638 41216 29644 41228
rect 29696 41216 29702 41268
rect 28368 41160 28994 41188
rect 28368 41132 28396 41160
rect 28350 41080 28356 41132
rect 28408 41080 28414 41132
rect 28966 41120 28994 41160
rect 28966 41092 29040 41120
rect 8110 41012 8116 41064
rect 8168 41012 8174 41064
rect 9122 41012 9128 41064
rect 9180 41012 9186 41064
rect 10042 41012 10048 41064
rect 10100 41012 10106 41064
rect 10781 41055 10839 41061
rect 10781 41021 10793 41055
rect 10827 41052 10839 41055
rect 11146 41052 11152 41064
rect 10827 41024 11152 41052
rect 10827 41021 10839 41024
rect 10781 41015 10839 41021
rect 11146 41012 11152 41024
rect 11204 41012 11210 41064
rect 12250 41012 12256 41064
rect 12308 41012 12314 41064
rect 12989 41055 13047 41061
rect 12989 41021 13001 41055
rect 13035 41052 13047 41055
rect 13538 41052 13544 41064
rect 13035 41024 13544 41052
rect 13035 41021 13047 41024
rect 12989 41015 13047 41021
rect 13538 41012 13544 41024
rect 13596 41012 13602 41064
rect 27798 41012 27804 41064
rect 27856 41052 27862 41064
rect 28718 41052 28724 41064
rect 27856 41024 28724 41052
rect 27856 41012 27862 41024
rect 28718 41012 28724 41024
rect 28776 41012 28782 41064
rect 28810 41012 28816 41064
rect 28868 41012 28874 41064
rect 29012 41061 29040 41092
rect 28905 41055 28963 41061
rect 28905 41021 28917 41055
rect 28951 41021 28963 41055
rect 28905 41015 28963 41021
rect 28997 41055 29055 41061
rect 28997 41021 29009 41055
rect 29043 41021 29055 41055
rect 28997 41015 29055 41021
rect 27706 40944 27712 40996
rect 27764 40984 27770 40996
rect 28920 40984 28948 41015
rect 29270 41012 29276 41064
rect 29328 41012 29334 41064
rect 27764 40956 30328 40984
rect 27764 40944 27770 40956
rect 8662 40876 8668 40928
rect 8720 40876 8726 40928
rect 9674 40876 9680 40928
rect 9732 40916 9738 40928
rect 9769 40919 9827 40925
rect 9769 40916 9781 40919
rect 9732 40888 9781 40916
rect 9732 40876 9738 40888
rect 9769 40885 9781 40888
rect 9815 40885 9827 40919
rect 9769 40879 9827 40885
rect 10594 40876 10600 40928
rect 10652 40876 10658 40928
rect 11330 40876 11336 40928
rect 11388 40876 11394 40928
rect 12802 40876 12808 40928
rect 12860 40876 12866 40928
rect 12986 40876 12992 40928
rect 13044 40916 13050 40928
rect 13541 40919 13599 40925
rect 13541 40916 13553 40919
rect 13044 40888 13553 40916
rect 13044 40876 13050 40888
rect 13541 40885 13553 40888
rect 13587 40885 13599 40919
rect 13541 40879 13599 40885
rect 25038 40876 25044 40928
rect 25096 40916 25102 40928
rect 28350 40916 28356 40928
rect 25096 40888 28356 40916
rect 25096 40876 25102 40888
rect 28350 40876 28356 40888
rect 28408 40876 28414 40928
rect 28537 40919 28595 40925
rect 28537 40885 28549 40919
rect 28583 40916 28595 40919
rect 29454 40916 29460 40928
rect 28583 40888 29460 40916
rect 28583 40885 28595 40888
rect 28537 40879 28595 40885
rect 29454 40876 29460 40888
rect 29512 40876 29518 40928
rect 29546 40876 29552 40928
rect 29604 40916 29610 40928
rect 30300 40925 30328 40956
rect 29917 40919 29975 40925
rect 29917 40916 29929 40919
rect 29604 40888 29929 40916
rect 29604 40876 29610 40888
rect 29917 40885 29929 40888
rect 29963 40885 29975 40919
rect 29917 40879 29975 40885
rect 30285 40919 30343 40925
rect 30285 40885 30297 40919
rect 30331 40916 30343 40919
rect 31202 40916 31208 40928
rect 30331 40888 31208 40916
rect 30331 40885 30343 40888
rect 30285 40879 30343 40885
rect 31202 40876 31208 40888
rect 31260 40876 31266 40928
rect 1104 40826 43884 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 43884 40826
rect 1104 40752 43884 40774
rect 12250 40672 12256 40724
rect 12308 40712 12314 40724
rect 12621 40715 12679 40721
rect 12621 40712 12633 40715
rect 12308 40684 12633 40712
rect 12308 40672 12314 40684
rect 12621 40681 12633 40684
rect 12667 40681 12679 40715
rect 29362 40712 29368 40724
rect 12621 40675 12679 40681
rect 28368 40684 29368 40712
rect 13262 40536 13268 40588
rect 13320 40536 13326 40588
rect 23658 40536 23664 40588
rect 23716 40576 23722 40588
rect 25038 40576 25044 40588
rect 23716 40548 25044 40576
rect 23716 40536 23722 40548
rect 25038 40536 25044 40548
rect 25096 40536 25102 40588
rect 27890 40576 27896 40588
rect 26988 40548 27896 40576
rect 934 40468 940 40520
rect 992 40508 998 40520
rect 1581 40511 1639 40517
rect 1581 40508 1593 40511
rect 992 40480 1593 40508
rect 992 40468 998 40480
rect 1581 40477 1593 40480
rect 1627 40477 1639 40511
rect 1581 40471 1639 40477
rect 8205 40511 8263 40517
rect 8205 40477 8217 40511
rect 8251 40508 8263 40511
rect 8570 40508 8576 40520
rect 8251 40480 8576 40508
rect 8251 40477 8263 40480
rect 8205 40471 8263 40477
rect 8570 40468 8576 40480
rect 8628 40468 8634 40520
rect 8938 40468 8944 40520
rect 8996 40468 9002 40520
rect 10410 40468 10416 40520
rect 10468 40468 10474 40520
rect 11238 40468 11244 40520
rect 11296 40468 11302 40520
rect 11882 40468 11888 40520
rect 11940 40468 11946 40520
rect 14090 40468 14096 40520
rect 14148 40468 14154 40520
rect 15102 40468 15108 40520
rect 15160 40468 15166 40520
rect 15930 40468 15936 40520
rect 15988 40468 15994 40520
rect 23474 40468 23480 40520
rect 23532 40508 23538 40520
rect 24397 40511 24455 40517
rect 24397 40508 24409 40511
rect 23532 40480 24409 40508
rect 23532 40468 23538 40480
rect 24397 40477 24409 40480
rect 24443 40477 24455 40511
rect 24397 40471 24455 40477
rect 24578 40468 24584 40520
rect 24636 40468 24642 40520
rect 26988 40517 27016 40548
rect 27890 40536 27896 40548
rect 27948 40536 27954 40588
rect 28261 40579 28319 40585
rect 28261 40545 28273 40579
rect 28307 40576 28319 40579
rect 28368 40576 28396 40684
rect 29362 40672 29368 40684
rect 29420 40712 29426 40724
rect 29730 40712 29736 40724
rect 29420 40684 29736 40712
rect 29420 40672 29426 40684
rect 29730 40672 29736 40684
rect 29788 40672 29794 40724
rect 29840 40616 30880 40644
rect 29840 40588 29868 40616
rect 29822 40576 29828 40588
rect 28307 40548 28396 40576
rect 29104 40548 29828 40576
rect 28307 40545 28319 40548
rect 28261 40539 28319 40545
rect 26881 40511 26939 40517
rect 26881 40477 26893 40511
rect 26927 40477 26939 40511
rect 26881 40471 26939 40477
rect 26973 40511 27031 40517
rect 26973 40477 26985 40511
rect 27019 40477 27031 40511
rect 26973 40471 27031 40477
rect 27341 40511 27399 40517
rect 27341 40477 27353 40511
rect 27387 40477 27399 40511
rect 27341 40471 27399 40477
rect 8018 40400 8024 40452
rect 8076 40440 8082 40452
rect 9585 40443 9643 40449
rect 9585 40440 9597 40443
rect 8076 40412 9597 40440
rect 8076 40400 8082 40412
rect 9585 40409 9597 40412
rect 9631 40409 9643 40443
rect 9585 40403 9643 40409
rect 10870 40400 10876 40452
rect 10928 40440 10934 40452
rect 11793 40443 11851 40449
rect 11793 40440 11805 40443
rect 10928 40412 11805 40440
rect 10928 40400 10934 40412
rect 11793 40409 11805 40412
rect 11839 40409 11851 40443
rect 11793 40403 11851 40409
rect 12989 40443 13047 40449
rect 12989 40409 13001 40443
rect 13035 40440 13047 40443
rect 14737 40443 14795 40449
rect 14737 40440 14749 40443
rect 13035 40412 14749 40440
rect 13035 40409 13047 40412
rect 12989 40403 13047 40409
rect 14737 40409 14749 40412
rect 14783 40409 14795 40443
rect 14737 40403 14795 40409
rect 24210 40400 24216 40452
rect 24268 40440 24274 40452
rect 24268 40412 25544 40440
rect 24268 40400 24274 40412
rect 8757 40375 8815 40381
rect 8757 40341 8769 40375
rect 8803 40372 8815 40375
rect 8846 40372 8852 40384
rect 8803 40344 8852 40372
rect 8803 40341 8815 40344
rect 8757 40335 8815 40341
rect 8846 40332 8852 40344
rect 8904 40332 8910 40384
rect 10962 40332 10968 40384
rect 11020 40332 11026 40384
rect 12434 40332 12440 40384
rect 12492 40372 12498 40384
rect 12529 40375 12587 40381
rect 12529 40372 12541 40375
rect 12492 40344 12541 40372
rect 12492 40332 12498 40344
rect 12529 40341 12541 40344
rect 12575 40341 12587 40375
rect 12529 40335 12587 40341
rect 13081 40375 13139 40381
rect 13081 40341 13093 40375
rect 13127 40372 13139 40375
rect 13170 40372 13176 40384
rect 13127 40344 13176 40372
rect 13127 40341 13139 40344
rect 13081 40335 13139 40341
rect 13170 40332 13176 40344
rect 13228 40332 13234 40384
rect 15746 40332 15752 40384
rect 15804 40332 15810 40384
rect 16482 40332 16488 40384
rect 16540 40332 16546 40384
rect 24762 40332 24768 40384
rect 24820 40332 24826 40384
rect 25516 40381 25544 40412
rect 26234 40400 26240 40452
rect 26292 40440 26298 40452
rect 26896 40440 26924 40471
rect 27356 40440 27384 40471
rect 27430 40468 27436 40520
rect 27488 40468 27494 40520
rect 29104 40517 29132 40548
rect 29822 40536 29828 40548
rect 29880 40536 29886 40588
rect 30098 40536 30104 40588
rect 30156 40576 30162 40588
rect 30852 40585 30880 40616
rect 30837 40579 30895 40585
rect 30156 40548 30512 40576
rect 30156 40536 30162 40548
rect 29089 40511 29147 40517
rect 29089 40510 29101 40511
rect 29012 40508 29101 40510
rect 27540 40482 29101 40508
rect 27540 40480 29040 40482
rect 27540 40440 27568 40480
rect 29089 40477 29101 40482
rect 29135 40477 29147 40511
rect 29089 40471 29147 40477
rect 29178 40468 29184 40520
rect 29236 40468 29242 40520
rect 30484 40517 30512 40548
rect 30837 40545 30849 40579
rect 30883 40576 30895 40579
rect 31297 40579 31355 40585
rect 31297 40576 31309 40579
rect 30883 40548 31309 40576
rect 30883 40545 30895 40548
rect 30837 40539 30895 40545
rect 31297 40545 31309 40548
rect 31343 40545 31355 40579
rect 31297 40539 31355 40545
rect 29641 40511 29699 40517
rect 29641 40477 29653 40511
rect 29687 40508 29699 40511
rect 30285 40511 30343 40517
rect 30285 40508 30297 40511
rect 29687 40480 30297 40508
rect 29687 40477 29699 40480
rect 29641 40471 29699 40477
rect 30285 40477 30297 40480
rect 30331 40477 30343 40511
rect 30285 40471 30343 40477
rect 30469 40511 30527 40517
rect 30469 40477 30481 40511
rect 30515 40477 30527 40511
rect 30469 40471 30527 40477
rect 30742 40468 30748 40520
rect 30800 40468 30806 40520
rect 31018 40468 31024 40520
rect 31076 40468 31082 40520
rect 31478 40468 31484 40520
rect 31536 40468 31542 40520
rect 26292 40412 27568 40440
rect 29012 40412 30328 40440
rect 26292 40400 26298 40412
rect 29012 40384 29040 40412
rect 25501 40375 25559 40381
rect 25501 40341 25513 40375
rect 25547 40372 25559 40375
rect 26602 40372 26608 40384
rect 25547 40344 26608 40372
rect 25547 40341 25559 40344
rect 25501 40335 25559 40341
rect 26602 40332 26608 40344
rect 26660 40332 26666 40384
rect 26694 40332 26700 40384
rect 26752 40332 26758 40384
rect 27154 40332 27160 40384
rect 27212 40332 27218 40384
rect 27614 40332 27620 40384
rect 27672 40332 27678 40384
rect 27890 40332 27896 40384
rect 27948 40332 27954 40384
rect 28810 40332 28816 40384
rect 28868 40332 28874 40384
rect 28994 40332 29000 40384
rect 29052 40332 29058 40384
rect 29362 40332 29368 40384
rect 29420 40332 29426 40384
rect 29730 40332 29736 40384
rect 29788 40372 29794 40384
rect 30193 40375 30251 40381
rect 30193 40372 30205 40375
rect 29788 40344 30205 40372
rect 29788 40332 29794 40344
rect 30193 40341 30205 40344
rect 30239 40341 30251 40375
rect 30300 40372 30328 40412
rect 30374 40400 30380 40452
rect 30432 40440 30438 40452
rect 31205 40443 31263 40449
rect 31205 40440 31217 40443
rect 30432 40412 31217 40440
rect 30432 40400 30438 40412
rect 31205 40409 31217 40412
rect 31251 40409 31263 40443
rect 31205 40403 31263 40409
rect 30558 40372 30564 40384
rect 30300 40344 30564 40372
rect 30193 40335 30251 40341
rect 30558 40332 30564 40344
rect 30616 40332 30622 40384
rect 30653 40375 30711 40381
rect 30653 40341 30665 40375
rect 30699 40372 30711 40375
rect 31294 40372 31300 40384
rect 30699 40344 31300 40372
rect 30699 40341 30711 40344
rect 30653 40335 30711 40341
rect 31294 40332 31300 40344
rect 31352 40332 31358 40384
rect 31662 40332 31668 40384
rect 31720 40332 31726 40384
rect 1104 40282 43884 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 43884 40282
rect 1104 40208 43884 40230
rect 8110 40128 8116 40180
rect 8168 40168 8174 40180
rect 8205 40171 8263 40177
rect 8205 40168 8217 40171
rect 8168 40140 8217 40168
rect 8168 40128 8174 40140
rect 8205 40137 8217 40140
rect 8251 40137 8263 40171
rect 8205 40131 8263 40137
rect 10042 40128 10048 40180
rect 10100 40168 10106 40180
rect 10413 40171 10471 40177
rect 10413 40168 10425 40171
rect 10100 40140 10425 40168
rect 10100 40128 10106 40140
rect 10413 40137 10425 40140
rect 10459 40137 10471 40171
rect 10413 40131 10471 40137
rect 10781 40171 10839 40177
rect 10781 40137 10793 40171
rect 10827 40168 10839 40171
rect 11330 40168 11336 40180
rect 10827 40140 11336 40168
rect 10827 40137 10839 40140
rect 10781 40131 10839 40137
rect 11330 40128 11336 40140
rect 11388 40128 11394 40180
rect 13541 40171 13599 40177
rect 13541 40137 13553 40171
rect 13587 40168 13599 40171
rect 14090 40168 14096 40180
rect 13587 40140 14096 40168
rect 13587 40137 13599 40140
rect 13541 40131 13599 40137
rect 14090 40128 14096 40140
rect 14148 40128 14154 40180
rect 15105 40171 15163 40177
rect 15105 40137 15117 40171
rect 15151 40137 15163 40171
rect 15105 40131 15163 40137
rect 15473 40171 15531 40177
rect 15473 40137 15485 40171
rect 15519 40168 15531 40171
rect 16482 40168 16488 40180
rect 15519 40140 16488 40168
rect 15519 40137 15531 40140
rect 15473 40131 15531 40137
rect 9582 40060 9588 40112
rect 9640 40100 9646 40112
rect 9953 40103 10011 40109
rect 9953 40100 9965 40103
rect 9640 40072 9965 40100
rect 9640 40060 9646 40072
rect 9953 40069 9965 40072
rect 9999 40069 10011 40103
rect 9953 40063 10011 40069
rect 12428 40103 12486 40109
rect 12428 40069 12440 40103
rect 12474 40100 12486 40103
rect 12802 40100 12808 40112
rect 12474 40072 12808 40100
rect 12474 40069 12486 40072
rect 12428 40063 12486 40069
rect 12802 40060 12808 40072
rect 12860 40060 12866 40112
rect 15120 40100 15148 40131
rect 16482 40128 16488 40140
rect 16540 40128 16546 40180
rect 25593 40171 25651 40177
rect 25593 40137 25605 40171
rect 25639 40168 25651 40171
rect 27246 40168 27252 40180
rect 25639 40140 27252 40168
rect 25639 40137 25651 40140
rect 25593 40131 25651 40137
rect 27246 40128 27252 40140
rect 27304 40128 27310 40180
rect 28997 40171 29055 40177
rect 27356 40140 28028 40168
rect 24210 40100 24216 40112
rect 14844 40072 15148 40100
rect 23860 40072 24216 40100
rect 6270 39992 6276 40044
rect 6328 40032 6334 40044
rect 7193 40035 7251 40041
rect 7193 40032 7205 40035
rect 6328 40004 7205 40032
rect 6328 39992 6334 40004
rect 7193 40001 7205 40004
rect 7239 40001 7251 40035
rect 7193 39995 7251 40001
rect 8573 40035 8631 40041
rect 8573 40001 8585 40035
rect 8619 40032 8631 40035
rect 8846 40032 8852 40044
rect 8619 40004 8852 40032
rect 8619 40001 8631 40004
rect 8573 39995 8631 40001
rect 8846 39992 8852 40004
rect 8904 40032 8910 40044
rect 9490 40032 9496 40044
rect 8904 40004 9496 40032
rect 8904 39992 8910 40004
rect 9490 39992 9496 40004
rect 9548 39992 9554 40044
rect 13262 39992 13268 40044
rect 13320 40032 13326 40044
rect 14734 40032 14740 40044
rect 13320 40004 14740 40032
rect 13320 39992 13326 40004
rect 14734 39992 14740 40004
rect 14792 39992 14798 40044
rect 6549 39967 6607 39973
rect 6549 39933 6561 39967
rect 6595 39964 6607 39967
rect 6730 39964 6736 39976
rect 6595 39936 6736 39964
rect 6595 39933 6607 39936
rect 6549 39927 6607 39933
rect 6730 39924 6736 39936
rect 6788 39924 6794 39976
rect 8665 39967 8723 39973
rect 8665 39933 8677 39967
rect 8711 39933 8723 39967
rect 8665 39927 8723 39933
rect 8757 39967 8815 39973
rect 8757 39933 8769 39967
rect 8803 39964 8815 39967
rect 9214 39964 9220 39976
rect 8803 39936 9220 39964
rect 8803 39933 8815 39936
rect 8757 39927 8815 39933
rect 8680 39896 8708 39927
rect 9214 39924 9220 39936
rect 9272 39924 9278 39976
rect 9306 39924 9312 39976
rect 9364 39924 9370 39976
rect 9398 39924 9404 39976
rect 9456 39924 9462 39976
rect 10778 39924 10784 39976
rect 10836 39964 10842 39976
rect 10873 39967 10931 39973
rect 10873 39964 10885 39967
rect 10836 39936 10885 39964
rect 10836 39924 10842 39936
rect 10873 39933 10885 39936
rect 10919 39933 10931 39967
rect 10873 39927 10931 39933
rect 10965 39967 11023 39973
rect 10965 39933 10977 39967
rect 11011 39933 11023 39967
rect 10965 39927 11023 39933
rect 9416 39896 9444 39924
rect 10980 39896 11008 39927
rect 11974 39924 11980 39976
rect 12032 39964 12038 39976
rect 12161 39967 12219 39973
rect 12161 39964 12173 39967
rect 12032 39936 12173 39964
rect 12032 39924 12038 39936
rect 12161 39933 12173 39936
rect 12207 39933 12219 39967
rect 12161 39927 12219 39933
rect 8680 39868 9444 39896
rect 9784 39868 11008 39896
rect 9784 39840 9812 39868
rect 7098 39788 7104 39840
rect 7156 39788 7162 39840
rect 7834 39788 7840 39840
rect 7892 39788 7898 39840
rect 9766 39788 9772 39840
rect 9824 39788 9830 39840
rect 10980 39828 11008 39868
rect 13280 39828 13308 39992
rect 13630 39924 13636 39976
rect 13688 39924 13694 39976
rect 14461 39967 14519 39973
rect 14461 39933 14473 39967
rect 14507 39964 14519 39967
rect 14844 39964 14872 40072
rect 22925 40035 22983 40041
rect 14507 39936 14872 39964
rect 15028 40004 15700 40032
rect 14507 39933 14519 39936
rect 14461 39927 14519 39933
rect 15028 39896 15056 40004
rect 15286 39924 15292 39976
rect 15344 39964 15350 39976
rect 15672 39973 15700 40004
rect 22925 40001 22937 40035
rect 22971 40032 22983 40035
rect 23860 40032 23888 40072
rect 24210 40060 24216 40072
rect 24268 40060 24274 40112
rect 24480 40103 24538 40109
rect 24480 40069 24492 40103
rect 24526 40100 24538 40103
rect 24762 40100 24768 40112
rect 24526 40072 24768 40100
rect 24526 40069 24538 40072
rect 24480 40063 24538 40069
rect 24762 40060 24768 40072
rect 24820 40060 24826 40112
rect 26694 40100 26700 40112
rect 26528 40072 26700 40100
rect 22971 40004 23888 40032
rect 22971 40001 22983 40004
rect 22925 39995 22983 40001
rect 23934 39992 23940 40044
rect 23992 39992 23998 40044
rect 26528 40041 26556 40072
rect 26694 40060 26700 40072
rect 26752 40100 26758 40112
rect 27356 40100 27384 40140
rect 28000 40112 28028 40140
rect 28997 40137 29009 40171
rect 29043 40137 29055 40171
rect 28997 40131 29055 40137
rect 26752 40072 27384 40100
rect 26752 40060 26758 40072
rect 27614 40060 27620 40112
rect 27672 40100 27678 40112
rect 27862 40103 27920 40109
rect 27862 40100 27874 40103
rect 27672 40072 27874 40100
rect 27672 40060 27678 40072
rect 27862 40069 27874 40072
rect 27908 40069 27920 40103
rect 27862 40063 27920 40069
rect 27982 40060 27988 40112
rect 28040 40060 28046 40112
rect 29012 40100 29040 40131
rect 29638 40128 29644 40180
rect 29696 40168 29702 40180
rect 30469 40171 30527 40177
rect 30469 40168 30481 40171
rect 29696 40140 30481 40168
rect 29696 40128 29702 40140
rect 30469 40137 30481 40140
rect 30515 40137 30527 40171
rect 30469 40131 30527 40137
rect 30558 40128 30564 40180
rect 30616 40168 30622 40180
rect 31205 40171 31263 40177
rect 31205 40168 31217 40171
rect 30616 40140 31217 40168
rect 30616 40128 30622 40140
rect 31205 40137 31217 40140
rect 31251 40137 31263 40171
rect 31205 40131 31263 40137
rect 29012 40072 30604 40100
rect 26513 40035 26571 40041
rect 24136 40004 26464 40032
rect 15565 39967 15623 39973
rect 15565 39964 15577 39967
rect 15344 39936 15577 39964
rect 15344 39924 15350 39936
rect 15565 39933 15577 39936
rect 15611 39933 15623 39967
rect 15565 39927 15623 39933
rect 15657 39967 15715 39973
rect 15657 39933 15669 39967
rect 15703 39933 15715 39967
rect 15657 39927 15715 39933
rect 16850 39924 16856 39976
rect 16908 39924 16914 39976
rect 17770 39924 17776 39976
rect 17828 39924 17834 39976
rect 23474 39924 23480 39976
rect 23532 39964 23538 39976
rect 23753 39967 23811 39973
rect 23753 39964 23765 39967
rect 23532 39936 23765 39964
rect 23532 39924 23538 39936
rect 23753 39933 23765 39936
rect 23799 39933 23811 39967
rect 23753 39927 23811 39933
rect 24136 39896 24164 40004
rect 24213 39967 24271 39973
rect 24213 39933 24225 39967
rect 24259 39933 24271 39967
rect 26436 39964 26464 40004
rect 26513 40001 26525 40035
rect 26559 40001 26571 40035
rect 26513 39995 26571 40001
rect 26602 39992 26608 40044
rect 26660 40032 26666 40044
rect 27430 40032 27436 40044
rect 26660 40004 27436 40032
rect 26660 39992 26666 40004
rect 27430 39992 27436 40004
rect 27488 39992 27494 40044
rect 27540 40030 29040 40032
rect 29178 40030 29184 40044
rect 27540 40004 29184 40030
rect 27540 39964 27568 40004
rect 29012 40002 29184 40004
rect 29178 39992 29184 40002
rect 29236 39992 29242 40044
rect 29356 40035 29414 40041
rect 29356 40001 29368 40035
rect 29402 40032 29414 40035
rect 30374 40032 30380 40044
rect 29402 40004 30380 40032
rect 29402 40001 29414 40004
rect 29356 39995 29414 40001
rect 30374 39992 30380 40004
rect 30432 39992 30438 40044
rect 30576 40041 30604 40072
rect 30668 40072 31524 40100
rect 30561 40035 30619 40041
rect 30561 40001 30573 40035
rect 30607 40001 30619 40035
rect 30561 39995 30619 40001
rect 26436 39936 27568 39964
rect 27617 39967 27675 39973
rect 24213 39927 24271 39933
rect 27617 39933 27629 39967
rect 27663 39933 27675 39967
rect 27617 39927 27675 39933
rect 13372 39868 15056 39896
rect 15580 39868 24164 39896
rect 13372 39840 13400 39868
rect 15580 39840 15608 39868
rect 10980 39800 13308 39828
rect 13354 39788 13360 39840
rect 13412 39788 13418 39840
rect 13814 39788 13820 39840
rect 13872 39828 13878 39840
rect 14277 39831 14335 39837
rect 14277 39828 14289 39831
rect 13872 39800 14289 39828
rect 13872 39788 13878 39800
rect 14277 39797 14289 39800
rect 14323 39797 14335 39831
rect 14277 39791 14335 39797
rect 15010 39788 15016 39840
rect 15068 39788 15074 39840
rect 15562 39788 15568 39840
rect 15620 39788 15626 39840
rect 17218 39788 17224 39840
rect 17276 39828 17282 39840
rect 17497 39831 17555 39837
rect 17497 39828 17509 39831
rect 17276 39800 17509 39828
rect 17276 39788 17282 39800
rect 17497 39797 17509 39800
rect 17543 39797 17555 39831
rect 17497 39791 17555 39797
rect 18322 39788 18328 39840
rect 18380 39788 18386 39840
rect 22557 39831 22615 39837
rect 22557 39797 22569 39831
rect 22603 39828 22615 39831
rect 23290 39828 23296 39840
rect 22603 39800 23296 39828
rect 22603 39797 22615 39800
rect 22557 39791 22615 39797
rect 23290 39788 23296 39800
rect 23348 39788 23354 39840
rect 23658 39788 23664 39840
rect 23716 39788 23722 39840
rect 24118 39788 24124 39840
rect 24176 39788 24182 39840
rect 24228 39828 24256 39927
rect 26697 39899 26755 39905
rect 26697 39896 26709 39899
rect 25332 39868 26709 39896
rect 25332 39840 25360 39868
rect 26697 39865 26709 39868
rect 26743 39865 26755 39899
rect 27522 39896 27528 39908
rect 26697 39859 26755 39865
rect 27172 39868 27528 39896
rect 24486 39828 24492 39840
rect 24228 39800 24492 39828
rect 24486 39788 24492 39800
rect 24544 39788 24550 39840
rect 25314 39788 25320 39840
rect 25372 39788 25378 39840
rect 25961 39831 26019 39837
rect 25961 39797 25973 39831
rect 26007 39828 26019 39831
rect 26329 39831 26387 39837
rect 26329 39828 26341 39831
rect 26007 39800 26341 39828
rect 26007 39797 26019 39800
rect 25961 39791 26019 39797
rect 26329 39797 26341 39800
rect 26375 39828 26387 39831
rect 27172 39828 27200 39868
rect 27522 39856 27528 39868
rect 27580 39856 27586 39908
rect 27632 39840 27660 39927
rect 28902 39924 28908 39976
rect 28960 39964 28966 39976
rect 29089 39967 29147 39973
rect 29089 39964 29101 39967
rect 28960 39936 29101 39964
rect 28960 39924 28966 39936
rect 29089 39933 29101 39936
rect 29135 39933 29147 39967
rect 30668 39964 30696 40072
rect 31496 40041 31524 40072
rect 31389 40035 31447 40041
rect 31389 40001 31401 40035
rect 31435 40001 31447 40035
rect 31389 39995 31447 40001
rect 31481 40035 31539 40041
rect 31481 40001 31493 40035
rect 31527 40032 31539 40035
rect 31527 40004 33364 40032
rect 31527 40001 31539 40004
rect 31481 39995 31539 40001
rect 29089 39927 29147 39933
rect 30116 39936 30696 39964
rect 26375 39800 27200 39828
rect 27249 39831 27307 39837
rect 26375 39797 26387 39800
rect 26329 39791 26387 39797
rect 27249 39797 27261 39831
rect 27295 39828 27307 39831
rect 27430 39828 27436 39840
rect 27295 39800 27436 39828
rect 27295 39797 27307 39800
rect 27249 39791 27307 39797
rect 27430 39788 27436 39800
rect 27488 39788 27494 39840
rect 27614 39788 27620 39840
rect 27672 39828 27678 39840
rect 28920 39828 28948 39924
rect 27672 39800 28948 39828
rect 27672 39788 27678 39800
rect 29086 39788 29092 39840
rect 29144 39828 29150 39840
rect 30116 39828 30144 39936
rect 30558 39856 30564 39908
rect 30616 39896 30622 39908
rect 31404 39896 31432 39995
rect 32401 39899 32459 39905
rect 32401 39896 32413 39899
rect 30616 39868 31340 39896
rect 31404 39868 32413 39896
rect 30616 39856 30622 39868
rect 29144 39800 30144 39828
rect 31312 39828 31340 39868
rect 32401 39865 32413 39868
rect 32447 39896 32459 39899
rect 33226 39896 33232 39908
rect 32447 39868 33232 39896
rect 32447 39865 32459 39868
rect 32401 39859 32459 39865
rect 33226 39856 33232 39868
rect 33284 39856 33290 39908
rect 31665 39831 31723 39837
rect 31665 39828 31677 39831
rect 31312 39800 31677 39828
rect 29144 39788 29150 39800
rect 31665 39797 31677 39800
rect 31711 39797 31723 39831
rect 31665 39791 31723 39797
rect 32769 39831 32827 39837
rect 32769 39797 32781 39831
rect 32815 39828 32827 39831
rect 33336 39828 33364 40004
rect 33502 39828 33508 39840
rect 32815 39800 33508 39828
rect 32815 39797 32827 39800
rect 32769 39791 32827 39797
rect 33502 39788 33508 39800
rect 33560 39788 33566 39840
rect 1104 39738 43884 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 43884 39738
rect 1104 39664 43884 39686
rect 8941 39627 8999 39633
rect 8941 39624 8953 39627
rect 7116 39596 8953 39624
rect 1210 39448 1216 39500
rect 1268 39488 1274 39500
rect 1857 39491 1915 39497
rect 1857 39488 1869 39491
rect 1268 39460 1869 39488
rect 1268 39448 1274 39460
rect 1857 39457 1869 39460
rect 1903 39457 1915 39491
rect 1857 39451 1915 39457
rect 6362 39448 6368 39500
rect 6420 39448 6426 39500
rect 6733 39491 6791 39497
rect 6733 39457 6745 39491
rect 6779 39488 6791 39491
rect 7116 39488 7144 39596
rect 8941 39593 8953 39596
rect 8987 39593 8999 39627
rect 8941 39587 8999 39593
rect 9122 39584 9128 39636
rect 9180 39584 9186 39636
rect 11146 39584 11152 39636
rect 11204 39624 11210 39636
rect 11241 39627 11299 39633
rect 11241 39624 11253 39627
rect 11204 39596 11253 39624
rect 11204 39584 11210 39596
rect 11241 39593 11253 39596
rect 11287 39593 11299 39627
rect 11241 39587 11299 39593
rect 13538 39584 13544 39636
rect 13596 39584 13602 39636
rect 20993 39627 21051 39633
rect 20993 39593 21005 39627
rect 21039 39624 21051 39627
rect 22370 39624 22376 39636
rect 21039 39596 22376 39624
rect 21039 39593 21051 39596
rect 20993 39587 21051 39593
rect 22370 39584 22376 39596
rect 22428 39624 22434 39636
rect 26234 39624 26240 39636
rect 22428 39596 25084 39624
rect 22428 39584 22434 39596
rect 8757 39559 8815 39565
rect 8757 39525 8769 39559
rect 8803 39556 8815 39559
rect 9140 39556 9168 39584
rect 9766 39556 9772 39568
rect 8803 39528 9168 39556
rect 9508 39528 9772 39556
rect 8803 39525 8815 39528
rect 8757 39519 8815 39525
rect 6779 39460 7144 39488
rect 6779 39457 6791 39460
rect 6733 39451 6791 39457
rect 7374 39448 7380 39500
rect 7432 39448 7438 39500
rect 9508 39497 9536 39528
rect 9766 39516 9772 39528
rect 9824 39516 9830 39568
rect 9493 39491 9551 39497
rect 9493 39488 9505 39491
rect 9140 39460 9505 39488
rect 1581 39423 1639 39429
rect 1581 39389 1593 39423
rect 1627 39420 1639 39423
rect 1627 39392 2774 39420
rect 1627 39389 1639 39392
rect 1581 39383 1639 39389
rect 2746 39352 2774 39392
rect 5994 39380 6000 39432
rect 6052 39380 6058 39432
rect 6380 39420 6408 39448
rect 9140 39420 9168 39460
rect 9493 39457 9505 39460
rect 9539 39457 9551 39491
rect 9493 39451 9551 39457
rect 24320 39460 24532 39488
rect 6380 39392 9168 39420
rect 9309 39423 9367 39429
rect 9309 39389 9321 39423
rect 9355 39420 9367 39423
rect 9674 39420 9680 39432
rect 9355 39392 9680 39420
rect 9355 39389 9367 39392
rect 9309 39383 9367 39389
rect 9674 39380 9680 39392
rect 9732 39380 9738 39432
rect 9766 39380 9772 39432
rect 9824 39420 9830 39432
rect 9861 39423 9919 39429
rect 9861 39420 9873 39423
rect 9824 39392 9873 39420
rect 9824 39380 9830 39392
rect 9861 39389 9873 39392
rect 9907 39389 9919 39423
rect 9861 39383 9919 39389
rect 10128 39423 10186 39429
rect 10128 39389 10140 39423
rect 10174 39420 10186 39423
rect 10594 39420 10600 39432
rect 10174 39392 10600 39420
rect 10174 39389 10186 39392
rect 10128 39383 10186 39389
rect 10594 39380 10600 39392
rect 10652 39380 10658 39432
rect 11514 39380 11520 39432
rect 11572 39380 11578 39432
rect 11974 39380 11980 39432
rect 12032 39420 12038 39432
rect 12434 39429 12440 39432
rect 12161 39423 12219 39429
rect 12161 39420 12173 39423
rect 12032 39392 12173 39420
rect 12032 39380 12038 39392
rect 12161 39389 12173 39392
rect 12207 39389 12219 39423
rect 12161 39383 12219 39389
rect 12428 39383 12440 39429
rect 12492 39420 12498 39432
rect 12492 39392 12528 39420
rect 12434 39380 12440 39383
rect 12492 39380 12498 39392
rect 14642 39380 14648 39432
rect 14700 39420 14706 39432
rect 16577 39423 16635 39429
rect 16577 39420 16589 39423
rect 14700 39392 16589 39420
rect 14700 39380 14706 39392
rect 16577 39389 16589 39392
rect 16623 39420 16635 39423
rect 17126 39420 17132 39432
rect 16623 39392 17132 39420
rect 16623 39389 16635 39392
rect 16577 39383 16635 39389
rect 17126 39380 17132 39392
rect 17184 39380 17190 39432
rect 17218 39380 17224 39432
rect 17276 39380 17282 39432
rect 18138 39380 18144 39432
rect 18196 39380 18202 39432
rect 22649 39423 22707 39429
rect 22649 39389 22661 39423
rect 22695 39420 22707 39423
rect 24320 39420 24348 39460
rect 24504 39432 24532 39460
rect 22695 39392 24348 39420
rect 22695 39389 22707 39392
rect 22649 39383 22707 39389
rect 24394 39380 24400 39432
rect 24452 39380 24458 39432
rect 24486 39380 24492 39432
rect 24544 39380 24550 39432
rect 25056 39420 25084 39596
rect 25148 39596 26240 39624
rect 25148 39497 25176 39596
rect 26234 39584 26240 39596
rect 26292 39584 26298 39636
rect 26326 39584 26332 39636
rect 26384 39624 26390 39636
rect 28169 39627 28227 39633
rect 28169 39624 28181 39627
rect 26384 39596 28181 39624
rect 26384 39584 26390 39596
rect 28169 39593 28181 39596
rect 28215 39593 28227 39627
rect 28169 39587 28227 39593
rect 27062 39516 27068 39568
rect 27120 39556 27126 39568
rect 27614 39556 27620 39568
rect 27120 39528 27620 39556
rect 27120 39516 27126 39528
rect 27614 39516 27620 39528
rect 27672 39516 27678 39568
rect 25133 39491 25191 39497
rect 25133 39457 25145 39491
rect 25179 39457 25191 39491
rect 25958 39488 25964 39500
rect 25133 39451 25191 39457
rect 25240 39460 25964 39488
rect 25240 39420 25268 39460
rect 25958 39448 25964 39460
rect 26016 39448 26022 39500
rect 27890 39488 27896 39500
rect 27080 39460 27896 39488
rect 27080 39432 27108 39460
rect 27890 39448 27896 39460
rect 27948 39488 27954 39500
rect 28718 39488 28724 39500
rect 27948 39460 28724 39488
rect 27948 39448 27954 39460
rect 28718 39448 28724 39460
rect 28776 39448 28782 39500
rect 25056 39392 25268 39420
rect 25314 39380 25320 39432
rect 25372 39380 25378 39432
rect 26053 39423 26111 39429
rect 26053 39389 26065 39423
rect 26099 39420 26111 39423
rect 26878 39420 26884 39432
rect 26099 39392 26884 39420
rect 26099 39389 26111 39392
rect 26053 39383 26111 39389
rect 26878 39380 26884 39392
rect 26936 39380 26942 39432
rect 27062 39380 27068 39432
rect 27120 39380 27126 39432
rect 27154 39380 27160 39432
rect 27212 39380 27218 39432
rect 27246 39380 27252 39432
rect 27304 39420 27310 39432
rect 27525 39423 27583 39429
rect 27525 39420 27537 39423
rect 27304 39392 27537 39420
rect 27304 39380 27310 39392
rect 27525 39389 27537 39392
rect 27571 39389 27583 39423
rect 27525 39383 27583 39389
rect 28261 39423 28319 39429
rect 28261 39389 28273 39423
rect 28307 39389 28319 39423
rect 28261 39383 28319 39389
rect 3145 39355 3203 39361
rect 3145 39352 3157 39355
rect 2746 39324 3157 39352
rect 3145 39321 3157 39324
rect 3191 39352 3203 39355
rect 7285 39355 7343 39361
rect 3191 39324 6684 39352
rect 3191 39321 3203 39324
rect 3145 39315 3203 39321
rect 6546 39244 6552 39296
rect 6604 39244 6610 39296
rect 6656 39284 6684 39324
rect 7285 39321 7297 39355
rect 7331 39352 7343 39355
rect 7622 39355 7680 39361
rect 7622 39352 7634 39355
rect 7331 39324 7634 39352
rect 7331 39321 7343 39324
rect 7285 39315 7343 39321
rect 7622 39321 7634 39324
rect 7668 39321 7680 39355
rect 14912 39355 14970 39361
rect 7622 39315 7680 39321
rect 7760 39324 11376 39352
rect 7760 39284 7788 39324
rect 11348 39296 11376 39324
rect 14912 39321 14924 39355
rect 14958 39352 14970 39355
rect 15746 39352 15752 39364
rect 14958 39324 15752 39352
rect 14958 39321 14970 39324
rect 14912 39315 14970 39321
rect 15746 39312 15752 39324
rect 15804 39312 15810 39364
rect 16844 39355 16902 39361
rect 16844 39321 16856 39355
rect 16890 39352 16902 39355
rect 17236 39352 17264 39380
rect 18969 39355 19027 39361
rect 18969 39352 18981 39355
rect 16890 39324 17264 39352
rect 17328 39324 18981 39352
rect 16890 39321 16902 39324
rect 16844 39315 16902 39321
rect 6656 39256 7788 39284
rect 9398 39244 9404 39296
rect 9456 39244 9462 39296
rect 11330 39244 11336 39296
rect 11388 39244 11394 39296
rect 12069 39287 12127 39293
rect 12069 39253 12081 39287
rect 12115 39284 12127 39287
rect 12526 39284 12532 39296
rect 12115 39256 12532 39284
rect 12115 39253 12127 39256
rect 12069 39247 12127 39253
rect 12526 39244 12532 39256
rect 12584 39244 12590 39296
rect 16022 39244 16028 39296
rect 16080 39244 16086 39296
rect 16390 39244 16396 39296
rect 16448 39284 16454 39296
rect 17328 39284 17356 39324
rect 18969 39321 18981 39324
rect 19015 39352 19027 39355
rect 22094 39352 22100 39364
rect 19015 39324 22100 39352
rect 19015 39321 19027 39324
rect 18969 39315 19027 39321
rect 22094 39312 22100 39324
rect 22152 39312 22158 39364
rect 22916 39355 22974 39361
rect 22916 39321 22928 39355
rect 22962 39352 22974 39355
rect 24118 39352 24124 39364
rect 22962 39324 24124 39352
rect 22962 39321 22974 39324
rect 22916 39315 22974 39321
rect 24118 39312 24124 39324
rect 24176 39312 24182 39364
rect 24854 39312 24860 39364
rect 24912 39352 24918 39364
rect 25332 39352 25360 39380
rect 24912 39324 25360 39352
rect 26320 39355 26378 39361
rect 24912 39312 24918 39324
rect 26320 39321 26332 39355
rect 26366 39352 26378 39355
rect 27172 39352 27200 39380
rect 28276 39352 28304 39383
rect 28902 39380 28908 39432
rect 28960 39420 28966 39432
rect 29549 39423 29607 39429
rect 29549 39420 29561 39423
rect 28960 39392 29561 39420
rect 28960 39380 28966 39392
rect 29549 39389 29561 39392
rect 29595 39420 29607 39423
rect 31021 39423 31079 39429
rect 31021 39420 31033 39423
rect 29595 39392 31033 39420
rect 29595 39389 29607 39392
rect 29549 39383 29607 39389
rect 31021 39389 31033 39392
rect 31067 39389 31079 39423
rect 31021 39383 31079 39389
rect 31288 39423 31346 39429
rect 31288 39389 31300 39423
rect 31334 39420 31346 39423
rect 31662 39420 31668 39432
rect 31334 39392 31668 39420
rect 31334 39389 31346 39392
rect 31288 39383 31346 39389
rect 31662 39380 31668 39392
rect 31720 39380 31726 39432
rect 43349 39423 43407 39429
rect 43349 39389 43361 39423
rect 43395 39420 43407 39423
rect 43395 39392 43852 39420
rect 43395 39389 43407 39392
rect 43349 39383 43407 39389
rect 43824 39364 43852 39392
rect 26366 39324 27200 39352
rect 27264 39324 28304 39352
rect 26366 39321 26378 39324
rect 26320 39315 26378 39321
rect 27264 39296 27292 39324
rect 29362 39312 29368 39364
rect 29420 39352 29426 39364
rect 29794 39355 29852 39361
rect 29794 39352 29806 39355
rect 29420 39324 29806 39352
rect 29420 39312 29426 39324
rect 29794 39321 29806 39324
rect 29840 39321 29852 39355
rect 32677 39355 32735 39361
rect 32677 39352 32689 39355
rect 29794 39315 29852 39321
rect 31956 39324 32689 39352
rect 31956 39296 31984 39324
rect 32677 39321 32689 39324
rect 32723 39321 32735 39355
rect 32677 39315 32735 39321
rect 43806 39312 43812 39364
rect 43864 39312 43870 39364
rect 16448 39256 17356 39284
rect 16448 39244 16454 39256
rect 17954 39244 17960 39296
rect 18012 39244 18018 39296
rect 18690 39244 18696 39296
rect 18748 39244 18754 39296
rect 21450 39244 21456 39296
rect 21508 39244 21514 39296
rect 22557 39287 22615 39293
rect 22557 39253 22569 39287
rect 22603 39284 22615 39287
rect 23198 39284 23204 39296
rect 22603 39256 23204 39284
rect 22603 39253 22615 39256
rect 22557 39247 22615 39253
rect 23198 39244 23204 39256
rect 23256 39244 23262 39296
rect 23382 39244 23388 39296
rect 23440 39284 23446 39296
rect 24029 39287 24087 39293
rect 24029 39284 24041 39287
rect 23440 39256 24041 39284
rect 23440 39244 23446 39256
rect 24029 39253 24041 39256
rect 24075 39253 24087 39287
rect 24029 39247 24087 39253
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 25041 39287 25099 39293
rect 25041 39284 25053 39287
rect 24360 39256 25053 39284
rect 24360 39244 24366 39256
rect 25041 39253 25053 39256
rect 25087 39253 25099 39287
rect 25041 39247 25099 39253
rect 25406 39244 25412 39296
rect 25464 39284 25470 39296
rect 25501 39287 25559 39293
rect 25501 39284 25513 39287
rect 25464 39256 25513 39284
rect 25464 39244 25470 39256
rect 25501 39253 25513 39256
rect 25547 39253 25559 39287
rect 25501 39247 25559 39253
rect 25869 39287 25927 39293
rect 25869 39253 25881 39287
rect 25915 39284 25927 39287
rect 26234 39284 26240 39296
rect 25915 39256 26240 39284
rect 25915 39253 25927 39256
rect 25869 39247 25927 39253
rect 26234 39244 26240 39256
rect 26292 39244 26298 39296
rect 27246 39244 27252 39296
rect 27304 39244 27310 39296
rect 27338 39244 27344 39296
rect 27396 39284 27402 39296
rect 27433 39287 27491 39293
rect 27433 39284 27445 39287
rect 27396 39256 27445 39284
rect 27396 39244 27402 39256
rect 27433 39253 27445 39256
rect 27479 39253 27491 39287
rect 27433 39247 27491 39253
rect 28258 39244 28264 39296
rect 28316 39284 28322 39296
rect 28905 39287 28963 39293
rect 28905 39284 28917 39287
rect 28316 39256 28917 39284
rect 28316 39244 28322 39256
rect 28905 39253 28917 39256
rect 28951 39253 28963 39287
rect 28905 39247 28963 39253
rect 29178 39244 29184 39296
rect 29236 39244 29242 39296
rect 30926 39244 30932 39296
rect 30984 39244 30990 39296
rect 31938 39244 31944 39296
rect 31996 39244 32002 39296
rect 32030 39244 32036 39296
rect 32088 39284 32094 39296
rect 32401 39287 32459 39293
rect 32401 39284 32413 39287
rect 32088 39256 32413 39284
rect 32088 39244 32094 39256
rect 32401 39253 32413 39256
rect 32447 39253 32459 39287
rect 32401 39247 32459 39253
rect 43530 39244 43536 39296
rect 43588 39244 43594 39296
rect 1104 39194 43884 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 43884 39194
rect 1104 39120 43884 39142
rect 5994 39040 6000 39092
rect 6052 39080 6058 39092
rect 6365 39083 6423 39089
rect 6365 39080 6377 39083
rect 6052 39052 6377 39080
rect 6052 39040 6058 39052
rect 6365 39049 6377 39052
rect 6411 39049 6423 39083
rect 6365 39043 6423 39049
rect 6733 39083 6791 39089
rect 6733 39049 6745 39083
rect 6779 39080 6791 39083
rect 7098 39080 7104 39092
rect 6779 39052 7104 39080
rect 6779 39049 6791 39052
rect 6733 39043 6791 39049
rect 7098 39040 7104 39052
rect 7156 39040 7162 39092
rect 8570 39040 8576 39092
rect 8628 39080 8634 39092
rect 8941 39083 8999 39089
rect 8941 39080 8953 39083
rect 8628 39052 8953 39080
rect 8628 39040 8634 39052
rect 8941 39049 8953 39052
rect 8987 39049 8999 39083
rect 8941 39043 8999 39049
rect 9401 39083 9459 39089
rect 9401 39049 9413 39083
rect 9447 39080 9459 39083
rect 9674 39080 9680 39092
rect 9447 39052 9680 39080
rect 9447 39049 9459 39052
rect 9401 39043 9459 39049
rect 9674 39040 9680 39052
rect 9732 39040 9738 39092
rect 11238 39040 11244 39092
rect 11296 39040 11302 39092
rect 11514 39040 11520 39092
rect 11572 39040 11578 39092
rect 11882 39040 11888 39092
rect 11940 39040 11946 39092
rect 12713 39083 12771 39089
rect 12713 39080 12725 39083
rect 11992 39052 12725 39080
rect 7828 39015 7886 39021
rect 7828 38981 7840 39015
rect 7874 39012 7886 39015
rect 8662 39012 8668 39024
rect 7874 38984 8668 39012
rect 7874 38981 7886 38984
rect 7828 38975 7886 38981
rect 8662 38972 8668 38984
rect 8720 38972 8726 39024
rect 9490 38972 9496 39024
rect 9548 38972 9554 39024
rect 10128 39015 10186 39021
rect 10128 38981 10140 39015
rect 10174 39012 10186 39015
rect 10962 39012 10968 39024
rect 10174 38984 10968 39012
rect 10174 38981 10186 38984
rect 10128 38975 10186 38981
rect 10962 38972 10968 38984
rect 11020 38972 11026 39024
rect 11532 39012 11560 39040
rect 11992 39012 12020 39052
rect 12713 39049 12725 39052
rect 12759 39049 12771 39083
rect 12713 39043 12771 39049
rect 13081 39083 13139 39089
rect 13081 39049 13093 39083
rect 13127 39080 13139 39083
rect 13814 39080 13820 39092
rect 13127 39052 13820 39080
rect 13127 39049 13139 39052
rect 13081 39043 13139 39049
rect 13814 39040 13820 39052
rect 13872 39040 13878 39092
rect 13909 39083 13967 39089
rect 13909 39049 13921 39083
rect 13955 39080 13967 39083
rect 14090 39080 14096 39092
rect 13955 39052 14096 39080
rect 13955 39049 13967 39052
rect 13909 39043 13967 39049
rect 14090 39040 14096 39052
rect 14148 39040 14154 39092
rect 15930 39040 15936 39092
rect 15988 39080 15994 39092
rect 16025 39083 16083 39089
rect 16025 39080 16037 39083
rect 15988 39052 16037 39080
rect 15988 39040 15994 39052
rect 16025 39049 16037 39052
rect 16071 39049 16083 39083
rect 16025 39043 16083 39049
rect 18138 39040 18144 39092
rect 18196 39040 18202 39092
rect 18322 39040 18328 39092
rect 18380 39080 18386 39092
rect 18509 39083 18567 39089
rect 18509 39080 18521 39083
rect 18380 39052 18521 39080
rect 18380 39040 18386 39052
rect 18509 39049 18521 39052
rect 18555 39049 18567 39083
rect 18509 39043 18567 39049
rect 18690 39040 18696 39092
rect 18748 39040 18754 39092
rect 23201 39083 23259 39089
rect 23201 39049 23213 39083
rect 23247 39080 23259 39083
rect 24394 39080 24400 39092
rect 23247 39052 24400 39080
rect 23247 39049 23259 39052
rect 23201 39043 23259 39049
rect 24394 39040 24400 39052
rect 24452 39040 24458 39092
rect 26513 39083 26571 39089
rect 26513 39049 26525 39083
rect 26559 39080 26571 39083
rect 27246 39080 27252 39092
rect 26559 39052 27252 39080
rect 26559 39049 26571 39052
rect 26513 39043 26571 39049
rect 27246 39040 27252 39052
rect 27304 39040 27310 39092
rect 27341 39083 27399 39089
rect 27341 39049 27353 39083
rect 27387 39049 27399 39083
rect 27341 39043 27399 39049
rect 28813 39083 28871 39089
rect 28813 39049 28825 39083
rect 28859 39080 28871 39083
rect 29270 39080 29276 39092
rect 28859 39052 29276 39080
rect 28859 39049 28871 39052
rect 28813 39043 28871 39049
rect 11532 38984 12020 39012
rect 12253 39015 12311 39021
rect 12253 38981 12265 39015
rect 12299 39012 12311 39015
rect 12986 39012 12992 39024
rect 12299 38984 12992 39012
rect 12299 38981 12311 38984
rect 12253 38975 12311 38981
rect 12986 38972 12992 38984
rect 13044 38972 13050 39024
rect 13170 38972 13176 39024
rect 13228 38972 13234 39024
rect 13538 38972 13544 39024
rect 13596 39012 13602 39024
rect 14001 39015 14059 39021
rect 14001 39012 14013 39015
rect 13596 38984 14013 39012
rect 13596 38972 13602 38984
rect 14001 38981 14013 38984
rect 14047 38981 14059 39015
rect 14001 38975 14059 38981
rect 14912 39015 14970 39021
rect 14912 38981 14924 39015
rect 14958 39012 14970 39015
rect 15010 39012 15016 39024
rect 14958 38984 15016 39012
rect 14958 38981 14970 38984
rect 14912 38975 14970 38981
rect 15010 38972 15016 38984
rect 15068 38972 15074 39024
rect 16936 39015 16994 39021
rect 16936 38981 16948 39015
rect 16982 39012 16994 39015
rect 18708 39012 18736 39040
rect 23474 39012 23480 39024
rect 16982 38984 18736 39012
rect 21376 38984 23480 39012
rect 16982 38981 16994 38984
rect 16936 38975 16994 38981
rect 13188 38944 13216 38972
rect 21376 38956 21404 38984
rect 23474 38972 23480 38984
rect 23532 38972 23538 39024
rect 24302 39012 24308 39024
rect 23584 38984 24308 39012
rect 7024 38916 9260 38944
rect 5626 38836 5632 38888
rect 5684 38836 5690 38888
rect 5902 38836 5908 38888
rect 5960 38876 5966 38888
rect 7024 38885 7052 38916
rect 9232 38888 9260 38916
rect 12360 38916 13216 38944
rect 12360 38888 12388 38916
rect 14642 38904 14648 38956
rect 14700 38904 14706 38956
rect 16669 38947 16727 38953
rect 16669 38913 16681 38947
rect 16715 38944 16727 38947
rect 17494 38944 17500 38956
rect 16715 38916 17500 38944
rect 16715 38913 16727 38916
rect 16669 38907 16727 38913
rect 17494 38904 17500 38916
rect 17552 38904 17558 38956
rect 17954 38904 17960 38956
rect 18012 38944 18018 38956
rect 18969 38947 19027 38953
rect 18969 38944 18981 38947
rect 18012 38916 18981 38944
rect 18012 38904 18018 38916
rect 18969 38913 18981 38916
rect 19015 38944 19027 38947
rect 19978 38944 19984 38956
rect 19015 38916 19984 38944
rect 19015 38913 19027 38916
rect 18969 38907 19027 38913
rect 19978 38904 19984 38916
rect 20036 38904 20042 38956
rect 21358 38904 21364 38956
rect 21416 38904 21422 38956
rect 21910 38904 21916 38956
rect 21968 38944 21974 38956
rect 23584 38953 23612 38984
rect 24302 38972 24308 38984
rect 24360 38972 24366 39024
rect 24486 38972 24492 39024
rect 24544 39012 24550 39024
rect 26878 39012 26884 39024
rect 24544 38984 26884 39012
rect 24544 38972 24550 38984
rect 22077 38947 22135 38953
rect 22077 38944 22089 38947
rect 21968 38916 22089 38944
rect 21968 38904 21974 38916
rect 22077 38913 22089 38916
rect 22123 38913 22135 38947
rect 22077 38907 22135 38913
rect 23569 38947 23627 38953
rect 23569 38913 23581 38947
rect 23615 38913 23627 38947
rect 23569 38907 23627 38913
rect 23661 38947 23719 38953
rect 23661 38913 23673 38947
rect 23707 38913 23719 38947
rect 23661 38907 23719 38913
rect 23845 38947 23903 38953
rect 23845 38913 23857 38947
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 6825 38879 6883 38885
rect 6825 38876 6837 38879
rect 5960 38848 6837 38876
rect 5960 38836 5966 38848
rect 6825 38845 6837 38848
rect 6871 38845 6883 38879
rect 6825 38839 6883 38845
rect 7009 38879 7067 38885
rect 7009 38845 7021 38879
rect 7055 38845 7067 38879
rect 7374 38876 7380 38888
rect 7009 38839 7067 38845
rect 7116 38848 7380 38876
rect 7116 38752 7144 38848
rect 7374 38836 7380 38848
rect 7432 38876 7438 38888
rect 7561 38879 7619 38885
rect 7561 38876 7573 38879
rect 7432 38848 7573 38876
rect 7432 38836 7438 38848
rect 7561 38845 7573 38848
rect 7607 38845 7619 38879
rect 7561 38839 7619 38845
rect 9214 38836 9220 38888
rect 9272 38836 9278 38888
rect 9490 38836 9496 38888
rect 9548 38876 9554 38888
rect 9585 38879 9643 38885
rect 9585 38876 9597 38879
rect 9548 38848 9597 38876
rect 9548 38836 9554 38848
rect 9585 38845 9597 38848
rect 9631 38845 9643 38879
rect 9585 38839 9643 38845
rect 9766 38836 9772 38888
rect 9824 38876 9830 38888
rect 9861 38879 9919 38885
rect 9861 38876 9873 38879
rect 9824 38848 9873 38876
rect 9824 38836 9830 38848
rect 9861 38845 9873 38848
rect 9907 38845 9919 38879
rect 9861 38839 9919 38845
rect 12342 38836 12348 38888
rect 12400 38836 12406 38888
rect 12437 38879 12495 38885
rect 12437 38845 12449 38879
rect 12483 38845 12495 38879
rect 12437 38839 12495 38845
rect 12452 38808 12480 38839
rect 13262 38836 13268 38888
rect 13320 38836 13326 38888
rect 14185 38879 14243 38885
rect 14185 38845 14197 38879
rect 14231 38876 14243 38879
rect 14274 38876 14280 38888
rect 14231 38848 14280 38876
rect 14231 38845 14243 38848
rect 14185 38839 14243 38845
rect 14274 38836 14280 38848
rect 14332 38836 14338 38888
rect 17678 38836 17684 38888
rect 17736 38876 17742 38888
rect 18601 38879 18659 38885
rect 18601 38876 18613 38879
rect 17736 38848 18613 38876
rect 17736 38836 17742 38848
rect 18601 38845 18613 38848
rect 18647 38845 18659 38879
rect 18601 38839 18659 38845
rect 18782 38836 18788 38888
rect 18840 38836 18846 38888
rect 21818 38836 21824 38888
rect 21876 38836 21882 38888
rect 23382 38876 23388 38888
rect 23032 38848 23388 38876
rect 12406 38780 14688 38808
rect 6178 38700 6184 38752
rect 6236 38700 6242 38752
rect 7098 38700 7104 38752
rect 7156 38700 7162 38752
rect 8202 38700 8208 38752
rect 8260 38740 8266 38752
rect 9033 38743 9091 38749
rect 9033 38740 9045 38743
rect 8260 38712 9045 38740
rect 8260 38700 8266 38712
rect 9033 38709 9045 38712
rect 9079 38709 9091 38743
rect 9033 38703 9091 38709
rect 11054 38700 11060 38752
rect 11112 38740 11118 38752
rect 12406 38740 12434 38780
rect 11112 38712 12434 38740
rect 11112 38700 11118 38712
rect 13354 38700 13360 38752
rect 13412 38740 13418 38752
rect 13541 38743 13599 38749
rect 13541 38740 13553 38743
rect 13412 38712 13553 38740
rect 13412 38700 13418 38712
rect 13541 38709 13553 38712
rect 13587 38709 13599 38743
rect 14660 38740 14688 38780
rect 15654 38740 15660 38752
rect 14660 38712 15660 38740
rect 13541 38703 13599 38709
rect 15654 38700 15660 38712
rect 15712 38700 15718 38752
rect 15838 38700 15844 38752
rect 15896 38740 15902 38752
rect 16390 38740 16396 38752
rect 15896 38712 16396 38740
rect 15896 38700 15902 38712
rect 16390 38700 16396 38712
rect 16448 38700 16454 38752
rect 17770 38700 17776 38752
rect 17828 38740 17834 38752
rect 18049 38743 18107 38749
rect 18049 38740 18061 38743
rect 17828 38712 18061 38740
rect 17828 38700 17834 38712
rect 18049 38709 18061 38712
rect 18095 38709 18107 38743
rect 18049 38703 18107 38709
rect 19610 38700 19616 38752
rect 19668 38700 19674 38752
rect 20254 38700 20260 38752
rect 20312 38700 20318 38752
rect 20438 38700 20444 38752
rect 20496 38740 20502 38752
rect 20533 38743 20591 38749
rect 20533 38740 20545 38743
rect 20496 38712 20545 38740
rect 20496 38700 20502 38712
rect 20533 38709 20545 38712
rect 20579 38709 20591 38743
rect 20533 38703 20591 38709
rect 21266 38700 21272 38752
rect 21324 38700 21330 38752
rect 21634 38700 21640 38752
rect 21692 38700 21698 38752
rect 22094 38700 22100 38752
rect 22152 38740 22158 38752
rect 23032 38740 23060 38848
rect 23382 38836 23388 38848
rect 23440 38876 23446 38888
rect 23676 38876 23704 38907
rect 23440 38848 23704 38876
rect 23860 38876 23888 38907
rect 24578 38904 24584 38956
rect 24636 38904 24642 38956
rect 24762 38904 24768 38956
rect 24820 38904 24826 38956
rect 25148 38953 25176 38984
rect 26878 38972 26884 38984
rect 26936 39012 26942 39024
rect 27356 39012 27384 39043
rect 29270 39040 29276 39052
rect 29328 39040 29334 39092
rect 29362 39040 29368 39092
rect 29420 39080 29426 39092
rect 29546 39080 29552 39092
rect 29420 39052 29552 39080
rect 29420 39040 29426 39052
rect 29546 39040 29552 39052
rect 29604 39040 29610 39092
rect 29638 39040 29644 39092
rect 29696 39040 29702 39092
rect 30926 39040 30932 39092
rect 30984 39080 30990 39092
rect 30984 39052 31754 39080
rect 30984 39040 30990 39052
rect 27678 39015 27736 39021
rect 27678 39012 27690 39015
rect 26936 38984 27292 39012
rect 27356 38984 27690 39012
rect 26936 38972 26942 38984
rect 27264 38956 27292 38984
rect 27678 38981 27690 38984
rect 27724 38981 27736 39015
rect 29656 39012 29684 39040
rect 27678 38975 27736 38981
rect 29288 38984 29684 39012
rect 31726 39012 31754 39052
rect 31726 38984 32168 39012
rect 25406 38953 25412 38956
rect 24857 38947 24915 38953
rect 24857 38913 24869 38947
rect 24903 38913 24915 38947
rect 24857 38907 24915 38913
rect 25133 38947 25191 38953
rect 25133 38913 25145 38947
rect 25179 38913 25191 38947
rect 25400 38944 25412 38953
rect 25367 38916 25412 38944
rect 25133 38907 25191 38913
rect 25400 38907 25412 38916
rect 23934 38876 23940 38888
rect 23860 38848 23940 38876
rect 23440 38836 23446 38848
rect 23934 38836 23940 38848
rect 23992 38876 23998 38888
rect 24210 38876 24216 38888
rect 23992 38848 24216 38876
rect 23992 38836 23998 38848
rect 24210 38836 24216 38848
rect 24268 38836 24274 38888
rect 24305 38879 24363 38885
rect 24305 38845 24317 38879
rect 24351 38845 24363 38879
rect 24305 38839 24363 38845
rect 24320 38808 24348 38839
rect 23216 38780 24348 38808
rect 23216 38752 23244 38780
rect 22152 38712 23060 38740
rect 22152 38700 22158 38712
rect 23198 38700 23204 38752
rect 23256 38700 23262 38752
rect 23474 38700 23480 38752
rect 23532 38740 23538 38752
rect 24397 38743 24455 38749
rect 24397 38740 24409 38743
rect 23532 38712 24409 38740
rect 23532 38700 23538 38712
rect 24397 38709 24409 38712
rect 24443 38709 24455 38743
rect 24872 38740 24900 38907
rect 25406 38904 25412 38907
rect 25464 38904 25470 38956
rect 25958 38904 25964 38956
rect 26016 38944 26022 38956
rect 26973 38947 27031 38953
rect 26973 38944 26985 38947
rect 26016 38916 26985 38944
rect 26016 38904 26022 38916
rect 26973 38913 26985 38916
rect 27019 38944 27031 38947
rect 27062 38944 27068 38956
rect 27019 38916 27068 38944
rect 27019 38913 27031 38916
rect 26973 38907 27031 38913
rect 27062 38904 27068 38916
rect 27120 38904 27126 38956
rect 27157 38947 27215 38953
rect 27157 38913 27169 38947
rect 27203 38913 27215 38947
rect 27157 38907 27215 38913
rect 25314 38740 25320 38752
rect 24872 38712 25320 38740
rect 24397 38703 24455 38709
rect 25314 38700 25320 38712
rect 25372 38700 25378 38752
rect 27172 38740 27200 38907
rect 27246 38904 27252 38956
rect 27304 38944 27310 38956
rect 27433 38947 27491 38953
rect 27433 38944 27445 38947
rect 27304 38916 27445 38944
rect 27304 38904 27310 38916
rect 27433 38913 27445 38916
rect 27479 38913 27491 38947
rect 27433 38907 27491 38913
rect 27522 38904 27528 38956
rect 27580 38944 27586 38956
rect 29288 38953 29316 38984
rect 29273 38947 29331 38953
rect 27580 38916 28948 38944
rect 27580 38904 27586 38916
rect 28810 38836 28816 38888
rect 28868 38836 28874 38888
rect 28828 38808 28856 38836
rect 28368 38780 28856 38808
rect 28920 38808 28948 38916
rect 29273 38913 29285 38947
rect 29319 38913 29331 38947
rect 29273 38907 29331 38913
rect 29362 38904 29368 38956
rect 29420 38904 29426 38956
rect 29457 38947 29515 38953
rect 29457 38913 29469 38947
rect 29503 38913 29515 38947
rect 29457 38907 29515 38913
rect 29181 38879 29239 38885
rect 29181 38845 29193 38879
rect 29227 38876 29239 38879
rect 29380 38876 29408 38904
rect 29227 38848 29408 38876
rect 29227 38845 29239 38848
rect 29181 38839 29239 38845
rect 29472 38808 29500 38907
rect 29638 38904 29644 38956
rect 29696 38944 29702 38956
rect 30009 38947 30067 38953
rect 30009 38944 30021 38947
rect 29696 38916 30021 38944
rect 29696 38904 29702 38916
rect 30009 38913 30021 38916
rect 30055 38913 30067 38947
rect 30009 38907 30067 38913
rect 31202 38904 31208 38956
rect 31260 38944 31266 38956
rect 31938 38944 31944 38956
rect 31260 38916 31944 38944
rect 31260 38904 31266 38916
rect 31938 38904 31944 38916
rect 31996 38904 32002 38956
rect 32140 38953 32168 38984
rect 32125 38947 32183 38953
rect 32125 38913 32137 38947
rect 32171 38913 32183 38947
rect 32125 38907 32183 38913
rect 29914 38836 29920 38888
rect 29972 38836 29978 38888
rect 31021 38879 31079 38885
rect 31021 38876 31033 38879
rect 30024 38848 31033 38876
rect 30024 38808 30052 38848
rect 31021 38845 31033 38848
rect 31067 38876 31079 38879
rect 31481 38879 31539 38885
rect 31481 38876 31493 38879
rect 31067 38848 31493 38876
rect 31067 38845 31079 38848
rect 31021 38839 31079 38845
rect 31404 38820 31432 38848
rect 31481 38845 31493 38848
rect 31527 38876 31539 38879
rect 31527 38848 33364 38876
rect 31527 38845 31539 38848
rect 31481 38839 31539 38845
rect 28920 38780 30052 38808
rect 30852 38780 31248 38808
rect 28368 38740 28396 38780
rect 30852 38752 30880 38780
rect 27172 38712 28396 38740
rect 29086 38700 29092 38752
rect 29144 38740 29150 38752
rect 30653 38743 30711 38749
rect 30653 38740 30665 38743
rect 29144 38712 30665 38740
rect 29144 38700 29150 38712
rect 30653 38709 30665 38712
rect 30699 38709 30711 38743
rect 30653 38703 30711 38709
rect 30834 38700 30840 38752
rect 30892 38700 30898 38752
rect 31220 38740 31248 38780
rect 31386 38768 31392 38820
rect 31444 38768 31450 38820
rect 31570 38768 31576 38820
rect 31628 38808 31634 38820
rect 33226 38808 33232 38820
rect 31628 38780 33232 38808
rect 31628 38768 31634 38780
rect 33226 38768 33232 38780
rect 33284 38768 33290 38820
rect 32769 38743 32827 38749
rect 32769 38740 32781 38743
rect 31220 38712 32781 38740
rect 32769 38709 32781 38712
rect 32815 38709 32827 38743
rect 32769 38703 32827 38709
rect 33137 38743 33195 38749
rect 33137 38709 33149 38743
rect 33183 38740 33195 38743
rect 33336 38740 33364 38848
rect 33594 38740 33600 38752
rect 33183 38712 33600 38740
rect 33183 38709 33195 38712
rect 33137 38703 33195 38709
rect 33594 38700 33600 38712
rect 33652 38700 33658 38752
rect 1104 38650 43884 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 43884 38650
rect 1104 38576 43884 38598
rect 3068 38508 6684 38536
rect 1210 38360 1216 38412
rect 1268 38400 1274 38412
rect 1857 38403 1915 38409
rect 1857 38400 1869 38403
rect 1268 38372 1869 38400
rect 1268 38360 1274 38372
rect 1857 38369 1869 38372
rect 1903 38369 1915 38403
rect 1857 38363 1915 38369
rect 3068 38341 3096 38508
rect 6656 38468 6684 38508
rect 6730 38496 6736 38548
rect 6788 38536 6794 38548
rect 6917 38539 6975 38545
rect 6917 38536 6929 38539
rect 6788 38508 6929 38536
rect 6788 38496 6794 38508
rect 6917 38505 6929 38508
rect 6963 38505 6975 38539
rect 10226 38536 10232 38548
rect 6917 38499 6975 38505
rect 7024 38508 10232 38536
rect 7024 38468 7052 38508
rect 10226 38496 10232 38508
rect 10284 38496 10290 38548
rect 10410 38496 10416 38548
rect 10468 38536 10474 38548
rect 10505 38539 10563 38545
rect 10505 38536 10517 38539
rect 10468 38508 10517 38536
rect 10468 38496 10474 38508
rect 10505 38505 10517 38508
rect 10551 38505 10563 38539
rect 11054 38536 11060 38548
rect 10505 38499 10563 38505
rect 10980 38508 11060 38536
rect 6656 38440 7052 38468
rect 9214 38428 9220 38480
rect 9272 38468 9278 38480
rect 10980 38468 11008 38508
rect 11054 38496 11060 38508
rect 11112 38536 11118 38548
rect 11112 38508 11192 38536
rect 11112 38496 11118 38508
rect 9272 38440 11008 38468
rect 9272 38428 9278 38440
rect 10778 38360 10784 38412
rect 10836 38400 10842 38412
rect 11164 38409 11192 38508
rect 12618 38496 12624 38548
rect 12676 38536 12682 38548
rect 13630 38536 13636 38548
rect 12676 38508 13636 38536
rect 12676 38496 12682 38508
rect 13630 38496 13636 38508
rect 13688 38496 13694 38548
rect 15102 38496 15108 38548
rect 15160 38536 15166 38548
rect 15197 38539 15255 38545
rect 15197 38536 15209 38539
rect 15160 38508 15209 38536
rect 15160 38496 15166 38508
rect 15197 38505 15209 38508
rect 15243 38505 15255 38539
rect 15197 38499 15255 38505
rect 16761 38539 16819 38545
rect 16761 38505 16773 38539
rect 16807 38536 16819 38539
rect 16850 38536 16856 38548
rect 16807 38508 16856 38536
rect 16807 38505 16819 38508
rect 16761 38499 16819 38505
rect 16850 38496 16856 38508
rect 16908 38496 16914 38548
rect 17589 38539 17647 38545
rect 17589 38505 17601 38539
rect 17635 38536 17647 38539
rect 17635 38508 17816 38536
rect 17635 38505 17647 38508
rect 17589 38499 17647 38505
rect 17788 38468 17816 38508
rect 17862 38496 17868 38548
rect 17920 38536 17926 38548
rect 17920 38508 20116 38536
rect 17920 38496 17926 38508
rect 20088 38468 20116 38508
rect 20162 38496 20168 38548
rect 20220 38496 20226 38548
rect 21174 38496 21180 38548
rect 21232 38536 21238 38548
rect 21269 38539 21327 38545
rect 21269 38536 21281 38539
rect 21232 38508 21281 38536
rect 21232 38496 21238 38508
rect 21269 38505 21281 38508
rect 21315 38505 21327 38539
rect 24578 38536 24584 38548
rect 21269 38499 21327 38505
rect 21928 38508 24584 38536
rect 20254 38468 20260 38480
rect 15856 38440 17623 38468
rect 17788 38440 19288 38468
rect 20088 38440 20260 38468
rect 10965 38403 11023 38409
rect 10965 38400 10977 38403
rect 10836 38372 10977 38400
rect 10836 38360 10842 38372
rect 10965 38369 10977 38372
rect 11011 38369 11023 38403
rect 10965 38363 11023 38369
rect 11149 38403 11207 38409
rect 11149 38369 11161 38403
rect 11195 38369 11207 38403
rect 11149 38363 11207 38369
rect 11974 38360 11980 38412
rect 12032 38400 12038 38412
rect 12250 38400 12256 38412
rect 12032 38372 12256 38400
rect 12032 38360 12038 38372
rect 12250 38360 12256 38372
rect 12308 38360 12314 38412
rect 14182 38360 14188 38412
rect 14240 38400 14246 38412
rect 15470 38400 15476 38412
rect 14240 38372 15476 38400
rect 14240 38360 14246 38372
rect 15470 38360 15476 38372
rect 15528 38400 15534 38412
rect 15856 38409 15884 38440
rect 15841 38403 15899 38409
rect 15841 38400 15853 38403
rect 15528 38372 15853 38400
rect 15528 38360 15534 38372
rect 15841 38369 15853 38372
rect 15887 38369 15899 38403
rect 15841 38363 15899 38369
rect 16022 38360 16028 38412
rect 16080 38360 16086 38412
rect 17405 38403 17463 38409
rect 17405 38369 17417 38403
rect 17451 38400 17463 38403
rect 17494 38400 17500 38412
rect 17451 38372 17500 38400
rect 17451 38369 17463 38372
rect 17405 38363 17463 38369
rect 17494 38360 17500 38372
rect 17552 38360 17558 38412
rect 17595 38400 17623 38440
rect 19260 38409 19288 38440
rect 20254 38428 20260 38440
rect 20312 38468 20318 38480
rect 20530 38468 20536 38480
rect 20312 38440 20536 38468
rect 20312 38428 20318 38440
rect 20530 38428 20536 38440
rect 20588 38428 20594 38480
rect 20809 38471 20867 38477
rect 20809 38437 20821 38471
rect 20855 38468 20867 38471
rect 21542 38468 21548 38480
rect 20855 38440 21548 38468
rect 20855 38437 20867 38440
rect 20809 38431 20867 38437
rect 21542 38428 21548 38440
rect 21600 38428 21606 38480
rect 21821 38471 21879 38477
rect 21821 38437 21833 38471
rect 21867 38468 21879 38471
rect 21928 38468 21956 38508
rect 24578 38496 24584 38508
rect 24636 38496 24642 38548
rect 29270 38536 29276 38548
rect 26896 38508 29276 38536
rect 23290 38468 23296 38480
rect 21867 38440 21956 38468
rect 22020 38440 23296 38468
rect 21867 38437 21879 38440
rect 21821 38431 21879 38437
rect 18141 38403 18199 38409
rect 18141 38400 18153 38403
rect 17595 38372 18153 38400
rect 18141 38369 18153 38372
rect 18187 38369 18199 38403
rect 19245 38403 19303 38409
rect 18141 38363 18199 38369
rect 18340 38372 18552 38400
rect 1581 38335 1639 38341
rect 1581 38301 1593 38335
rect 1627 38332 1639 38335
rect 3053 38335 3111 38341
rect 3053 38332 3065 38335
rect 1627 38304 3065 38332
rect 1627 38301 1639 38304
rect 1581 38295 1639 38301
rect 3053 38301 3065 38304
rect 3099 38301 3111 38335
rect 3053 38295 3111 38301
rect 4154 38292 4160 38344
rect 4212 38292 4218 38344
rect 4890 38292 4896 38344
rect 4948 38292 4954 38344
rect 5537 38335 5595 38341
rect 5537 38301 5549 38335
rect 5583 38332 5595 38335
rect 7009 38335 7067 38341
rect 7009 38332 7021 38335
rect 5583 38304 7021 38332
rect 5583 38301 5595 38304
rect 5537 38295 5595 38301
rect 7009 38301 7021 38304
rect 7055 38301 7067 38335
rect 7009 38295 7067 38301
rect 7276 38335 7334 38341
rect 7276 38301 7288 38335
rect 7322 38332 7334 38335
rect 7834 38332 7840 38344
rect 7322 38304 7840 38332
rect 7322 38301 7334 38304
rect 7276 38295 7334 38301
rect 5804 38267 5862 38273
rect 5804 38233 5816 38267
rect 5850 38264 5862 38267
rect 6546 38264 6552 38276
rect 5850 38236 6552 38264
rect 5850 38233 5862 38236
rect 5804 38227 5862 38233
rect 6546 38224 6552 38236
rect 6604 38224 6610 38276
rect 7024 38264 7052 38295
rect 7834 38292 7840 38304
rect 7892 38292 7898 38344
rect 9030 38292 9036 38344
rect 9088 38292 9094 38344
rect 9861 38335 9919 38341
rect 9861 38301 9873 38335
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 7098 38264 7104 38276
rect 7024 38236 7104 38264
rect 7098 38224 7104 38236
rect 7156 38264 7162 38276
rect 7466 38264 7472 38276
rect 7156 38236 7472 38264
rect 7156 38224 7162 38236
rect 7466 38224 7472 38236
rect 7524 38224 7530 38276
rect 9876 38264 9904 38295
rect 10870 38292 10876 38344
rect 10928 38292 10934 38344
rect 12526 38341 12532 38344
rect 11609 38335 11667 38341
rect 11609 38301 11621 38335
rect 11655 38301 11667 38335
rect 11609 38295 11667 38301
rect 12509 38335 12532 38341
rect 12509 38301 12521 38335
rect 12509 38295 12532 38301
rect 11054 38264 11060 38276
rect 9876 38236 11060 38264
rect 11054 38224 11060 38236
rect 11112 38224 11118 38276
rect 11624 38264 11652 38295
rect 12526 38292 12532 38295
rect 12584 38292 12590 38344
rect 13814 38292 13820 38344
rect 13872 38332 13878 38344
rect 14461 38335 14519 38341
rect 14461 38332 14473 38335
rect 13872 38304 14473 38332
rect 13872 38292 13878 38304
rect 14461 38301 14473 38304
rect 14507 38301 14519 38335
rect 14461 38295 14519 38301
rect 17129 38335 17187 38341
rect 17129 38301 17141 38335
rect 17175 38332 17187 38335
rect 18340 38332 18368 38372
rect 17175 38304 18368 38332
rect 17175 38301 17187 38304
rect 17129 38295 17187 38301
rect 14366 38264 14372 38276
rect 11624 38236 14372 38264
rect 14366 38224 14372 38236
rect 14424 38224 14430 38276
rect 14476 38264 14504 38295
rect 18414 38292 18420 38344
rect 18472 38292 18478 38344
rect 18524 38332 18552 38372
rect 19245 38369 19257 38403
rect 19291 38369 19303 38403
rect 19245 38363 19303 38369
rect 20714 38360 20720 38412
rect 20772 38360 20778 38412
rect 22020 38409 22048 38440
rect 23290 38428 23296 38440
rect 23348 38428 23354 38480
rect 20901 38403 20959 38409
rect 20901 38369 20913 38403
rect 20947 38400 20959 38403
rect 22005 38403 22063 38409
rect 20947 38372 21404 38400
rect 20947 38369 20959 38372
rect 20901 38363 20959 38369
rect 19610 38332 19616 38344
rect 18524 38304 19616 38332
rect 19610 38292 19616 38304
rect 19668 38292 19674 38344
rect 20732 38332 20760 38360
rect 21376 38344 21404 38372
rect 22005 38369 22017 38403
rect 22051 38369 22063 38403
rect 22005 38363 22063 38369
rect 22278 38360 22284 38412
rect 22336 38400 22342 38412
rect 23658 38400 23664 38412
rect 22336 38372 23664 38400
rect 22336 38360 22342 38372
rect 23658 38360 23664 38372
rect 23716 38400 23722 38412
rect 26896 38409 26924 38508
rect 29270 38496 29276 38508
rect 29328 38496 29334 38548
rect 31110 38536 31116 38548
rect 30852 38508 31116 38536
rect 27264 38440 28304 38468
rect 27264 38409 27292 38440
rect 28276 38412 28304 38440
rect 28718 38428 28724 38480
rect 28776 38468 28782 38480
rect 30852 38468 30880 38508
rect 31110 38496 31116 38508
rect 31168 38536 31174 38548
rect 31570 38536 31576 38548
rect 31168 38508 31576 38536
rect 31168 38496 31174 38508
rect 31570 38496 31576 38508
rect 31628 38496 31634 38548
rect 28776 38440 30880 38468
rect 28776 38428 28782 38440
rect 26881 38403 26939 38409
rect 26881 38400 26893 38403
rect 23716 38372 24164 38400
rect 23716 38360 23722 38372
rect 24136 38344 24164 38372
rect 25424 38372 26893 38400
rect 21085 38335 21143 38341
rect 21085 38332 21097 38335
rect 20732 38304 21097 38332
rect 21085 38301 21097 38304
rect 21131 38301 21143 38335
rect 21085 38295 21143 38301
rect 14826 38264 14832 38276
rect 14476 38236 14832 38264
rect 14826 38224 14832 38236
rect 14884 38224 14890 38276
rect 15565 38267 15623 38273
rect 15565 38233 15577 38267
rect 15611 38264 15623 38267
rect 16669 38267 16727 38273
rect 16669 38264 16681 38267
rect 15611 38236 16681 38264
rect 15611 38233 15623 38236
rect 15565 38227 15623 38233
rect 16669 38233 16681 38236
rect 16715 38233 16727 38267
rect 16669 38227 16727 38233
rect 16850 38224 16856 38276
rect 16908 38264 16914 38276
rect 17862 38264 17868 38276
rect 16908 38236 17868 38264
rect 16908 38224 16914 38236
rect 17862 38224 17868 38236
rect 17920 38224 17926 38276
rect 17957 38267 18015 38273
rect 17957 38233 17969 38267
rect 18003 38264 18015 38267
rect 19061 38267 19119 38273
rect 19061 38264 19073 38267
rect 18003 38236 19073 38264
rect 18003 38233 18015 38236
rect 17957 38227 18015 38233
rect 19061 38233 19073 38236
rect 19107 38233 19119 38267
rect 19061 38227 19119 38233
rect 19978 38224 19984 38276
rect 20036 38224 20042 38276
rect 4706 38156 4712 38208
rect 4764 38156 4770 38208
rect 5442 38156 5448 38208
rect 5500 38156 5506 38208
rect 6822 38156 6828 38208
rect 6880 38196 6886 38208
rect 8389 38199 8447 38205
rect 8389 38196 8401 38199
rect 6880 38168 8401 38196
rect 6880 38156 6886 38168
rect 8389 38165 8401 38168
rect 8435 38165 8447 38199
rect 8389 38159 8447 38165
rect 8754 38156 8760 38208
rect 8812 38156 8818 38208
rect 9674 38156 9680 38208
rect 9732 38156 9738 38208
rect 10410 38156 10416 38208
rect 10468 38156 10474 38208
rect 12161 38199 12219 38205
rect 12161 38165 12173 38199
rect 12207 38196 12219 38199
rect 12802 38196 12808 38208
rect 12207 38168 12808 38196
rect 12207 38165 12219 38168
rect 12161 38159 12219 38165
rect 12802 38156 12808 38168
rect 12860 38156 12866 38208
rect 15102 38156 15108 38208
rect 15160 38156 15166 38208
rect 15286 38156 15292 38208
rect 15344 38196 15350 38208
rect 15657 38199 15715 38205
rect 15657 38196 15669 38199
rect 15344 38168 15669 38196
rect 15344 38156 15350 38168
rect 15657 38165 15669 38168
rect 15703 38196 15715 38199
rect 17221 38199 17279 38205
rect 17221 38196 17233 38199
rect 15703 38168 17233 38196
rect 15703 38165 15715 38168
rect 15657 38159 15715 38165
rect 17221 38165 17233 38168
rect 17267 38196 17279 38199
rect 17678 38196 17684 38208
rect 17267 38168 17684 38196
rect 17267 38165 17279 38168
rect 17221 38159 17279 38165
rect 17678 38156 17684 38168
rect 17736 38156 17742 38208
rect 18049 38199 18107 38205
rect 18049 38165 18061 38199
rect 18095 38196 18107 38199
rect 18598 38196 18604 38208
rect 18095 38168 18604 38196
rect 18095 38165 18107 38168
rect 18049 38159 18107 38165
rect 18598 38156 18604 38168
rect 18656 38156 18662 38208
rect 18690 38156 18696 38208
rect 18748 38196 18754 38208
rect 19889 38199 19947 38205
rect 19889 38196 19901 38199
rect 18748 38168 19901 38196
rect 18748 38156 18754 38168
rect 19889 38165 19901 38168
rect 19935 38165 19947 38199
rect 19889 38159 19947 38165
rect 20070 38156 20076 38208
rect 20128 38196 20134 38208
rect 20181 38199 20239 38205
rect 20181 38196 20193 38199
rect 20128 38168 20193 38196
rect 20128 38156 20134 38168
rect 20181 38165 20193 38168
rect 20227 38165 20239 38199
rect 20181 38159 20239 38165
rect 20346 38156 20352 38208
rect 20404 38156 20410 38208
rect 21100 38196 21128 38295
rect 21358 38292 21364 38344
rect 21416 38292 21422 38344
rect 21545 38335 21603 38341
rect 21545 38301 21557 38335
rect 21591 38301 21603 38335
rect 21545 38295 21603 38301
rect 21266 38224 21272 38276
rect 21324 38264 21330 38276
rect 21560 38264 21588 38295
rect 21910 38292 21916 38344
rect 21968 38332 21974 38344
rect 22097 38335 22155 38341
rect 22097 38332 22109 38335
rect 21968 38304 22109 38332
rect 21968 38292 21974 38304
rect 22097 38301 22109 38304
rect 22143 38301 22155 38335
rect 22097 38295 22155 38301
rect 22186 38292 22192 38344
rect 22244 38292 22250 38344
rect 22465 38335 22523 38341
rect 22465 38301 22477 38335
rect 22511 38332 22523 38335
rect 23198 38332 23204 38344
rect 22511 38304 23204 38332
rect 22511 38301 22523 38304
rect 22465 38295 22523 38301
rect 23198 38292 23204 38304
rect 23256 38292 23262 38344
rect 23385 38335 23443 38341
rect 23385 38301 23397 38335
rect 23431 38332 23443 38335
rect 23474 38332 23480 38344
rect 23431 38304 23480 38332
rect 23431 38301 23443 38304
rect 23385 38295 23443 38301
rect 23474 38292 23480 38304
rect 23532 38292 23538 38344
rect 24118 38292 24124 38344
rect 24176 38292 24182 38344
rect 24397 38335 24455 38341
rect 24397 38301 24409 38335
rect 24443 38332 24455 38335
rect 24486 38332 24492 38344
rect 24443 38304 24492 38332
rect 24443 38301 24455 38304
rect 24397 38295 24455 38301
rect 24486 38292 24492 38304
rect 24544 38292 24550 38344
rect 25424 38276 25452 38372
rect 26881 38369 26893 38372
rect 26927 38369 26939 38403
rect 26881 38363 26939 38369
rect 27249 38403 27307 38409
rect 27249 38369 27261 38403
rect 27295 38369 27307 38403
rect 27249 38363 27307 38369
rect 28258 38360 28264 38412
rect 28316 38360 28322 38412
rect 28902 38360 28908 38412
rect 28960 38360 28966 38412
rect 29288 38409 29316 38440
rect 30926 38428 30932 38480
rect 30984 38468 30990 38480
rect 33689 38471 33747 38477
rect 33689 38468 33701 38471
rect 30984 38440 33701 38468
rect 30984 38428 30990 38440
rect 33689 38437 33701 38440
rect 33735 38437 33747 38471
rect 33689 38431 33747 38437
rect 29273 38403 29331 38409
rect 29273 38369 29285 38403
rect 29319 38369 29331 38403
rect 29273 38363 29331 38369
rect 29362 38360 29368 38412
rect 29420 38400 29426 38412
rect 30282 38400 30288 38412
rect 29420 38372 30288 38400
rect 29420 38360 29426 38372
rect 30282 38360 30288 38372
rect 30340 38400 30346 38412
rect 37642 38400 37648 38412
rect 30340 38372 30972 38400
rect 30340 38360 30346 38372
rect 30760 38344 30788 38372
rect 26142 38292 26148 38344
rect 26200 38292 26206 38344
rect 26237 38335 26295 38341
rect 26237 38301 26249 38335
rect 26283 38332 26295 38335
rect 26326 38332 26332 38344
rect 26283 38304 26332 38332
rect 26283 38301 26295 38304
rect 26237 38295 26295 38301
rect 26326 38292 26332 38304
rect 26384 38292 26390 38344
rect 26421 38335 26479 38341
rect 26421 38301 26433 38335
rect 26467 38301 26479 38335
rect 26421 38295 26479 38301
rect 21324 38236 21588 38264
rect 21729 38267 21787 38273
rect 21324 38224 21330 38236
rect 21729 38233 21741 38267
rect 21775 38264 21787 38267
rect 24642 38267 24700 38273
rect 24642 38264 24654 38267
rect 21775 38236 24654 38264
rect 21775 38233 21787 38236
rect 21729 38227 21787 38233
rect 24642 38233 24654 38236
rect 24688 38233 24700 38267
rect 24642 38227 24700 38233
rect 25406 38224 25412 38276
rect 25464 38224 25470 38276
rect 21450 38196 21456 38208
rect 21100 38168 21456 38196
rect 21450 38156 21456 38168
rect 21508 38196 21514 38208
rect 22695 38199 22753 38205
rect 22695 38196 22707 38199
rect 21508 38168 22707 38196
rect 21508 38156 21514 38168
rect 22695 38165 22707 38168
rect 22741 38165 22753 38199
rect 22695 38159 22753 38165
rect 24026 38156 24032 38208
rect 24084 38156 24090 38208
rect 25774 38156 25780 38208
rect 25832 38156 25838 38208
rect 26344 38196 26372 38292
rect 26436 38264 26464 38295
rect 26510 38292 26516 38344
rect 26568 38332 26574 38344
rect 27338 38332 27344 38344
rect 26568 38304 27344 38332
rect 26568 38292 26574 38304
rect 27338 38292 27344 38304
rect 27396 38292 27402 38344
rect 27522 38292 27528 38344
rect 27580 38292 27586 38344
rect 28074 38292 28080 38344
rect 28132 38332 28138 38344
rect 29178 38332 29184 38344
rect 28132 38304 29184 38332
rect 28132 38292 28138 38304
rect 29178 38292 29184 38304
rect 29236 38332 29242 38344
rect 29549 38335 29607 38341
rect 29549 38332 29561 38335
rect 29236 38304 29561 38332
rect 29236 38292 29242 38304
rect 29549 38301 29561 38304
rect 29595 38332 29607 38335
rect 29595 38304 30420 38332
rect 29595 38301 29607 38304
rect 29549 38295 29607 38301
rect 27540 38264 27568 38292
rect 26436 38236 27568 38264
rect 27982 38224 27988 38276
rect 28040 38224 28046 38276
rect 30006 38224 30012 38276
rect 30064 38264 30070 38276
rect 30285 38267 30343 38273
rect 30285 38264 30297 38267
rect 30064 38236 30297 38264
rect 30064 38224 30070 38236
rect 30285 38233 30297 38236
rect 30331 38233 30343 38267
rect 30392 38264 30420 38304
rect 30742 38292 30748 38344
rect 30800 38292 30806 38344
rect 30834 38292 30840 38344
rect 30892 38292 30898 38344
rect 30944 38341 30972 38372
rect 31726 38372 37648 38400
rect 30929 38335 30987 38341
rect 30929 38301 30941 38335
rect 30975 38301 30987 38335
rect 30929 38295 30987 38301
rect 31018 38292 31024 38344
rect 31076 38292 31082 38344
rect 31110 38292 31116 38344
rect 31168 38332 31174 38344
rect 31205 38335 31263 38341
rect 31205 38332 31217 38335
rect 31168 38304 31217 38332
rect 31168 38292 31174 38304
rect 31205 38301 31217 38304
rect 31251 38301 31263 38335
rect 31205 38295 31263 38301
rect 31573 38335 31631 38341
rect 31573 38301 31585 38335
rect 31619 38332 31631 38335
rect 31726 38332 31754 38372
rect 37642 38360 37648 38372
rect 37700 38360 37706 38412
rect 31619 38304 31754 38332
rect 31619 38301 31631 38304
rect 31573 38295 31631 38301
rect 32306 38292 32312 38344
rect 32364 38292 32370 38344
rect 32398 38292 32404 38344
rect 32456 38332 32462 38344
rect 33045 38335 33103 38341
rect 33045 38332 33057 38335
rect 32456 38304 33057 38332
rect 32456 38292 32462 38304
rect 33045 38301 33057 38304
rect 33091 38301 33103 38335
rect 33045 38295 33103 38301
rect 30392 38236 31892 38264
rect 30285 38227 30343 38233
rect 31864 38208 31892 38236
rect 31938 38224 31944 38276
rect 31996 38264 32002 38276
rect 32122 38264 32128 38276
rect 31996 38236 32128 38264
rect 31996 38224 32002 38236
rect 32122 38224 32128 38236
rect 32180 38224 32186 38276
rect 27154 38196 27160 38208
rect 26344 38168 27160 38196
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 30561 38199 30619 38205
rect 30561 38165 30573 38199
rect 30607 38196 30619 38199
rect 31754 38196 31760 38208
rect 30607 38168 31760 38196
rect 30607 38165 30619 38168
rect 30561 38159 30619 38165
rect 31754 38156 31760 38168
rect 31812 38156 31818 38208
rect 31846 38156 31852 38208
rect 31904 38156 31910 38208
rect 32950 38156 32956 38208
rect 33008 38156 33014 38208
rect 1104 38106 43884 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 43884 38106
rect 1104 38032 43884 38054
rect 4154 37952 4160 38004
rect 4212 37992 4218 38004
rect 4617 37995 4675 38001
rect 4617 37992 4629 37995
rect 4212 37964 4629 37992
rect 4212 37952 4218 37964
rect 4617 37961 4629 37964
rect 4663 37961 4675 37995
rect 4617 37955 4675 37961
rect 5626 37952 5632 38004
rect 5684 37952 5690 38004
rect 5813 37995 5871 38001
rect 5813 37961 5825 37995
rect 5859 37992 5871 37995
rect 6178 37992 6184 38004
rect 5859 37964 6184 37992
rect 5859 37961 5871 37964
rect 5813 37955 5871 37961
rect 6178 37952 6184 37964
rect 6236 37952 6242 38004
rect 6730 37952 6736 38004
rect 6788 37992 6794 38004
rect 6917 37995 6975 38001
rect 6917 37992 6929 37995
rect 6788 37964 6929 37992
rect 6788 37952 6794 37964
rect 6917 37961 6929 37964
rect 6963 37961 6975 37995
rect 9033 37995 9091 38001
rect 6917 37955 6975 37961
rect 7208 37964 8156 37992
rect 5644 37924 5672 37952
rect 6822 37924 6828 37936
rect 5644 37896 6828 37924
rect 6822 37884 6828 37896
rect 6880 37884 6886 37936
rect 4525 37859 4583 37865
rect 4525 37825 4537 37859
rect 4571 37856 4583 37859
rect 4985 37859 5043 37865
rect 4985 37856 4997 37859
rect 4571 37828 4997 37856
rect 4571 37825 4583 37828
rect 4525 37819 4583 37825
rect 4985 37825 4997 37828
rect 5031 37825 5043 37859
rect 4985 37819 5043 37825
rect 5077 37859 5135 37865
rect 5077 37825 5089 37859
rect 5123 37856 5135 37859
rect 7208 37856 7236 37964
rect 8128 37936 8156 37964
rect 9033 37961 9045 37995
rect 9079 37992 9091 37995
rect 9306 37992 9312 38004
rect 9079 37964 9312 37992
rect 9079 37961 9091 37964
rect 9033 37955 9091 37961
rect 9306 37952 9312 37964
rect 9364 37952 9370 38004
rect 9493 37995 9551 38001
rect 9493 37961 9505 37995
rect 9539 37992 9551 37995
rect 9582 37992 9588 38004
rect 9539 37964 9588 37992
rect 9539 37961 9551 37964
rect 9493 37955 9551 37961
rect 9582 37952 9588 37964
rect 9640 37952 9646 38004
rect 10410 37952 10416 38004
rect 10468 37992 10474 38004
rect 10781 37995 10839 38001
rect 10781 37992 10793 37995
rect 10468 37964 10793 37992
rect 10468 37952 10474 37964
rect 10781 37961 10793 37964
rect 10827 37961 10839 37995
rect 10781 37955 10839 37961
rect 11238 37952 11244 38004
rect 11296 37992 11302 38004
rect 11885 37995 11943 38001
rect 11885 37992 11897 37995
rect 11296 37964 11897 37992
rect 11296 37952 11302 37964
rect 11885 37961 11897 37964
rect 11931 37961 11943 37995
rect 15657 37995 15715 38001
rect 11885 37955 11943 37961
rect 12452 37964 15047 37992
rect 7920 37927 7978 37933
rect 7920 37893 7932 37927
rect 7966 37924 7978 37927
rect 8018 37924 8024 37936
rect 7966 37896 8024 37924
rect 7966 37893 7978 37896
rect 7920 37887 7978 37893
rect 8018 37884 8024 37896
rect 8076 37884 8082 37936
rect 8110 37884 8116 37936
rect 8168 37884 8174 37936
rect 5123 37828 5948 37856
rect 5123 37825 5135 37828
rect 5077 37819 5135 37825
rect 5920 37800 5948 37828
rect 7024 37828 7236 37856
rect 7561 37859 7619 37865
rect 7024 37800 7052 37828
rect 7561 37825 7573 37859
rect 7607 37856 7619 37859
rect 8294 37856 8300 37868
rect 7607 37828 8300 37856
rect 7607 37825 7619 37828
rect 7561 37819 7619 37825
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 10778 37816 10784 37868
rect 10836 37856 10842 37868
rect 10873 37859 10931 37865
rect 10873 37856 10885 37859
rect 10836 37828 10885 37856
rect 10836 37816 10842 37828
rect 10873 37825 10885 37828
rect 10919 37856 10931 37859
rect 11790 37856 11796 37868
rect 10919 37828 11796 37856
rect 10919 37825 10931 37828
rect 10873 37819 10931 37825
rect 11790 37816 11796 37828
rect 11848 37816 11854 37868
rect 12452 37865 12480 37964
rect 14642 37924 14648 37936
rect 12728 37896 14648 37924
rect 12437 37859 12495 37865
rect 12437 37856 12449 37859
rect 12176 37828 12449 37856
rect 12176 37800 12204 37828
rect 12437 37825 12449 37828
rect 12483 37825 12495 37859
rect 12437 37819 12495 37825
rect 12618 37816 12624 37868
rect 12676 37816 12682 37868
rect 3973 37791 4031 37797
rect 3973 37757 3985 37791
rect 4019 37757 4031 37791
rect 3973 37751 4031 37757
rect 3988 37720 4016 37751
rect 5258 37748 5264 37800
rect 5316 37788 5322 37800
rect 5316 37760 5856 37788
rect 5316 37748 5322 37760
rect 5626 37720 5632 37732
rect 3988 37692 5632 37720
rect 5626 37680 5632 37692
rect 5684 37680 5690 37732
rect 5828 37720 5856 37760
rect 5902 37748 5908 37800
rect 5960 37748 5966 37800
rect 6089 37791 6147 37797
rect 6089 37757 6101 37791
rect 6135 37788 6147 37791
rect 6362 37788 6368 37800
rect 6135 37760 6368 37788
rect 6135 37757 6147 37760
rect 6089 37751 6147 37757
rect 6362 37748 6368 37760
rect 6420 37788 6426 37800
rect 6914 37788 6920 37800
rect 6420 37760 6920 37788
rect 6420 37748 6426 37760
rect 6914 37748 6920 37760
rect 6972 37748 6978 37800
rect 7006 37748 7012 37800
rect 7064 37748 7070 37800
rect 7466 37748 7472 37800
rect 7524 37788 7530 37800
rect 7653 37791 7711 37797
rect 7653 37788 7665 37791
rect 7524 37760 7665 37788
rect 7524 37748 7530 37760
rect 7653 37757 7665 37760
rect 7699 37757 7711 37791
rect 7653 37751 7711 37757
rect 8938 37748 8944 37800
rect 8996 37748 9002 37800
rect 9398 37748 9404 37800
rect 9456 37788 9462 37800
rect 9585 37791 9643 37797
rect 9585 37788 9597 37791
rect 9456 37760 9597 37788
rect 9456 37748 9462 37760
rect 9585 37757 9597 37760
rect 9631 37757 9643 37791
rect 9585 37751 9643 37757
rect 9769 37791 9827 37797
rect 9769 37757 9781 37791
rect 9815 37788 9827 37791
rect 9815 37760 10640 37788
rect 9815 37757 9827 37760
rect 9769 37751 9827 37757
rect 8956 37720 8984 37748
rect 9125 37723 9183 37729
rect 9125 37720 9137 37723
rect 5828 37692 6592 37720
rect 8956 37692 9137 37720
rect 5445 37655 5503 37661
rect 5445 37621 5457 37655
rect 5491 37652 5503 37655
rect 6270 37652 6276 37664
rect 5491 37624 6276 37652
rect 5491 37621 5503 37624
rect 5445 37615 5503 37621
rect 6270 37612 6276 37624
rect 6328 37612 6334 37664
rect 6454 37612 6460 37664
rect 6512 37612 6518 37664
rect 6564 37652 6592 37692
rect 9125 37689 9137 37692
rect 9171 37689 9183 37723
rect 9125 37683 9183 37689
rect 9784 37652 9812 37751
rect 10612 37720 10640 37760
rect 10962 37748 10968 37800
rect 11020 37748 11026 37800
rect 11146 37748 11152 37800
rect 11204 37788 11210 37800
rect 11977 37791 12035 37797
rect 11977 37788 11989 37791
rect 11204 37760 11989 37788
rect 11204 37748 11210 37760
rect 11977 37757 11989 37760
rect 12023 37757 12035 37791
rect 11977 37751 12035 37757
rect 12158 37748 12164 37800
rect 12216 37748 12222 37800
rect 12728 37797 12756 37896
rect 14642 37884 14648 37896
rect 14700 37884 14706 37936
rect 12802 37816 12808 37868
rect 12860 37856 12866 37868
rect 12969 37859 13027 37865
rect 12969 37856 12981 37859
rect 12860 37828 12981 37856
rect 12860 37816 12866 37828
rect 12969 37825 12981 37828
rect 13015 37825 13027 37859
rect 12969 37819 13027 37825
rect 14553 37859 14611 37865
rect 14553 37825 14565 37859
rect 14599 37856 14611 37859
rect 14918 37856 14924 37868
rect 14599 37828 14924 37856
rect 14599 37825 14611 37828
rect 14553 37819 14611 37825
rect 14918 37816 14924 37828
rect 14976 37816 14982 37868
rect 15019 37856 15047 37964
rect 15657 37961 15669 37995
rect 15703 37992 15715 37995
rect 16022 37992 16028 38004
rect 15703 37964 16028 37992
rect 15703 37961 15715 37964
rect 15657 37955 15715 37961
rect 16022 37952 16028 37964
rect 16080 37952 16086 38004
rect 16206 37952 16212 38004
rect 16264 37992 16270 38004
rect 16264 37964 17540 37992
rect 16264 37952 16270 37964
rect 15102 37884 15108 37936
rect 15160 37924 15166 37936
rect 16945 37927 17003 37933
rect 16945 37924 16957 37927
rect 15160 37896 16957 37924
rect 15160 37884 15166 37896
rect 16945 37893 16957 37896
rect 16991 37893 17003 37927
rect 16945 37887 17003 37893
rect 15378 37856 15384 37868
rect 15019 37828 15384 37856
rect 15378 37816 15384 37828
rect 15436 37816 15442 37868
rect 15565 37859 15623 37865
rect 15565 37825 15577 37859
rect 15611 37856 15623 37859
rect 15930 37856 15936 37868
rect 15611 37828 15936 37856
rect 15611 37825 15623 37828
rect 15565 37819 15623 37825
rect 15930 37816 15936 37828
rect 15988 37816 15994 37868
rect 16117 37859 16175 37865
rect 16117 37825 16129 37859
rect 16163 37825 16175 37859
rect 16117 37819 16175 37825
rect 12713 37791 12771 37797
rect 12713 37757 12725 37791
rect 12759 37757 12771 37791
rect 12713 37751 12771 37757
rect 10612 37692 11468 37720
rect 11440 37664 11468 37692
rect 12250 37680 12256 37732
rect 12308 37720 12314 37732
rect 12728 37720 12756 37751
rect 15746 37748 15752 37800
rect 15804 37748 15810 37800
rect 16132 37788 16160 37819
rect 16206 37816 16212 37868
rect 16264 37816 16270 37868
rect 16669 37859 16727 37865
rect 16669 37825 16681 37859
rect 16715 37825 16727 37859
rect 16669 37819 16727 37825
rect 16853 37859 16911 37865
rect 16853 37825 16865 37859
rect 16899 37825 16911 37859
rect 16853 37819 16911 37825
rect 16390 37788 16396 37800
rect 16132 37760 16396 37788
rect 16390 37748 16396 37760
rect 16448 37748 16454 37800
rect 12308 37692 12756 37720
rect 12308 37680 12314 37692
rect 14458 37680 14464 37732
rect 14516 37720 14522 37732
rect 16684 37720 16712 37819
rect 16868 37788 16896 37819
rect 17034 37816 17040 37868
rect 17092 37816 17098 37868
rect 17126 37816 17132 37868
rect 17184 37856 17190 37868
rect 17313 37859 17371 37865
rect 17313 37856 17325 37859
rect 17184 37828 17325 37856
rect 17184 37816 17190 37828
rect 17313 37825 17325 37828
rect 17359 37825 17371 37859
rect 17512 37856 17540 37964
rect 18322 37952 18328 38004
rect 18380 37992 18386 38004
rect 18380 37964 20208 37992
rect 18380 37952 18386 37964
rect 17580 37927 17638 37933
rect 17580 37893 17592 37927
rect 17626 37924 17638 37927
rect 18690 37924 18696 37936
rect 17626 37896 18696 37924
rect 17626 37893 17638 37896
rect 17580 37887 17638 37893
rect 18690 37884 18696 37896
rect 18748 37884 18754 37936
rect 19426 37924 19432 37936
rect 18800 37896 19432 37924
rect 18800 37856 18828 37896
rect 19426 37884 19432 37896
rect 19484 37924 19490 37936
rect 20070 37924 20076 37936
rect 19484 37896 20076 37924
rect 19484 37884 19490 37896
rect 20070 37884 20076 37896
rect 20128 37884 20134 37936
rect 20180 37924 20208 37964
rect 20714 37952 20720 38004
rect 20772 37992 20778 38004
rect 22370 37992 22376 38004
rect 20772 37964 22376 37992
rect 20772 37952 20778 37964
rect 22370 37952 22376 37964
rect 22428 37952 22434 38004
rect 24026 37952 24032 38004
rect 24084 37952 24090 38004
rect 24854 37992 24860 38004
rect 24780 37964 24860 37992
rect 22732 37927 22790 37933
rect 20180 37896 22692 37924
rect 17512 37828 18828 37856
rect 17313 37819 17371 37825
rect 19242 37816 19248 37868
rect 19300 37856 19306 37868
rect 19705 37859 19763 37865
rect 19705 37856 19717 37859
rect 19300 37828 19717 37856
rect 19300 37816 19306 37828
rect 19705 37825 19717 37828
rect 19751 37825 19763 37859
rect 19705 37819 19763 37825
rect 19889 37859 19947 37865
rect 19889 37825 19901 37859
rect 19935 37825 19947 37859
rect 19889 37819 19947 37825
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37856 20039 37859
rect 20088 37856 20116 37884
rect 20027 37828 20116 37856
rect 20027 37825 20039 37828
rect 19981 37819 20039 37825
rect 16942 37788 16948 37800
rect 16868 37760 16948 37788
rect 16942 37748 16948 37760
rect 17000 37748 17006 37800
rect 18414 37748 18420 37800
rect 18472 37788 18478 37800
rect 18785 37791 18843 37797
rect 18785 37788 18797 37791
rect 18472 37760 18797 37788
rect 18472 37748 18478 37760
rect 18785 37757 18797 37760
rect 18831 37757 18843 37791
rect 18785 37751 18843 37757
rect 18874 37748 18880 37800
rect 18932 37788 18938 37800
rect 19904 37788 19932 37819
rect 20162 37816 20168 37868
rect 20220 37816 20226 37868
rect 20441 37859 20499 37865
rect 20441 37825 20453 37859
rect 20487 37856 20499 37859
rect 20530 37856 20536 37868
rect 20487 37828 20536 37856
rect 20487 37825 20499 37828
rect 20441 37819 20499 37825
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 20714 37816 20720 37868
rect 20772 37816 20778 37868
rect 20809 37859 20867 37865
rect 20809 37825 20821 37859
rect 20855 37825 20867 37859
rect 20809 37819 20867 37825
rect 20901 37859 20959 37865
rect 20901 37825 20913 37859
rect 20947 37856 20959 37859
rect 22554 37856 22560 37868
rect 20947 37828 22560 37856
rect 20947 37825 20959 37828
rect 20901 37819 20959 37825
rect 20180 37788 20208 37816
rect 18932 37760 19847 37788
rect 19904 37760 20208 37788
rect 20257 37791 20315 37797
rect 18932 37748 18938 37760
rect 14516 37692 16712 37720
rect 14516 37680 14522 37692
rect 17218 37680 17224 37732
rect 17276 37680 17282 37732
rect 18322 37680 18328 37732
rect 18380 37720 18386 37732
rect 19521 37723 19579 37729
rect 19521 37720 19533 37723
rect 18380 37692 19533 37720
rect 18380 37680 18386 37692
rect 19521 37689 19533 37692
rect 19567 37689 19579 37723
rect 19819 37720 19847 37760
rect 20257 37757 20269 37791
rect 20303 37788 20315 37791
rect 20732 37788 20760 37816
rect 20303 37760 20760 37788
rect 20824 37788 20852 37819
rect 22554 37816 22560 37828
rect 22612 37816 22618 37868
rect 22664 37856 22692 37896
rect 22732 37893 22744 37927
rect 22778 37924 22790 37927
rect 24044 37924 24072 37952
rect 22778 37896 24072 37924
rect 22778 37893 22790 37896
rect 22732 37887 22790 37893
rect 24780 37856 24808 37964
rect 24854 37952 24860 37964
rect 24912 37952 24918 38004
rect 25774 37952 25780 38004
rect 25832 37952 25838 38004
rect 26053 37995 26111 38001
rect 26053 37961 26065 37995
rect 26099 37992 26111 37995
rect 26142 37992 26148 38004
rect 26099 37964 26148 37992
rect 26099 37961 26111 37964
rect 26053 37955 26111 37961
rect 26142 37952 26148 37964
rect 26200 37952 26206 38004
rect 28810 37952 28816 38004
rect 28868 37952 28874 38004
rect 29638 37952 29644 38004
rect 29696 37952 29702 38004
rect 30009 37995 30067 38001
rect 30009 37961 30021 37995
rect 30055 37992 30067 37995
rect 31573 37995 31631 38001
rect 30055 37964 30512 37992
rect 30055 37961 30067 37964
rect 30009 37955 30067 37961
rect 25225 37927 25283 37933
rect 25225 37924 25237 37927
rect 24872 37896 25237 37924
rect 24872 37868 24900 37896
rect 25225 37893 25237 37896
rect 25271 37893 25283 37927
rect 25225 37887 25283 37893
rect 22664 37828 24808 37856
rect 24854 37816 24860 37868
rect 24912 37816 24918 37868
rect 25038 37816 25044 37868
rect 25096 37816 25102 37868
rect 25314 37816 25320 37868
rect 25372 37816 25378 37868
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37856 25559 37859
rect 25792 37856 25820 37952
rect 28442 37884 28448 37936
rect 28500 37924 28506 37936
rect 30024 37924 30052 37955
rect 28500 37896 30052 37924
rect 30484 37924 30512 37964
rect 31573 37961 31585 37995
rect 31619 37992 31631 37995
rect 32398 37992 32404 38004
rect 31619 37964 32404 37992
rect 31619 37961 31631 37964
rect 31573 37955 31631 37961
rect 32398 37952 32404 37964
rect 32456 37952 32462 38004
rect 32950 37952 32956 38004
rect 33008 37952 33014 38004
rect 33502 37952 33508 38004
rect 33560 37952 33566 38004
rect 32968 37924 32996 37952
rect 34241 37927 34299 37933
rect 34241 37924 34253 37927
rect 30484 37896 32996 37924
rect 33336 37896 34253 37924
rect 28500 37884 28506 37896
rect 25547 37828 25820 37856
rect 25547 37825 25559 37828
rect 25501 37819 25559 37825
rect 27430 37816 27436 37868
rect 27488 37816 27494 37868
rect 27522 37816 27528 37868
rect 27580 37816 27586 37868
rect 27700 37859 27758 37865
rect 27700 37825 27712 37859
rect 27746 37856 27758 37859
rect 29086 37856 29092 37868
rect 27746 37828 29092 37856
rect 27746 37825 27758 37828
rect 27700 37819 27758 37825
rect 29086 37816 29092 37828
rect 29144 37816 29150 37868
rect 29454 37816 29460 37868
rect 29512 37856 29518 37868
rect 29825 37859 29883 37865
rect 29825 37856 29837 37859
rect 29512 37828 29837 37856
rect 29512 37816 29518 37828
rect 29825 37825 29837 37828
rect 29871 37825 29883 37859
rect 29825 37819 29883 37825
rect 30101 37859 30159 37865
rect 30101 37825 30113 37859
rect 30147 37856 30159 37859
rect 30282 37856 30288 37868
rect 30147 37828 30288 37856
rect 30147 37825 30159 37828
rect 30101 37819 30159 37825
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 30466 37865 30472 37868
rect 30460 37856 30472 37865
rect 30427 37828 30472 37856
rect 30460 37819 30472 37828
rect 30466 37816 30472 37819
rect 30524 37816 30530 37868
rect 33134 37816 33140 37868
rect 33192 37856 33198 37868
rect 33336 37865 33364 37896
rect 34241 37893 34253 37896
rect 34287 37893 34299 37927
rect 34241 37887 34299 37893
rect 33321 37859 33379 37865
rect 33321 37856 33333 37859
rect 33192 37828 33333 37856
rect 33192 37816 33198 37828
rect 33321 37825 33333 37828
rect 33367 37825 33379 37859
rect 33781 37859 33839 37865
rect 33781 37856 33793 37859
rect 33321 37819 33379 37825
rect 33428 37828 33793 37856
rect 21358 37788 21364 37800
rect 20824 37760 21364 37788
rect 20303 37757 20315 37760
rect 20257 37751 20315 37757
rect 21358 37748 21364 37760
rect 21416 37748 21422 37800
rect 21818 37748 21824 37800
rect 21876 37788 21882 37800
rect 22094 37788 22100 37800
rect 21876 37760 22100 37788
rect 21876 37748 21882 37760
rect 22094 37748 22100 37760
rect 22152 37788 22158 37800
rect 22465 37791 22523 37797
rect 22465 37788 22477 37791
rect 22152 37760 22477 37788
rect 22152 37748 22158 37760
rect 22465 37757 22477 37760
rect 22511 37757 22523 37791
rect 24121 37791 24179 37797
rect 24121 37788 24133 37791
rect 22465 37751 22523 37757
rect 23860 37760 24133 37788
rect 19819 37692 20760 37720
rect 19521 37683 19579 37689
rect 6564 37624 9812 37652
rect 9858 37612 9864 37664
rect 9916 37652 9922 37664
rect 10229 37655 10287 37661
rect 10229 37652 10241 37655
rect 9916 37624 10241 37652
rect 9916 37612 9922 37624
rect 10229 37621 10241 37624
rect 10275 37621 10287 37655
rect 10229 37615 10287 37621
rect 10410 37612 10416 37664
rect 10468 37612 10474 37664
rect 11422 37612 11428 37664
rect 11480 37612 11486 37664
rect 11514 37612 11520 37664
rect 11572 37612 11578 37664
rect 12529 37655 12587 37661
rect 12529 37621 12541 37655
rect 12575 37652 12587 37655
rect 13630 37652 13636 37664
rect 12575 37624 13636 37652
rect 12575 37621 12587 37624
rect 12529 37615 12587 37621
rect 13630 37612 13636 37624
rect 13688 37612 13694 37664
rect 14090 37612 14096 37664
rect 14148 37612 14154 37664
rect 14918 37612 14924 37664
rect 14976 37652 14982 37664
rect 15105 37655 15163 37661
rect 15105 37652 15117 37655
rect 14976 37624 15117 37652
rect 14976 37612 14982 37624
rect 15105 37621 15117 37624
rect 15151 37621 15163 37655
rect 15105 37615 15163 37621
rect 15194 37612 15200 37664
rect 15252 37612 15258 37664
rect 15378 37612 15384 37664
rect 15436 37652 15442 37664
rect 16393 37655 16451 37661
rect 16393 37652 16405 37655
rect 15436 37624 16405 37652
rect 15436 37612 15442 37624
rect 16393 37621 16405 37624
rect 16439 37652 16451 37655
rect 16482 37652 16488 37664
rect 16439 37624 16488 37652
rect 16439 37621 16451 37624
rect 16393 37615 16451 37621
rect 16482 37612 16488 37624
rect 16540 37612 16546 37664
rect 16666 37612 16672 37664
rect 16724 37652 16730 37664
rect 18506 37652 18512 37664
rect 16724 37624 18512 37652
rect 16724 37612 16730 37624
rect 18506 37612 18512 37624
rect 18564 37652 18570 37664
rect 18693 37655 18751 37661
rect 18693 37652 18705 37655
rect 18564 37624 18705 37652
rect 18564 37612 18570 37624
rect 18693 37621 18705 37624
rect 18739 37621 18751 37655
rect 18693 37615 18751 37621
rect 18782 37612 18788 37664
rect 18840 37652 18846 37664
rect 19429 37655 19487 37661
rect 19429 37652 19441 37655
rect 18840 37624 19441 37652
rect 18840 37612 18846 37624
rect 19429 37621 19441 37624
rect 19475 37621 19487 37655
rect 19429 37615 19487 37621
rect 20530 37612 20536 37664
rect 20588 37652 20594 37664
rect 20625 37655 20683 37661
rect 20625 37652 20637 37655
rect 20588 37624 20637 37652
rect 20588 37612 20594 37624
rect 20625 37621 20637 37624
rect 20671 37621 20683 37655
rect 20732 37652 20760 37692
rect 20806 37680 20812 37732
rect 20864 37720 20870 37732
rect 22186 37720 22192 37732
rect 20864 37692 22192 37720
rect 20864 37680 20870 37692
rect 22186 37680 22192 37692
rect 22244 37720 22250 37732
rect 23860 37729 23888 37760
rect 24121 37757 24133 37760
rect 24167 37757 24179 37791
rect 25332 37788 25360 37816
rect 25774 37788 25780 37800
rect 25332 37760 25780 37788
rect 24121 37751 24179 37757
rect 25774 37748 25780 37760
rect 25832 37748 25838 37800
rect 26237 37791 26295 37797
rect 26237 37757 26249 37791
rect 26283 37757 26295 37791
rect 26237 37751 26295 37757
rect 22373 37723 22431 37729
rect 22373 37720 22385 37723
rect 22244 37692 22385 37720
rect 22244 37680 22250 37692
rect 22373 37689 22385 37692
rect 22419 37689 22431 37723
rect 22373 37683 22431 37689
rect 23845 37723 23903 37729
rect 23845 37689 23857 37723
rect 23891 37689 23903 37723
rect 23845 37683 23903 37689
rect 24210 37680 24216 37732
rect 24268 37720 24274 37732
rect 24857 37723 24915 37729
rect 24857 37720 24869 37723
rect 24268 37692 24869 37720
rect 24268 37680 24274 37692
rect 24857 37689 24869 37692
rect 24903 37689 24915 37723
rect 26252 37720 26280 37751
rect 26326 37748 26332 37800
rect 26384 37788 26390 37800
rect 27249 37791 27307 37797
rect 27249 37788 27261 37791
rect 26384 37760 27261 37788
rect 26384 37748 26390 37760
rect 27249 37757 27261 37760
rect 27295 37788 27307 37791
rect 27540 37788 27568 37816
rect 27295 37760 27568 37788
rect 27295 37757 27307 37760
rect 27249 37751 27307 37757
rect 28902 37748 28908 37800
rect 28960 37748 28966 37800
rect 30193 37791 30251 37797
rect 30193 37788 30205 37791
rect 30024 37760 30205 37788
rect 26252 37692 27476 37720
rect 24857 37683 24915 37689
rect 21266 37652 21272 37664
rect 20732 37624 21272 37652
rect 20625 37615 20683 37621
rect 21266 37612 21272 37624
rect 21324 37612 21330 37664
rect 21542 37612 21548 37664
rect 21600 37612 21606 37664
rect 23750 37612 23756 37664
rect 23808 37652 23814 37664
rect 24762 37652 24768 37664
rect 23808 37624 24768 37652
rect 23808 37612 23814 37624
rect 24762 37612 24768 37624
rect 24820 37612 24826 37664
rect 25222 37612 25228 37664
rect 25280 37652 25286 37664
rect 26234 37652 26240 37664
rect 25280 37624 26240 37652
rect 25280 37612 25286 37624
rect 26234 37612 26240 37624
rect 26292 37612 26298 37664
rect 26694 37612 26700 37664
rect 26752 37652 26758 37664
rect 26789 37655 26847 37661
rect 26789 37652 26801 37655
rect 26752 37624 26801 37652
rect 26752 37612 26758 37624
rect 26789 37621 26801 37624
rect 26835 37621 26847 37655
rect 27448 37652 27476 37692
rect 30024 37664 30052 37760
rect 30193 37757 30205 37760
rect 30239 37757 30251 37791
rect 30193 37751 30251 37757
rect 31202 37748 31208 37800
rect 31260 37788 31266 37800
rect 32125 37791 32183 37797
rect 32125 37788 32137 37791
rect 31260 37760 32137 37788
rect 31260 37748 31266 37760
rect 32125 37757 32137 37760
rect 32171 37757 32183 37791
rect 32125 37751 32183 37757
rect 32674 37748 32680 37800
rect 32732 37788 32738 37800
rect 33428 37788 33456 37828
rect 33781 37825 33793 37828
rect 33827 37825 33839 37859
rect 33781 37819 33839 37825
rect 32732 37760 33456 37788
rect 33597 37791 33655 37797
rect 32732 37748 32738 37760
rect 33597 37757 33609 37791
rect 33643 37757 33655 37791
rect 33597 37751 33655 37757
rect 31294 37680 31300 37732
rect 31352 37720 31358 37732
rect 32769 37723 32827 37729
rect 32769 37720 32781 37723
rect 31352 37692 32781 37720
rect 31352 37680 31358 37692
rect 32769 37689 32781 37692
rect 32815 37689 32827 37723
rect 33612 37720 33640 37751
rect 32769 37683 32827 37689
rect 32876 37692 33640 37720
rect 27706 37652 27712 37664
rect 27448 37624 27712 37652
rect 26789 37615 26847 37621
rect 27706 37612 27712 37624
rect 27764 37612 27770 37664
rect 29546 37612 29552 37664
rect 29604 37612 29610 37664
rect 30006 37612 30012 37664
rect 30064 37612 30070 37664
rect 31846 37612 31852 37664
rect 31904 37612 31910 37664
rect 32214 37612 32220 37664
rect 32272 37652 32278 37664
rect 32876 37652 32904 37692
rect 32272 37624 32904 37652
rect 33137 37655 33195 37661
rect 32272 37612 32278 37624
rect 33137 37621 33149 37655
rect 33183 37652 33195 37655
rect 33226 37652 33232 37664
rect 33183 37624 33232 37652
rect 33183 37621 33195 37624
rect 33137 37615 33195 37621
rect 33226 37612 33232 37624
rect 33284 37612 33290 37664
rect 33962 37612 33968 37664
rect 34020 37612 34026 37664
rect 1104 37562 43884 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 43884 37562
rect 1104 37488 43884 37510
rect 5537 37451 5595 37457
rect 5537 37417 5549 37451
rect 5583 37448 5595 37451
rect 5626 37448 5632 37460
rect 5583 37420 5632 37448
rect 5583 37417 5595 37420
rect 5537 37411 5595 37417
rect 5626 37408 5632 37420
rect 5684 37408 5690 37460
rect 7285 37451 7343 37457
rect 7285 37417 7297 37451
rect 7331 37448 7343 37451
rect 8386 37448 8392 37460
rect 7331 37420 8392 37448
rect 7331 37417 7343 37420
rect 7285 37411 7343 37417
rect 8386 37408 8392 37420
rect 8444 37408 8450 37460
rect 8757 37451 8815 37457
rect 8757 37417 8769 37451
rect 8803 37448 8815 37451
rect 9030 37448 9036 37460
rect 8803 37420 9036 37448
rect 8803 37417 8815 37420
rect 8757 37411 8815 37417
rect 9030 37408 9036 37420
rect 9088 37408 9094 37460
rect 11054 37408 11060 37460
rect 11112 37448 11118 37460
rect 11241 37451 11299 37457
rect 11241 37448 11253 37451
rect 11112 37420 11253 37448
rect 11112 37408 11118 37420
rect 11241 37417 11253 37420
rect 11287 37417 11299 37451
rect 11241 37411 11299 37417
rect 6730 37272 6736 37324
rect 6788 37272 6794 37324
rect 8478 37272 8484 37324
rect 8536 37312 8542 37324
rect 9493 37315 9551 37321
rect 9493 37312 9505 37315
rect 8536 37284 9505 37312
rect 8536 37272 8542 37284
rect 9493 37281 9505 37284
rect 9539 37312 9551 37315
rect 9539 37284 9996 37312
rect 9539 37281 9551 37284
rect 9493 37275 9551 37281
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 1627 37216 2774 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 2317 37179 2375 37185
rect 2317 37145 2329 37179
rect 2363 37145 2375 37179
rect 2317 37139 2375 37145
rect 1210 37068 1216 37120
rect 1268 37108 1274 37120
rect 2332 37108 2360 37139
rect 1268 37080 2360 37108
rect 2746 37108 2774 37216
rect 4154 37204 4160 37256
rect 4212 37244 4218 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 4212 37216 7389 37244
rect 4212 37204 4218 37216
rect 7377 37213 7389 37216
rect 7423 37244 7435 37247
rect 7466 37244 7472 37256
rect 7423 37216 7472 37244
rect 7423 37213 7435 37216
rect 7377 37207 7435 37213
rect 7466 37204 7472 37216
rect 7524 37244 7530 37256
rect 8570 37244 8576 37256
rect 7524 37216 8576 37244
rect 7524 37204 7530 37216
rect 8570 37204 8576 37216
rect 8628 37244 8634 37256
rect 9766 37244 9772 37256
rect 8628 37216 9082 37244
rect 8628 37204 8634 37216
rect 4424 37179 4482 37185
rect 4424 37145 4436 37179
rect 4470 37176 4482 37179
rect 4706 37176 4712 37188
rect 4470 37148 4712 37176
rect 4470 37145 4482 37148
rect 4424 37139 4482 37145
rect 4706 37136 4712 37148
rect 4764 37136 4770 37188
rect 5718 37136 5724 37188
rect 5776 37176 5782 37188
rect 5776 37148 6224 37176
rect 5776 37136 5782 37148
rect 3145 37111 3203 37117
rect 3145 37108 3157 37111
rect 2746 37080 3157 37108
rect 1268 37068 1274 37080
rect 3145 37077 3157 37080
rect 3191 37108 3203 37111
rect 5810 37108 5816 37120
rect 3191 37080 5816 37108
rect 3191 37077 3203 37080
rect 3145 37071 3203 37077
rect 5810 37068 5816 37080
rect 5868 37068 5874 37120
rect 6086 37068 6092 37120
rect 6144 37068 6150 37120
rect 6196 37117 6224 37148
rect 6454 37136 6460 37188
rect 6512 37176 6518 37188
rect 6549 37179 6607 37185
rect 6549 37176 6561 37179
rect 6512 37148 6561 37176
rect 6512 37136 6518 37148
rect 6549 37145 6561 37148
rect 6595 37145 6607 37179
rect 6549 37139 6607 37145
rect 7644 37179 7702 37185
rect 7644 37145 7656 37179
rect 7690 37176 7702 37179
rect 8662 37176 8668 37188
rect 7690 37148 8668 37176
rect 7690 37145 7702 37148
rect 7644 37139 7702 37145
rect 8662 37136 8668 37148
rect 8720 37136 8726 37188
rect 9054 37176 9082 37216
rect 9201 37216 9772 37244
rect 9201 37176 9229 37216
rect 9766 37204 9772 37216
rect 9824 37244 9830 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9824 37216 9873 37244
rect 9824 37204 9830 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9968 37244 9996 37284
rect 11256 37244 11284 37411
rect 11330 37408 11336 37460
rect 11388 37448 11394 37460
rect 12894 37448 12900 37460
rect 11388 37420 12900 37448
rect 11388 37408 11394 37420
rect 12894 37408 12900 37420
rect 12952 37408 12958 37460
rect 13817 37451 13875 37457
rect 13817 37417 13829 37451
rect 13863 37448 13875 37451
rect 13998 37448 14004 37460
rect 13863 37420 14004 37448
rect 13863 37417 13875 37420
rect 13817 37411 13875 37417
rect 13998 37408 14004 37420
rect 14056 37448 14062 37460
rect 14056 37420 14228 37448
rect 14056 37408 14062 37420
rect 11422 37340 11428 37392
rect 11480 37380 11486 37392
rect 11480 37352 12434 37380
rect 11480 37340 11486 37352
rect 11977 37315 12035 37321
rect 11977 37281 11989 37315
rect 12023 37312 12035 37315
rect 12158 37312 12164 37324
rect 12023 37284 12164 37312
rect 12023 37281 12035 37284
rect 11977 37275 12035 37281
rect 12158 37272 12164 37284
rect 12216 37272 12222 37324
rect 12406 37312 12434 37352
rect 13262 37340 13268 37392
rect 13320 37340 13326 37392
rect 13906 37380 13912 37392
rect 13556 37352 13912 37380
rect 12805 37315 12863 37321
rect 12805 37312 12817 37315
rect 12406 37284 12817 37312
rect 12805 37281 12817 37284
rect 12851 37312 12863 37315
rect 13280 37312 13308 37340
rect 13556 37321 13584 37352
rect 13906 37340 13912 37352
rect 13964 37340 13970 37392
rect 14200 37380 14228 37420
rect 14274 37408 14280 37460
rect 14332 37408 14338 37460
rect 14458 37408 14464 37460
rect 14516 37408 14522 37460
rect 17034 37448 17040 37460
rect 14660 37420 17040 37448
rect 14660 37380 14688 37420
rect 17034 37408 17040 37420
rect 17092 37408 17098 37460
rect 18046 37408 18052 37460
rect 18104 37448 18110 37460
rect 18104 37420 19334 37448
rect 18104 37408 18110 37420
rect 14200 37352 14688 37380
rect 17494 37340 17500 37392
rect 17552 37340 17558 37392
rect 19061 37383 19119 37389
rect 19061 37349 19073 37383
rect 19107 37349 19119 37383
rect 19306 37380 19334 37420
rect 19794 37408 19800 37460
rect 19852 37448 19858 37460
rect 29546 37448 29552 37460
rect 19852 37420 20392 37448
rect 19852 37408 19858 37420
rect 20364 37389 20392 37420
rect 23124 37420 29552 37448
rect 20349 37383 20407 37389
rect 19306 37352 20024 37380
rect 19061 37343 19119 37349
rect 12851 37284 13308 37312
rect 13541 37315 13599 37321
rect 12851 37281 12863 37284
rect 12805 37275 12863 37281
rect 13541 37281 13553 37315
rect 13587 37281 13599 37315
rect 13541 37275 13599 37281
rect 13630 37272 13636 37324
rect 13688 37272 13694 37324
rect 14182 37272 14188 37324
rect 14240 37272 14246 37324
rect 14642 37272 14648 37324
rect 14700 37272 14706 37324
rect 16482 37272 16488 37324
rect 16540 37312 16546 37324
rect 16853 37315 16911 37321
rect 16540 37284 16804 37312
rect 16540 37272 16546 37284
rect 11701 37247 11759 37253
rect 11701 37244 11713 37247
rect 9968 37216 11100 37244
rect 11256 37216 11713 37244
rect 9861 37207 9919 37213
rect 11072 37188 11100 37216
rect 11701 37213 11713 37216
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 11790 37204 11796 37256
rect 11848 37244 11854 37256
rect 12621 37247 12679 37253
rect 12621 37244 12633 37247
rect 11848 37216 12633 37244
rect 11848 37204 11854 37216
rect 12621 37213 12633 37216
rect 12667 37213 12679 37247
rect 12621 37207 12679 37213
rect 13170 37204 13176 37256
rect 13228 37204 13234 37256
rect 13265 37247 13323 37253
rect 13265 37213 13277 37247
rect 13311 37244 13323 37247
rect 13354 37244 13360 37256
rect 13311 37216 13360 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 13354 37204 13360 37216
rect 13412 37204 13418 37256
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 14200 37244 14228 37272
rect 14918 37253 14924 37256
rect 14912 37244 14924 37253
rect 13771 37216 14228 37244
rect 14879 37216 14924 37244
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 14912 37207 14924 37216
rect 9054 37148 9229 37176
rect 9309 37179 9367 37185
rect 9309 37145 9321 37179
rect 9355 37176 9367 37179
rect 9674 37176 9680 37188
rect 9355 37148 9680 37176
rect 9355 37145 9367 37148
rect 9309 37139 9367 37145
rect 9674 37136 9680 37148
rect 9732 37136 9738 37188
rect 10128 37179 10186 37185
rect 10128 37145 10140 37179
rect 10174 37176 10186 37179
rect 10962 37176 10968 37188
rect 10174 37148 10968 37176
rect 10174 37145 10186 37148
rect 10128 37139 10186 37145
rect 10962 37136 10968 37148
rect 11020 37136 11026 37188
rect 11054 37136 11060 37188
rect 11112 37176 11118 37188
rect 13740 37176 13768 37207
rect 14918 37204 14924 37207
rect 14976 37204 14982 37256
rect 16669 37247 16727 37253
rect 16669 37213 16681 37247
rect 16715 37213 16727 37247
rect 16669 37207 16727 37213
rect 11112 37148 13768 37176
rect 14093 37179 14151 37185
rect 11112 37136 11118 37148
rect 14093 37145 14105 37179
rect 14139 37145 14151 37179
rect 14093 37139 14151 37145
rect 14309 37179 14367 37185
rect 14309 37145 14321 37179
rect 14355 37176 14367 37179
rect 14550 37176 14556 37188
rect 14355 37148 14556 37176
rect 14355 37145 14367 37148
rect 14309 37139 14367 37145
rect 6181 37111 6239 37117
rect 6181 37077 6193 37111
rect 6227 37077 6239 37111
rect 6181 37071 6239 37077
rect 6638 37068 6644 37120
rect 6696 37068 6702 37120
rect 8938 37068 8944 37120
rect 8996 37068 9002 37120
rect 9398 37068 9404 37120
rect 9456 37068 9462 37120
rect 11330 37068 11336 37120
rect 11388 37068 11394 37120
rect 11793 37111 11851 37117
rect 11793 37077 11805 37111
rect 11839 37108 11851 37111
rect 11882 37108 11888 37120
rect 11839 37080 11888 37108
rect 11839 37077 11851 37080
rect 11793 37071 11851 37077
rect 11882 37068 11888 37080
rect 11940 37068 11946 37120
rect 12158 37068 12164 37120
rect 12216 37068 12222 37120
rect 12526 37068 12532 37120
rect 12584 37068 12590 37120
rect 12986 37068 12992 37120
rect 13044 37068 13050 37120
rect 13170 37068 13176 37120
rect 13228 37108 13234 37120
rect 14108 37108 14136 37139
rect 14550 37136 14556 37148
rect 14608 37136 14614 37188
rect 14752 37148 16344 37176
rect 14752 37108 14780 37148
rect 16316 37120 16344 37148
rect 13228 37080 14780 37108
rect 13228 37068 13234 37080
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 16025 37111 16083 37117
rect 16025 37108 16037 37111
rect 14884 37080 16037 37108
rect 14884 37068 14890 37080
rect 16025 37077 16037 37080
rect 16071 37077 16083 37111
rect 16025 37071 16083 37077
rect 16298 37068 16304 37120
rect 16356 37068 16362 37120
rect 16482 37068 16488 37120
rect 16540 37108 16546 37120
rect 16684 37108 16712 37207
rect 16776 37185 16804 37284
rect 16853 37281 16865 37315
rect 16899 37312 16911 37315
rect 19076 37312 19104 37343
rect 19242 37312 19248 37324
rect 16899 37284 17264 37312
rect 19076 37284 19248 37312
rect 16899 37281 16911 37284
rect 16853 37275 16911 37281
rect 17236 37256 17264 37284
rect 19242 37272 19248 37284
rect 19300 37312 19306 37324
rect 19996 37321 20024 37352
rect 20349 37349 20361 37383
rect 20395 37349 20407 37383
rect 23124 37380 23152 37420
rect 29546 37408 29552 37420
rect 29604 37408 29610 37460
rect 33134 37448 33140 37460
rect 31726 37420 33140 37448
rect 24210 37380 24216 37392
rect 20349 37343 20407 37349
rect 21284 37352 23152 37380
rect 23216 37352 24216 37380
rect 19337 37315 19395 37321
rect 19337 37312 19349 37315
rect 19300 37284 19349 37312
rect 19300 37272 19306 37284
rect 19337 37281 19349 37284
rect 19383 37281 19395 37315
rect 19337 37275 19395 37281
rect 19981 37315 20039 37321
rect 19981 37281 19993 37315
rect 20027 37312 20039 37315
rect 20438 37312 20444 37324
rect 20027 37284 20444 37312
rect 20027 37281 20039 37284
rect 19981 37275 20039 37281
rect 20438 37272 20444 37284
rect 20496 37272 20502 37324
rect 21284 37321 21312 37352
rect 21269 37315 21327 37321
rect 21269 37281 21281 37315
rect 21315 37281 21327 37315
rect 21269 37275 21327 37281
rect 21453 37315 21511 37321
rect 21453 37281 21465 37315
rect 21499 37312 21511 37315
rect 21542 37312 21548 37324
rect 21499 37284 21548 37312
rect 21499 37281 21511 37284
rect 21453 37275 21511 37281
rect 21542 37272 21548 37284
rect 21600 37312 21606 37324
rect 21600 37284 21864 37312
rect 21600 37272 21606 37284
rect 17218 37204 17224 37256
rect 17276 37204 17282 37256
rect 17586 37204 17592 37256
rect 17644 37244 17650 37256
rect 17681 37247 17739 37253
rect 17681 37244 17693 37247
rect 17644 37216 17693 37244
rect 17644 37204 17650 37216
rect 17681 37213 17693 37216
rect 17727 37213 17739 37247
rect 17681 37207 17739 37213
rect 17948 37247 18006 37253
rect 17948 37213 17960 37247
rect 17994 37244 18006 37247
rect 18782 37244 18788 37256
rect 17994 37216 18788 37244
rect 17994 37213 18006 37216
rect 17948 37207 18006 37213
rect 18782 37204 18788 37216
rect 18840 37204 18846 37256
rect 19794 37244 19800 37256
rect 18892 37216 19800 37244
rect 16761 37179 16819 37185
rect 16761 37145 16773 37179
rect 16807 37176 16819 37179
rect 16850 37176 16856 37188
rect 16807 37148 16856 37176
rect 16807 37145 16819 37148
rect 16761 37139 16819 37145
rect 16850 37136 16856 37148
rect 16908 37136 16914 37188
rect 17034 37136 17040 37188
rect 17092 37176 17098 37188
rect 17129 37179 17187 37185
rect 17129 37176 17141 37179
rect 17092 37148 17141 37176
rect 17092 37136 17098 37148
rect 17129 37145 17141 37148
rect 17175 37176 17187 37179
rect 17402 37176 17408 37188
rect 17175 37148 17408 37176
rect 17175 37145 17187 37148
rect 17129 37139 17187 37145
rect 17402 37136 17408 37148
rect 17460 37136 17466 37188
rect 17862 37108 17868 37120
rect 16540 37080 17868 37108
rect 16540 37068 16546 37080
rect 17862 37068 17868 37080
rect 17920 37068 17926 37120
rect 17954 37068 17960 37120
rect 18012 37108 18018 37120
rect 18892 37108 18920 37216
rect 19794 37204 19800 37216
rect 19852 37204 19858 37256
rect 20165 37247 20223 37253
rect 20165 37246 20177 37247
rect 20088 37244 20177 37246
rect 19904 37218 20177 37244
rect 19904 37216 20116 37218
rect 19242 37136 19248 37188
rect 19300 37176 19306 37188
rect 19904 37176 19932 37216
rect 20165 37213 20177 37218
rect 20211 37213 20223 37247
rect 21836 37244 21864 37284
rect 22204 37253 22232 37352
rect 22925 37315 22983 37321
rect 22925 37281 22937 37315
rect 22971 37312 22983 37315
rect 23216 37312 23244 37352
rect 24210 37340 24216 37352
rect 24268 37340 24274 37392
rect 25222 37380 25228 37392
rect 24780 37352 25228 37380
rect 24780 37324 24808 37352
rect 25222 37340 25228 37352
rect 25280 37340 25286 37392
rect 26234 37340 26240 37392
rect 26292 37380 26298 37392
rect 27341 37383 27399 37389
rect 27341 37380 27353 37383
rect 26292 37352 27353 37380
rect 26292 37340 26298 37352
rect 27341 37349 27353 37352
rect 27387 37349 27399 37383
rect 27341 37343 27399 37349
rect 28718 37340 28724 37392
rect 28776 37380 28782 37392
rect 31726 37380 31754 37420
rect 33134 37408 33140 37420
rect 33192 37408 33198 37460
rect 33594 37408 33600 37460
rect 33652 37408 33658 37460
rect 28776 37352 31800 37380
rect 28776 37340 28782 37352
rect 22971 37284 23244 37312
rect 22971 37281 22983 37284
rect 22925 37275 22983 37281
rect 23290 37272 23296 37324
rect 23348 37312 23354 37324
rect 23845 37315 23903 37321
rect 23845 37312 23857 37315
rect 23348 37284 23857 37312
rect 23348 37272 23354 37284
rect 23845 37281 23857 37284
rect 23891 37312 23903 37315
rect 24762 37312 24768 37324
rect 23891 37284 24768 37312
rect 23891 37281 23903 37284
rect 23845 37275 23903 37281
rect 24762 37272 24768 37284
rect 24820 37272 24826 37324
rect 24857 37315 24915 37321
rect 24857 37281 24869 37315
rect 24903 37312 24915 37315
rect 27430 37312 27436 37324
rect 24903 37284 25176 37312
rect 24903 37281 24915 37284
rect 24857 37275 24915 37281
rect 20165 37207 20223 37213
rect 21008 37216 21864 37244
rect 19300 37148 19932 37176
rect 19300 37136 19306 37148
rect 21008 37120 21036 37216
rect 18012 37080 18920 37108
rect 18012 37068 18018 37080
rect 19150 37068 19156 37120
rect 19208 37108 19214 37120
rect 19889 37111 19947 37117
rect 19889 37108 19901 37111
rect 19208 37080 19901 37108
rect 19208 37068 19214 37080
rect 19889 37077 19901 37080
rect 19935 37077 19947 37111
rect 19889 37071 19947 37077
rect 20806 37068 20812 37120
rect 20864 37068 20870 37120
rect 20990 37068 20996 37120
rect 21048 37068 21054 37120
rect 21177 37111 21235 37117
rect 21177 37077 21189 37111
rect 21223 37108 21235 37111
rect 21726 37108 21732 37120
rect 21223 37080 21732 37108
rect 21223 37077 21235 37080
rect 21177 37071 21235 37077
rect 21726 37068 21732 37080
rect 21784 37068 21790 37120
rect 21836 37108 21864 37216
rect 22097 37247 22155 37253
rect 22097 37213 22109 37247
rect 22143 37213 22155 37247
rect 22097 37207 22155 37213
rect 22189 37247 22247 37253
rect 22189 37213 22201 37247
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22112 37176 22140 37207
rect 22278 37204 22284 37256
rect 22336 37244 22342 37256
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 22336 37216 22385 37244
rect 22336 37204 22342 37216
rect 22373 37213 22385 37216
rect 22419 37244 22431 37247
rect 23938 37247 23996 37253
rect 22419 37216 23888 37244
rect 22419 37213 22431 37216
rect 22373 37207 22431 37213
rect 23860 37188 23888 37216
rect 23938 37213 23950 37247
rect 23984 37213 23996 37247
rect 23938 37207 23996 37213
rect 22462 37176 22468 37188
rect 22112 37148 22468 37176
rect 22462 37136 22468 37148
rect 22520 37136 22526 37188
rect 22830 37136 22836 37188
rect 22888 37136 22894 37188
rect 23842 37136 23848 37188
rect 23900 37136 23906 37188
rect 23952 37176 23980 37207
rect 24026 37204 24032 37256
rect 24084 37204 24090 37256
rect 24118 37204 24124 37256
rect 24176 37244 24182 37256
rect 24394 37244 24400 37256
rect 24176 37216 24400 37244
rect 24176 37204 24182 37216
rect 24394 37204 24400 37216
rect 24452 37244 24458 37256
rect 24452 37216 24905 37244
rect 24452 37204 24458 37216
rect 24210 37176 24216 37188
rect 23952 37148 24216 37176
rect 24210 37136 24216 37148
rect 24268 37136 24274 37188
rect 24877 37176 24905 37216
rect 24946 37204 24952 37256
rect 25004 37204 25010 37256
rect 25041 37247 25099 37253
rect 25041 37213 25053 37247
rect 25087 37213 25099 37247
rect 25041 37207 25099 37213
rect 25056 37176 25084 37207
rect 24320 37148 24716 37176
rect 24877 37148 25084 37176
rect 22278 37108 22284 37120
rect 21836 37080 22284 37108
rect 22278 37068 22284 37080
rect 22336 37068 22342 37120
rect 22554 37068 22560 37120
rect 22612 37108 22618 37120
rect 23106 37108 23112 37120
rect 22612 37080 23112 37108
rect 22612 37068 22618 37080
rect 23106 37068 23112 37080
rect 23164 37068 23170 37120
rect 23566 37068 23572 37120
rect 23624 37068 23630 37120
rect 23661 37111 23719 37117
rect 23661 37077 23673 37111
rect 23707 37108 23719 37111
rect 24320 37108 24348 37148
rect 23707 37080 24348 37108
rect 23707 37077 23719 37080
rect 23661 37071 23719 37077
rect 24578 37068 24584 37120
rect 24636 37068 24642 37120
rect 24688 37108 24716 37148
rect 25038 37108 25044 37120
rect 24688 37080 25044 37108
rect 25038 37068 25044 37080
rect 25096 37068 25102 37120
rect 25148 37108 25176 37284
rect 26620 37284 27436 37312
rect 25225 37247 25283 37253
rect 25225 37213 25237 37247
rect 25271 37244 25283 37247
rect 26620 37244 26648 37284
rect 27430 37272 27436 37284
rect 27488 37272 27494 37324
rect 29270 37272 29276 37324
rect 29328 37312 29334 37324
rect 29546 37312 29552 37324
rect 29328 37284 29552 37312
rect 29328 37272 29334 37284
rect 29546 37272 29552 37284
rect 29604 37272 29610 37324
rect 31202 37312 31208 37324
rect 29932 37284 31208 37312
rect 25271 37216 26648 37244
rect 25271 37213 25283 37216
rect 25225 37207 25283 37213
rect 26694 37204 26700 37256
rect 26752 37204 26758 37256
rect 26786 37204 26792 37256
rect 26844 37204 26850 37256
rect 26970 37204 26976 37256
rect 27028 37244 27034 37256
rect 27709 37247 27767 37253
rect 27709 37244 27721 37247
rect 27028 37216 27721 37244
rect 27028 37204 27034 37216
rect 27709 37213 27721 37216
rect 27755 37213 27767 37247
rect 27709 37207 27767 37213
rect 27976 37247 28034 37253
rect 27976 37213 27988 37247
rect 28022 37244 28034 37247
rect 29638 37244 29644 37256
rect 28022 37216 29644 37244
rect 28022 37213 28034 37216
rect 27976 37207 28034 37213
rect 29638 37204 29644 37216
rect 29696 37204 29702 37256
rect 29730 37204 29736 37256
rect 29788 37204 29794 37256
rect 25492 37179 25550 37185
rect 25492 37145 25504 37179
rect 25538 37176 25550 37179
rect 26712 37176 26740 37204
rect 29932 37176 29960 37284
rect 31202 37272 31208 37284
rect 31260 37272 31266 37324
rect 31772 37321 31800 37352
rect 31757 37315 31815 37321
rect 31757 37281 31769 37315
rect 31803 37281 31815 37315
rect 31757 37275 31815 37281
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31021 37247 31079 37253
rect 31021 37244 31033 37247
rect 30984 37216 31033 37244
rect 30984 37204 30990 37216
rect 31021 37213 31033 37216
rect 31067 37213 31079 37247
rect 31021 37207 31079 37213
rect 31110 37204 31116 37256
rect 31168 37204 31174 37256
rect 31297 37247 31355 37253
rect 31297 37213 31309 37247
rect 31343 37244 31355 37247
rect 31386 37244 31392 37256
rect 31343 37216 31392 37244
rect 31343 37213 31355 37216
rect 31297 37207 31355 37213
rect 31386 37204 31392 37216
rect 31444 37204 31450 37256
rect 31941 37247 31999 37253
rect 31941 37213 31953 37247
rect 31987 37213 31999 37247
rect 31941 37207 31999 37213
rect 32208 37247 32266 37253
rect 32208 37213 32220 37247
rect 32254 37244 32266 37247
rect 33962 37244 33968 37256
rect 32254 37216 33968 37244
rect 32254 37213 32266 37216
rect 32208 37207 32266 37213
rect 25538 37148 26740 37176
rect 29104 37148 29960 37176
rect 25538 37145 25550 37148
rect 25492 37139 25550 37145
rect 26510 37108 26516 37120
rect 25148 37080 26516 37108
rect 26510 37068 26516 37080
rect 26568 37068 26574 37120
rect 26602 37068 26608 37120
rect 26660 37068 26666 37120
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27614 37108 27620 37120
rect 27120 37080 27620 37108
rect 27120 37068 27126 37080
rect 27614 37068 27620 37080
rect 27672 37068 27678 37120
rect 29104 37117 29132 37148
rect 30006 37136 30012 37188
rect 30064 37176 30070 37188
rect 31956 37176 31984 37207
rect 33962 37204 33968 37216
rect 34020 37204 34026 37256
rect 30064 37148 31984 37176
rect 30064 37136 30070 37148
rect 29089 37111 29147 37117
rect 29089 37077 29101 37111
rect 29135 37077 29147 37111
rect 29089 37071 29147 37077
rect 29270 37068 29276 37120
rect 29328 37108 29334 37120
rect 30285 37111 30343 37117
rect 30285 37108 30297 37111
rect 29328 37080 30297 37108
rect 29328 37068 29334 37080
rect 30285 37077 30297 37080
rect 30331 37077 30343 37111
rect 30285 37071 30343 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30561 37111 30619 37117
rect 30561 37108 30573 37111
rect 30432 37080 30573 37108
rect 30432 37068 30438 37080
rect 30561 37077 30573 37080
rect 30607 37077 30619 37111
rect 30561 37071 30619 37077
rect 31110 37068 31116 37120
rect 31168 37108 31174 37120
rect 32030 37108 32036 37120
rect 31168 37080 32036 37108
rect 31168 37068 31174 37080
rect 32030 37068 32036 37080
rect 32088 37068 32094 37120
rect 33318 37068 33324 37120
rect 33376 37068 33382 37120
rect 1104 37018 43884 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 43884 37018
rect 1104 36944 43884 36966
rect 5537 36907 5595 36913
rect 5537 36904 5549 36907
rect 3528 36876 5549 36904
rect 3528 36777 3556 36876
rect 5537 36873 5549 36876
rect 5583 36873 5595 36907
rect 5537 36867 5595 36873
rect 6365 36907 6423 36913
rect 6365 36873 6377 36907
rect 6411 36904 6423 36907
rect 6638 36904 6644 36916
rect 6411 36876 6644 36904
rect 6411 36873 6423 36876
rect 6365 36867 6423 36873
rect 4424 36839 4482 36845
rect 4424 36805 4436 36839
rect 4470 36836 4482 36839
rect 5442 36836 5448 36848
rect 4470 36808 5448 36836
rect 4470 36805 4482 36808
rect 4424 36799 4482 36805
rect 5442 36796 5448 36808
rect 5500 36796 5506 36848
rect 5552 36836 5580 36867
rect 6638 36864 6644 36876
rect 6696 36864 6702 36916
rect 7929 36907 7987 36913
rect 7929 36873 7941 36907
rect 7975 36904 7987 36907
rect 8297 36907 8355 36913
rect 8297 36904 8309 36907
rect 7975 36876 8309 36904
rect 7975 36873 7987 36876
rect 7929 36867 7987 36873
rect 8297 36873 8309 36876
rect 8343 36873 8355 36907
rect 8297 36867 8355 36873
rect 8757 36907 8815 36913
rect 8757 36873 8769 36907
rect 8803 36904 8815 36907
rect 9674 36904 9680 36916
rect 8803 36876 9680 36904
rect 8803 36873 8815 36876
rect 8757 36867 8815 36873
rect 9674 36864 9680 36876
rect 9732 36864 9738 36916
rect 11330 36864 11336 36916
rect 11388 36904 11394 36916
rect 11977 36907 12035 36913
rect 11977 36904 11989 36907
rect 11388 36876 11989 36904
rect 11388 36864 11394 36876
rect 11977 36873 11989 36876
rect 12023 36873 12035 36907
rect 12986 36904 12992 36916
rect 11977 36867 12035 36873
rect 12406 36876 12992 36904
rect 6825 36839 6883 36845
rect 6825 36836 6837 36839
rect 5552 36808 6837 36836
rect 6825 36805 6837 36808
rect 6871 36805 6883 36839
rect 6825 36799 6883 36805
rect 7208 36808 11468 36836
rect 3513 36771 3571 36777
rect 3513 36737 3525 36771
rect 3559 36737 3571 36771
rect 3513 36731 3571 36737
rect 4154 36728 4160 36780
rect 4212 36728 4218 36780
rect 5626 36728 5632 36780
rect 5684 36768 5690 36780
rect 6733 36771 6791 36777
rect 6733 36768 6745 36771
rect 5684 36740 6745 36768
rect 5684 36728 5690 36740
rect 6733 36737 6745 36740
rect 6779 36737 6791 36771
rect 7006 36768 7012 36780
rect 6733 36731 6791 36737
rect 6932 36740 7012 36768
rect 6638 36660 6644 36712
rect 6696 36660 6702 36712
rect 6932 36709 6960 36740
rect 7006 36728 7012 36740
rect 7064 36728 7070 36780
rect 7208 36777 7236 36808
rect 7193 36771 7251 36777
rect 7193 36737 7205 36771
rect 7239 36737 7251 36771
rect 7193 36731 7251 36737
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 8202 36768 8208 36780
rect 7883 36740 8208 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 8202 36728 8208 36740
rect 8260 36728 8266 36780
rect 8665 36771 8723 36777
rect 8665 36737 8677 36771
rect 8711 36768 8723 36771
rect 9582 36768 9588 36780
rect 8711 36740 9588 36768
rect 8711 36737 8723 36740
rect 8665 36731 8723 36737
rect 9582 36728 9588 36740
rect 9640 36728 9646 36780
rect 9766 36728 9772 36780
rect 9824 36728 9830 36780
rect 10036 36771 10094 36777
rect 10036 36737 10048 36771
rect 10082 36768 10094 36771
rect 11054 36768 11060 36780
rect 10082 36740 11060 36768
rect 10082 36737 10094 36740
rect 10036 36731 10094 36737
rect 11054 36728 11060 36740
rect 11112 36728 11118 36780
rect 11440 36768 11468 36808
rect 11514 36796 11520 36848
rect 11572 36836 11578 36848
rect 11885 36839 11943 36845
rect 11885 36836 11897 36839
rect 11572 36808 11897 36836
rect 11572 36796 11578 36808
rect 11885 36805 11897 36808
rect 11931 36805 11943 36839
rect 11885 36799 11943 36805
rect 12406 36768 12434 36876
rect 12986 36864 12992 36876
rect 13044 36864 13050 36916
rect 13538 36864 13544 36916
rect 13596 36904 13602 36916
rect 14550 36904 14556 36916
rect 13596 36876 14556 36904
rect 13596 36864 13602 36876
rect 14550 36864 14556 36876
rect 14608 36904 14614 36916
rect 17586 36904 17592 36916
rect 14608 36876 17592 36904
rect 14608 36864 14614 36876
rect 13906 36796 13912 36848
rect 13964 36796 13970 36848
rect 14921 36839 14979 36845
rect 14921 36836 14933 36839
rect 14108 36808 14933 36836
rect 11440 36740 12434 36768
rect 12529 36771 12587 36777
rect 12529 36737 12541 36771
rect 12575 36768 12587 36771
rect 13354 36768 13360 36780
rect 12575 36740 13360 36768
rect 12575 36737 12587 36740
rect 12529 36731 12587 36737
rect 13354 36728 13360 36740
rect 13412 36728 13418 36780
rect 6917 36703 6975 36709
rect 6917 36669 6929 36703
rect 6963 36669 6975 36703
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 6917 36663 6975 36669
rect 7024 36672 8033 36700
rect 6656 36632 6684 36660
rect 7024 36632 7052 36672
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 6656 36604 7052 36632
rect 7098 36592 7104 36644
rect 7156 36632 7162 36644
rect 8036 36632 8064 36663
rect 8110 36660 8116 36712
rect 8168 36700 8174 36712
rect 8941 36703 8999 36709
rect 8941 36700 8953 36703
rect 8168 36672 8953 36700
rect 8168 36660 8174 36672
rect 8941 36669 8953 36672
rect 8987 36700 8999 36703
rect 9490 36700 9496 36712
rect 8987 36672 9496 36700
rect 8987 36669 8999 36672
rect 8941 36663 8999 36669
rect 9490 36660 9496 36672
rect 9548 36660 9554 36712
rect 12066 36700 12072 36712
rect 10796 36672 12072 36700
rect 7156 36604 7512 36632
rect 8036 36604 9812 36632
rect 7156 36592 7162 36604
rect 4062 36524 4068 36576
rect 4120 36524 4126 36576
rect 6086 36524 6092 36576
rect 6144 36524 6150 36576
rect 6730 36524 6736 36576
rect 6788 36564 6794 36576
rect 7484 36573 7512 36604
rect 7285 36567 7343 36573
rect 7285 36564 7297 36567
rect 6788 36536 7297 36564
rect 6788 36524 6794 36536
rect 7285 36533 7297 36536
rect 7331 36533 7343 36567
rect 7285 36527 7343 36533
rect 7469 36567 7527 36573
rect 7469 36533 7481 36567
rect 7515 36533 7527 36567
rect 7469 36527 7527 36533
rect 8754 36524 8760 36576
rect 8812 36564 8818 36576
rect 9030 36564 9036 36576
rect 8812 36536 9036 36564
rect 8812 36524 8818 36536
rect 9030 36524 9036 36536
rect 9088 36564 9094 36576
rect 9585 36567 9643 36573
rect 9585 36564 9597 36567
rect 9088 36536 9597 36564
rect 9088 36524 9094 36536
rect 9585 36533 9597 36536
rect 9631 36533 9643 36567
rect 9784 36564 9812 36604
rect 10796 36564 10824 36672
rect 12066 36660 12072 36672
rect 12124 36660 12130 36712
rect 12618 36660 12624 36712
rect 12676 36700 12682 36712
rect 13265 36703 13323 36709
rect 13265 36700 13277 36703
rect 12676 36672 13277 36700
rect 12676 36660 12682 36672
rect 13265 36669 13277 36672
rect 13311 36669 13323 36703
rect 13924 36700 13952 36796
rect 14108 36780 14136 36808
rect 14921 36805 14933 36808
rect 14967 36805 14979 36839
rect 14921 36799 14979 36805
rect 14090 36728 14096 36780
rect 14148 36728 14154 36780
rect 15212 36777 15240 36876
rect 17586 36864 17592 36876
rect 17644 36904 17650 36916
rect 17954 36904 17960 36916
rect 17644 36876 17960 36904
rect 17644 36864 17650 36876
rect 17954 36864 17960 36876
rect 18012 36864 18018 36916
rect 18141 36907 18199 36913
rect 18141 36873 18153 36907
rect 18187 36904 18199 36907
rect 18414 36904 18420 36916
rect 18187 36876 18420 36904
rect 18187 36873 18199 36876
rect 18141 36867 18199 36873
rect 18414 36864 18420 36876
rect 18472 36864 18478 36916
rect 18509 36907 18567 36913
rect 18509 36873 18521 36907
rect 18555 36904 18567 36907
rect 19150 36904 19156 36916
rect 18555 36876 19156 36904
rect 18555 36873 18567 36876
rect 18509 36867 18567 36873
rect 19150 36864 19156 36876
rect 19208 36864 19214 36916
rect 20806 36904 20812 36916
rect 20088 36876 20812 36904
rect 15488 36808 16528 36836
rect 15488 36777 15516 36808
rect 16500 36780 16528 36808
rect 16850 36796 16856 36848
rect 16908 36836 16914 36848
rect 17221 36839 17279 36845
rect 17221 36836 17233 36839
rect 16908 36808 17233 36836
rect 16908 36796 16914 36808
rect 17221 36805 17233 36808
rect 17267 36836 17279 36839
rect 17267 36808 19012 36836
rect 17267 36805 17279 36808
rect 17221 36799 17279 36805
rect 14737 36771 14795 36777
rect 14737 36737 14749 36771
rect 14783 36766 14795 36771
rect 15013 36771 15071 36777
rect 15013 36768 15025 36771
rect 14783 36738 14872 36766
rect 14783 36737 14795 36738
rect 14737 36731 14795 36737
rect 13924 36672 14228 36700
rect 13265 36663 13323 36669
rect 11149 36635 11207 36641
rect 11149 36601 11161 36635
rect 11195 36632 11207 36635
rect 11195 36604 11928 36632
rect 11195 36601 11207 36604
rect 11149 36595 11207 36601
rect 11900 36576 11928 36604
rect 13630 36592 13636 36644
rect 13688 36632 13694 36644
rect 14200 36632 14228 36672
rect 14550 36660 14556 36712
rect 14608 36700 14614 36712
rect 14844 36700 14872 36738
rect 14936 36740 15025 36768
rect 14936 36712 14964 36740
rect 15013 36737 15025 36740
rect 15059 36737 15071 36771
rect 15013 36731 15071 36737
rect 15197 36771 15255 36777
rect 15197 36737 15209 36771
rect 15243 36737 15255 36771
rect 15197 36731 15255 36737
rect 15473 36771 15531 36777
rect 15473 36737 15485 36771
rect 15519 36737 15531 36771
rect 15473 36731 15531 36737
rect 15565 36771 15623 36777
rect 15565 36737 15577 36771
rect 15611 36768 15623 36771
rect 15746 36768 15752 36780
rect 15611 36740 15752 36768
rect 15611 36737 15623 36740
rect 15565 36731 15623 36737
rect 14608 36672 14872 36700
rect 14608 36660 14614 36672
rect 14737 36635 14795 36641
rect 14737 36632 14749 36635
rect 13688 36604 14044 36632
rect 14200 36604 14749 36632
rect 13688 36592 13694 36604
rect 9784 36536 10824 36564
rect 9585 36527 9643 36533
rect 11514 36524 11520 36576
rect 11572 36524 11578 36576
rect 11882 36524 11888 36576
rect 11940 36524 11946 36576
rect 13170 36524 13176 36576
rect 13228 36524 13234 36576
rect 13906 36524 13912 36576
rect 13964 36524 13970 36576
rect 14016 36564 14044 36604
rect 14737 36601 14749 36604
rect 14783 36601 14795 36635
rect 14844 36632 14872 36672
rect 14918 36660 14924 36712
rect 14976 36660 14982 36712
rect 15488 36632 15516 36731
rect 15580 36700 15608 36731
rect 15746 36728 15752 36740
rect 15804 36728 15810 36780
rect 15838 36728 15844 36780
rect 15896 36768 15902 36780
rect 15933 36771 15991 36777
rect 15933 36768 15945 36771
rect 15896 36740 15945 36768
rect 15896 36728 15902 36740
rect 15933 36737 15945 36740
rect 15979 36737 15991 36771
rect 15933 36731 15991 36737
rect 16482 36728 16488 36780
rect 16540 36728 16546 36780
rect 17129 36771 17187 36777
rect 17129 36737 17141 36771
rect 17175 36768 17187 36771
rect 17175 36740 17356 36768
rect 17175 36737 17187 36740
rect 17129 36731 17187 36737
rect 14844 36604 15516 36632
rect 15544 36672 15608 36700
rect 14737 36595 14795 36601
rect 14645 36567 14703 36573
rect 14645 36564 14657 36567
rect 14016 36536 14657 36564
rect 14645 36533 14657 36536
rect 14691 36533 14703 36567
rect 14645 36527 14703 36533
rect 14918 36524 14924 36576
rect 14976 36564 14982 36576
rect 15544 36564 15572 36672
rect 16298 36660 16304 36712
rect 16356 36700 16362 36712
rect 17144 36700 17172 36731
rect 16356 36672 17172 36700
rect 16356 36660 16362 36672
rect 17218 36660 17224 36712
rect 17276 36660 17282 36712
rect 17328 36700 17356 36740
rect 17402 36728 17408 36780
rect 17460 36768 17466 36780
rect 18984 36777 19012 36808
rect 20088 36777 20116 36876
rect 20806 36864 20812 36876
rect 20864 36864 20870 36916
rect 22186 36864 22192 36916
rect 22244 36904 22250 36916
rect 22830 36904 22836 36916
rect 22244 36876 22836 36904
rect 22244 36864 22250 36876
rect 22830 36864 22836 36876
rect 22888 36864 22894 36916
rect 24578 36864 24584 36916
rect 24636 36904 24642 36916
rect 28721 36907 28779 36913
rect 24636 36876 27936 36904
rect 24636 36864 24642 36876
rect 20717 36839 20775 36845
rect 20717 36805 20729 36839
rect 20763 36836 20775 36839
rect 21634 36836 21640 36848
rect 20763 36808 21640 36836
rect 20763 36805 20775 36808
rect 20717 36799 20775 36805
rect 21634 36796 21640 36808
rect 21692 36796 21698 36848
rect 22204 36777 22232 36864
rect 24765 36839 24823 36845
rect 24765 36836 24777 36839
rect 22296 36808 24777 36836
rect 22296 36777 22324 36808
rect 24765 36805 24777 36808
rect 24811 36836 24823 36839
rect 24854 36836 24860 36848
rect 24811 36808 24860 36836
rect 24811 36805 24823 36808
rect 24765 36799 24823 36805
rect 24854 36796 24860 36808
rect 24912 36796 24918 36848
rect 26970 36836 26976 36848
rect 24964 36808 26976 36836
rect 17589 36771 17647 36777
rect 17589 36768 17601 36771
rect 17460 36740 17601 36768
rect 17460 36728 17466 36740
rect 17589 36737 17601 36740
rect 17635 36737 17647 36771
rect 17589 36731 17647 36737
rect 18969 36771 19027 36777
rect 18969 36737 18981 36771
rect 19015 36737 19027 36771
rect 18969 36731 19027 36737
rect 19153 36771 19211 36777
rect 19153 36737 19165 36771
rect 19199 36737 19211 36771
rect 19153 36731 19211 36737
rect 20073 36771 20131 36777
rect 20073 36737 20085 36771
rect 20119 36737 20131 36771
rect 20073 36731 20131 36737
rect 22189 36771 22247 36777
rect 22189 36737 22201 36771
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 22281 36771 22339 36777
rect 22281 36737 22293 36771
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 22465 36771 22523 36777
rect 22465 36737 22477 36771
rect 22511 36768 22523 36771
rect 22511 36740 23060 36768
rect 22511 36737 22523 36740
rect 22465 36731 22523 36737
rect 17328 36672 18000 36700
rect 17972 36644 18000 36672
rect 18598 36660 18604 36712
rect 18656 36660 18662 36712
rect 18690 36660 18696 36712
rect 18748 36660 18754 36712
rect 15654 36592 15660 36644
rect 15712 36632 15718 36644
rect 16393 36635 16451 36641
rect 16393 36632 16405 36635
rect 15712 36604 16405 36632
rect 15712 36592 15718 36604
rect 16393 36601 16405 36604
rect 16439 36601 16451 36635
rect 16393 36595 16451 36601
rect 14976 36536 15572 36564
rect 16408 36564 16436 36595
rect 17126 36592 17132 36644
rect 17184 36632 17190 36644
rect 17773 36635 17831 36641
rect 17773 36632 17785 36635
rect 17184 36604 17785 36632
rect 17184 36592 17190 36604
rect 17773 36601 17785 36604
rect 17819 36601 17831 36635
rect 17773 36595 17831 36601
rect 17954 36592 17960 36644
rect 18012 36592 18018 36644
rect 18708 36632 18736 36660
rect 19168 36644 19196 36731
rect 19242 36660 19248 36712
rect 19300 36660 19306 36712
rect 21450 36660 21456 36712
rect 21508 36660 21514 36712
rect 22925 36703 22983 36709
rect 22925 36669 22937 36703
rect 22971 36669 22983 36703
rect 22925 36663 22983 36669
rect 18064 36604 18736 36632
rect 18064 36564 18092 36604
rect 19150 36592 19156 36644
rect 19208 36632 19214 36644
rect 19208 36604 20392 36632
rect 19208 36592 19214 36604
rect 20364 36576 20392 36604
rect 16408 36536 18092 36564
rect 14976 36524 14982 36536
rect 18506 36524 18512 36576
rect 18564 36564 18570 36576
rect 19061 36567 19119 36573
rect 19061 36564 19073 36567
rect 18564 36536 19073 36564
rect 18564 36524 18570 36536
rect 19061 36533 19073 36536
rect 19107 36533 19119 36567
rect 19061 36527 19119 36533
rect 19334 36524 19340 36576
rect 19392 36564 19398 36576
rect 19889 36567 19947 36573
rect 19889 36564 19901 36567
rect 19392 36536 19901 36564
rect 19392 36524 19398 36536
rect 19889 36533 19901 36536
rect 19935 36533 19947 36567
rect 19889 36527 19947 36533
rect 20346 36524 20352 36576
rect 20404 36524 20410 36576
rect 20622 36524 20628 36576
rect 20680 36524 20686 36576
rect 22940 36564 22968 36663
rect 23032 36632 23060 36740
rect 23106 36728 23112 36780
rect 23164 36728 23170 36780
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 24964 36777 24992 36808
rect 26970 36796 26976 36808
rect 27028 36796 27034 36848
rect 27356 36808 27568 36836
rect 24121 36771 24179 36777
rect 24121 36768 24133 36771
rect 23256 36740 24133 36768
rect 23256 36728 23262 36740
rect 24121 36737 24133 36740
rect 24167 36737 24179 36771
rect 24121 36731 24179 36737
rect 24949 36771 25007 36777
rect 24949 36737 24961 36771
rect 24995 36737 25007 36771
rect 24949 36731 25007 36737
rect 25216 36771 25274 36777
rect 25216 36737 25228 36771
rect 25262 36768 25274 36771
rect 26234 36768 26240 36780
rect 25262 36740 26240 36768
rect 25262 36737 25274 36740
rect 25216 36731 25274 36737
rect 26234 36728 26240 36740
rect 26292 36728 26298 36780
rect 26418 36728 26424 36780
rect 26476 36728 26482 36780
rect 26605 36771 26663 36777
rect 26605 36737 26617 36771
rect 26651 36737 26663 36771
rect 26605 36731 26663 36737
rect 26618 36730 26648 36731
rect 23937 36703 23995 36709
rect 23937 36669 23949 36703
rect 23983 36700 23995 36703
rect 24394 36700 24400 36712
rect 23983 36672 24400 36700
rect 23983 36669 23995 36672
rect 23937 36663 23995 36669
rect 24394 36660 24400 36672
rect 24452 36660 24458 36712
rect 23032 36604 24348 36632
rect 24320 36576 24348 36604
rect 26326 36592 26332 36644
rect 26384 36632 26390 36644
rect 26618 36632 26646 36730
rect 26786 36728 26792 36780
rect 26844 36728 26850 36780
rect 27154 36728 27160 36780
rect 27212 36768 27218 36780
rect 27356 36777 27384 36808
rect 27249 36771 27307 36777
rect 27249 36768 27261 36771
rect 27212 36740 27261 36768
rect 27212 36728 27218 36740
rect 27249 36737 27261 36740
rect 27295 36737 27307 36771
rect 27249 36731 27307 36737
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 27433 36771 27491 36777
rect 27433 36737 27445 36771
rect 27479 36737 27491 36771
rect 27433 36731 27491 36737
rect 26804 36700 26832 36728
rect 26973 36703 27031 36709
rect 26973 36700 26985 36703
rect 26804 36672 26985 36700
rect 26973 36669 26985 36672
rect 27019 36669 27031 36703
rect 26973 36663 27031 36669
rect 26384 36604 26646 36632
rect 26789 36635 26847 36641
rect 26384 36592 26390 36604
rect 26789 36601 26801 36635
rect 26835 36632 26847 36635
rect 27448 36632 27476 36731
rect 26835 36604 27476 36632
rect 27540 36632 27568 36808
rect 27614 36728 27620 36780
rect 27672 36768 27678 36780
rect 27908 36777 27936 36876
rect 28721 36873 28733 36907
rect 28767 36904 28779 36907
rect 28767 36876 29684 36904
rect 28767 36873 28779 36876
rect 28721 36867 28779 36873
rect 28000 36808 28764 36836
rect 27893 36771 27951 36777
rect 27672 36740 27844 36768
rect 27672 36728 27678 36740
rect 27706 36660 27712 36712
rect 27764 36660 27770 36712
rect 27816 36700 27844 36740
rect 27893 36737 27905 36771
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 28000 36700 28028 36808
rect 28074 36728 28080 36780
rect 28132 36728 28138 36780
rect 28169 36771 28227 36777
rect 28169 36737 28181 36771
rect 28215 36768 28227 36771
rect 28350 36768 28356 36780
rect 28215 36740 28356 36768
rect 28215 36737 28227 36740
rect 28169 36731 28227 36737
rect 27816 36672 28028 36700
rect 28184 36632 28212 36731
rect 28350 36728 28356 36740
rect 28408 36728 28414 36780
rect 28626 36728 28632 36780
rect 28684 36728 28690 36780
rect 28736 36768 28764 36808
rect 29178 36796 29184 36848
rect 29236 36836 29242 36848
rect 29656 36836 29684 36876
rect 29730 36864 29736 36916
rect 29788 36904 29794 36916
rect 30190 36904 30196 36916
rect 29788 36876 30196 36904
rect 29788 36864 29794 36876
rect 30190 36864 30196 36876
rect 30248 36904 30254 36916
rect 31389 36907 31447 36913
rect 31389 36904 31401 36907
rect 30248 36876 31401 36904
rect 30248 36864 30254 36876
rect 31389 36873 31401 36876
rect 31435 36873 31447 36907
rect 31389 36867 31447 36873
rect 33134 36864 33140 36916
rect 33192 36864 33198 36916
rect 33226 36864 33232 36916
rect 33284 36904 33290 36916
rect 33413 36907 33471 36913
rect 33413 36904 33425 36907
rect 33284 36876 33425 36904
rect 33284 36864 33290 36876
rect 33413 36873 33425 36876
rect 33459 36873 33471 36907
rect 33413 36867 33471 36873
rect 31294 36836 31300 36848
rect 29236 36808 29592 36836
rect 29656 36808 31300 36836
rect 29236 36796 29242 36808
rect 28736 36740 28948 36768
rect 28534 36660 28540 36712
rect 28592 36700 28598 36712
rect 28813 36703 28871 36709
rect 28813 36700 28825 36703
rect 28592 36672 28825 36700
rect 28592 36660 28598 36672
rect 28813 36669 28825 36672
rect 28859 36669 28871 36703
rect 28920 36700 28948 36740
rect 28994 36728 29000 36780
rect 29052 36768 29058 36780
rect 29362 36768 29368 36780
rect 29052 36740 29368 36768
rect 29052 36728 29058 36740
rect 29362 36728 29368 36740
rect 29420 36728 29426 36780
rect 29454 36728 29460 36780
rect 29512 36728 29518 36780
rect 29564 36777 29592 36808
rect 31294 36796 31300 36808
rect 31352 36796 31358 36848
rect 29549 36771 29607 36777
rect 29549 36737 29561 36771
rect 29595 36737 29607 36771
rect 29549 36731 29607 36737
rect 29733 36771 29791 36777
rect 29733 36737 29745 36771
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 29748 36700 29776 36731
rect 30006 36728 30012 36780
rect 30064 36728 30070 36780
rect 30276 36771 30334 36777
rect 30276 36737 30288 36771
rect 30322 36768 30334 36771
rect 32769 36771 32827 36777
rect 32769 36768 32781 36771
rect 30322 36740 32781 36768
rect 30322 36737 30334 36740
rect 30276 36731 30334 36737
rect 32769 36737 32781 36740
rect 32815 36737 32827 36771
rect 32769 36731 32827 36737
rect 28920 36672 29776 36700
rect 28813 36663 28871 36669
rect 27540 36604 28212 36632
rect 26835 36601 26847 36604
rect 26789 36595 26847 36601
rect 23658 36564 23664 36576
rect 22940 36536 23664 36564
rect 23658 36524 23664 36536
rect 23716 36524 23722 36576
rect 24302 36524 24308 36576
rect 24360 36524 24366 36576
rect 25866 36524 25872 36576
rect 25924 36564 25930 36576
rect 27540 36564 27568 36604
rect 28902 36592 28908 36644
rect 28960 36632 28966 36644
rect 28960 36604 29500 36632
rect 28960 36592 28966 36604
rect 25924 36536 27568 36564
rect 28261 36567 28319 36573
rect 25924 36524 25930 36536
rect 28261 36533 28273 36567
rect 28307 36564 28319 36567
rect 28994 36564 29000 36576
rect 28307 36536 29000 36564
rect 28307 36533 28319 36536
rect 28261 36527 28319 36533
rect 28994 36524 29000 36536
rect 29052 36524 29058 36576
rect 29086 36524 29092 36576
rect 29144 36524 29150 36576
rect 29472 36564 29500 36604
rect 29730 36592 29736 36644
rect 29788 36632 29794 36644
rect 30024 36632 30052 36728
rect 31754 36660 31760 36712
rect 31812 36700 31818 36712
rect 32125 36703 32183 36709
rect 32125 36700 32137 36703
rect 31812 36672 32137 36700
rect 31812 36660 31818 36672
rect 32125 36669 32137 36672
rect 32171 36669 32183 36703
rect 32125 36663 32183 36669
rect 29788 36604 30052 36632
rect 29788 36592 29794 36604
rect 30374 36564 30380 36576
rect 29472 36536 30380 36564
rect 30374 36524 30380 36536
rect 30432 36564 30438 36576
rect 31757 36567 31815 36573
rect 31757 36564 31769 36567
rect 30432 36536 31769 36564
rect 30432 36524 30438 36536
rect 31757 36533 31769 36536
rect 31803 36533 31815 36567
rect 31757 36527 31815 36533
rect 1104 36474 43884 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 43884 36474
rect 1104 36400 43884 36422
rect 4062 36320 4068 36372
rect 4120 36320 4126 36372
rect 4890 36320 4896 36372
rect 4948 36360 4954 36372
rect 5077 36363 5135 36369
rect 5077 36360 5089 36363
rect 4948 36332 5089 36360
rect 4948 36320 4954 36332
rect 5077 36329 5089 36332
rect 5123 36329 5135 36363
rect 5077 36323 5135 36329
rect 5626 36320 5632 36372
rect 5684 36360 5690 36372
rect 8478 36360 8484 36372
rect 5684 36332 8484 36360
rect 5684 36320 5690 36332
rect 8478 36320 8484 36332
rect 8536 36320 8542 36372
rect 10962 36320 10968 36372
rect 11020 36320 11026 36372
rect 11054 36320 11060 36372
rect 11112 36360 11118 36372
rect 11793 36363 11851 36369
rect 11793 36360 11805 36363
rect 11112 36332 11805 36360
rect 11112 36320 11118 36332
rect 11793 36329 11805 36332
rect 11839 36329 11851 36363
rect 12158 36360 12164 36372
rect 11793 36323 11851 36329
rect 11900 36332 12164 36360
rect 4080 36292 4108 36320
rect 8941 36295 8999 36301
rect 8941 36292 8953 36295
rect 4080 36264 5488 36292
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1581 36159 1639 36165
rect 1581 36156 1593 36159
rect 992 36128 1593 36156
rect 992 36116 998 36128
rect 1581 36125 1593 36128
rect 1627 36125 1639 36159
rect 1581 36119 1639 36125
rect 4430 36116 4436 36168
rect 4488 36116 4494 36168
rect 5460 36165 5488 36264
rect 6288 36264 8953 36292
rect 5626 36184 5632 36236
rect 5684 36184 5690 36236
rect 5445 36159 5503 36165
rect 5445 36125 5457 36159
rect 5491 36125 5503 36159
rect 5445 36119 5503 36125
rect 5994 36116 6000 36168
rect 6052 36116 6058 36168
rect 5537 36091 5595 36097
rect 5537 36057 5549 36091
rect 5583 36088 5595 36091
rect 5902 36088 5908 36100
rect 5583 36060 5908 36088
rect 5583 36057 5595 36060
rect 5537 36051 5595 36057
rect 5902 36048 5908 36060
rect 5960 36088 5966 36100
rect 6288 36088 6316 36264
rect 8941 36261 8953 36264
rect 8987 36261 8999 36295
rect 8941 36255 8999 36261
rect 9030 36252 9036 36304
rect 9088 36292 9094 36304
rect 9766 36292 9772 36304
rect 9088 36264 9772 36292
rect 9088 36252 9094 36264
rect 9766 36252 9772 36264
rect 9824 36252 9830 36304
rect 7650 36184 7656 36236
rect 7708 36224 7714 36236
rect 7708 36196 9628 36224
rect 7708 36184 7714 36196
rect 6733 36159 6791 36165
rect 6733 36125 6745 36159
rect 6779 36156 6791 36159
rect 7374 36156 7380 36168
rect 6779 36128 7380 36156
rect 6779 36125 6791 36128
rect 6733 36119 6791 36125
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 7466 36116 7472 36168
rect 7524 36116 7530 36168
rect 8110 36116 8116 36168
rect 8168 36116 8174 36168
rect 9030 36116 9036 36168
rect 9088 36156 9094 36168
rect 9217 36159 9275 36165
rect 9217 36156 9229 36159
rect 9088 36128 9229 36156
rect 9088 36116 9094 36128
rect 9217 36125 9229 36128
rect 9263 36125 9275 36159
rect 9217 36119 9275 36125
rect 9306 36116 9312 36168
rect 9364 36116 9370 36168
rect 9600 36165 9628 36196
rect 10410 36184 10416 36236
rect 10468 36184 10474 36236
rect 11241 36227 11299 36233
rect 11241 36193 11253 36227
rect 11287 36224 11299 36227
rect 11900 36224 11928 36332
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 13354 36320 13360 36372
rect 13412 36320 13418 36372
rect 13906 36320 13912 36372
rect 13964 36320 13970 36372
rect 16206 36360 16212 36372
rect 14292 36332 16212 36360
rect 11287 36196 11928 36224
rect 11287 36193 11299 36196
rect 11241 36187 11299 36193
rect 11974 36184 11980 36236
rect 12032 36184 12038 36236
rect 13924 36224 13952 36320
rect 13188 36196 13952 36224
rect 9401 36159 9459 36165
rect 9401 36125 9413 36159
rect 9447 36125 9459 36159
rect 9401 36119 9459 36125
rect 9585 36159 9643 36165
rect 9585 36125 9597 36159
rect 9631 36125 9643 36159
rect 9585 36119 9643 36125
rect 10229 36159 10287 36165
rect 10229 36125 10241 36159
rect 10275 36156 10287 36159
rect 10275 36128 11008 36156
rect 10275 36125 10287 36128
rect 10229 36119 10287 36125
rect 5960 36060 6316 36088
rect 5960 36048 5966 36060
rect 6914 36048 6920 36100
rect 6972 36088 6978 36100
rect 8021 36091 8079 36097
rect 8021 36088 8033 36091
rect 6972 36060 8033 36088
rect 6972 36048 6978 36060
rect 8021 36057 8033 36060
rect 8067 36057 8079 36091
rect 9416 36088 9444 36119
rect 10980 36100 11008 36128
rect 12066 36116 12072 36168
rect 12124 36116 12130 36168
rect 12244 36159 12302 36165
rect 12244 36125 12256 36159
rect 12290 36156 12302 36159
rect 13188 36156 13216 36196
rect 12290 36128 13216 36156
rect 13633 36159 13691 36165
rect 12290 36125 12302 36128
rect 12244 36119 12302 36125
rect 13633 36125 13645 36159
rect 13679 36156 13691 36159
rect 13814 36156 13820 36168
rect 13679 36128 13820 36156
rect 13679 36125 13691 36128
rect 13633 36119 13691 36125
rect 13814 36116 13820 36128
rect 13872 36116 13878 36168
rect 13909 36159 13967 36165
rect 13909 36125 13921 36159
rect 13955 36156 13967 36159
rect 14292 36156 14320 36332
rect 16206 36320 16212 36332
rect 16264 36320 16270 36372
rect 16850 36320 16856 36372
rect 16908 36360 16914 36372
rect 17310 36360 17316 36372
rect 16908 36332 17316 36360
rect 16908 36320 16914 36332
rect 17310 36320 17316 36332
rect 17368 36320 17374 36372
rect 19242 36320 19248 36372
rect 19300 36320 19306 36372
rect 20254 36320 20260 36372
rect 20312 36320 20318 36372
rect 22462 36320 22468 36372
rect 22520 36320 22526 36372
rect 24489 36363 24547 36369
rect 24489 36329 24501 36363
rect 24535 36360 24547 36363
rect 25866 36360 25872 36372
rect 24535 36332 25872 36360
rect 24535 36329 24547 36332
rect 24489 36323 24547 36329
rect 25866 36320 25872 36332
rect 25924 36320 25930 36372
rect 26602 36320 26608 36372
rect 26660 36320 26666 36372
rect 27525 36363 27583 36369
rect 27525 36329 27537 36363
rect 27571 36360 27583 36363
rect 28074 36360 28080 36372
rect 27571 36332 28080 36360
rect 27571 36329 27583 36332
rect 27525 36323 27583 36329
rect 15105 36295 15163 36301
rect 15105 36261 15117 36295
rect 15151 36292 15163 36295
rect 20272 36292 20300 36320
rect 15151 36264 16712 36292
rect 15151 36261 15163 36264
rect 15105 36255 15163 36261
rect 14734 36184 14740 36236
rect 14792 36184 14798 36236
rect 15654 36184 15660 36236
rect 15712 36184 15718 36236
rect 16684 36233 16712 36264
rect 17880 36264 20300 36292
rect 24121 36295 24179 36301
rect 16669 36227 16727 36233
rect 15764 36196 16252 36224
rect 14553 36159 14611 36165
rect 14553 36156 14565 36159
rect 13955 36128 14320 36156
rect 14384 36128 14565 36156
rect 13955 36125 13967 36128
rect 13909 36119 13967 36125
rect 10134 36088 10140 36100
rect 9416 36060 10140 36088
rect 8021 36051 8079 36057
rect 10134 36048 10140 36060
rect 10192 36048 10198 36100
rect 10962 36048 10968 36100
rect 11020 36048 11026 36100
rect 12084 36088 12112 36116
rect 12084 36060 13124 36088
rect 13096 36032 13124 36060
rect 13722 36048 13728 36100
rect 13780 36088 13786 36100
rect 14384 36088 14412 36128
rect 14553 36125 14565 36128
rect 14599 36156 14611 36159
rect 15565 36159 15623 36165
rect 15565 36156 15577 36159
rect 14599 36128 15577 36156
rect 14599 36125 14611 36128
rect 14553 36119 14611 36125
rect 15565 36125 15577 36128
rect 15611 36156 15623 36159
rect 15764 36156 15792 36196
rect 15611 36128 15792 36156
rect 16025 36159 16083 36165
rect 15611 36125 15623 36128
rect 15565 36119 15623 36125
rect 16025 36125 16037 36159
rect 16071 36156 16083 36159
rect 16114 36156 16120 36168
rect 16071 36128 16120 36156
rect 16071 36125 16083 36128
rect 16025 36119 16083 36125
rect 16114 36116 16120 36128
rect 16172 36116 16178 36168
rect 16224 36156 16252 36196
rect 16669 36193 16681 36227
rect 16715 36193 16727 36227
rect 16669 36187 16727 36193
rect 16942 36184 16948 36236
rect 17000 36184 17006 36236
rect 16960 36156 16988 36184
rect 17589 36159 17647 36165
rect 17589 36156 17601 36159
rect 16224 36128 16988 36156
rect 17052 36128 17601 36156
rect 17052 36100 17080 36128
rect 17589 36125 17601 36128
rect 17635 36125 17647 36159
rect 17589 36119 17647 36125
rect 17681 36159 17739 36165
rect 17681 36125 17693 36159
rect 17727 36156 17739 36159
rect 17770 36156 17776 36168
rect 17727 36128 17776 36156
rect 17727 36125 17739 36128
rect 17681 36119 17739 36125
rect 17770 36116 17776 36128
rect 17828 36116 17834 36168
rect 17880 36165 17908 36264
rect 24121 36261 24133 36295
rect 24167 36261 24179 36295
rect 24121 36255 24179 36261
rect 19797 36227 19855 36233
rect 19797 36193 19809 36227
rect 19843 36193 19855 36227
rect 22094 36224 22100 36236
rect 19797 36187 19855 36193
rect 21468 36196 22100 36224
rect 17865 36159 17923 36165
rect 17865 36125 17877 36159
rect 17911 36125 17923 36159
rect 17865 36119 17923 36125
rect 17954 36116 17960 36168
rect 18012 36116 18018 36168
rect 18506 36116 18512 36168
rect 18564 36116 18570 36168
rect 18598 36116 18604 36168
rect 18656 36156 18662 36168
rect 19705 36159 19763 36165
rect 19705 36156 19717 36159
rect 18656 36128 19717 36156
rect 18656 36116 18662 36128
rect 19705 36125 19717 36128
rect 19751 36125 19763 36159
rect 19705 36119 19763 36125
rect 13780 36060 14412 36088
rect 14461 36091 14519 36097
rect 13780 36048 13786 36060
rect 14461 36057 14473 36091
rect 14507 36088 14519 36091
rect 15378 36088 15384 36100
rect 14507 36060 15384 36088
rect 14507 36057 14519 36060
rect 14461 36051 14519 36057
rect 15378 36048 15384 36060
rect 15436 36048 15442 36100
rect 15473 36091 15531 36097
rect 15473 36057 15485 36091
rect 15519 36088 15531 36091
rect 16577 36091 16635 36097
rect 16577 36088 16589 36091
rect 15519 36060 16589 36088
rect 15519 36057 15531 36060
rect 15473 36051 15531 36057
rect 16577 36057 16589 36060
rect 16623 36057 16635 36091
rect 16577 36051 16635 36057
rect 17034 36048 17040 36100
rect 17092 36048 17098 36100
rect 17494 36048 17500 36100
rect 17552 36088 17558 36100
rect 19812 36088 19840 36187
rect 21468 36168 21496 36196
rect 22094 36184 22100 36196
rect 22152 36224 22158 36236
rect 22741 36227 22799 36233
rect 22741 36224 22753 36227
rect 22152 36196 22753 36224
rect 22152 36184 22158 36196
rect 22741 36193 22753 36196
rect 22787 36193 22799 36227
rect 24136 36224 24164 36255
rect 25590 36252 25596 36304
rect 25648 36292 25654 36304
rect 26620 36292 26648 36320
rect 25648 36264 26480 36292
rect 26620 36264 26924 36292
rect 25648 36252 25654 36264
rect 24302 36224 24308 36236
rect 24136 36196 24308 36224
rect 22741 36187 22799 36193
rect 24302 36184 24308 36196
rect 24360 36224 24366 36236
rect 25869 36227 25927 36233
rect 25869 36224 25881 36227
rect 24360 36196 25881 36224
rect 24360 36184 24366 36196
rect 25869 36193 25881 36196
rect 25915 36224 25927 36227
rect 25958 36224 25964 36236
rect 25915 36196 25964 36224
rect 25915 36193 25927 36196
rect 25869 36187 25927 36193
rect 25958 36184 25964 36196
rect 26016 36184 26022 36236
rect 20257 36159 20315 36165
rect 20257 36156 20269 36159
rect 17552 36060 19840 36088
rect 20180 36128 20269 36156
rect 17552 36048 17558 36060
rect 20180 36032 20208 36128
rect 20257 36125 20269 36128
rect 20303 36156 20315 36159
rect 21450 36156 21456 36168
rect 20303 36128 21456 36156
rect 20303 36125 20315 36128
rect 20257 36119 20315 36125
rect 21450 36116 21456 36128
rect 21508 36116 21514 36168
rect 21818 36116 21824 36168
rect 21876 36116 21882 36168
rect 24673 36159 24731 36165
rect 24673 36125 24685 36159
rect 24719 36156 24731 36159
rect 24762 36156 24768 36168
rect 24719 36128 24768 36156
rect 24719 36125 24731 36128
rect 24673 36119 24731 36125
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 25038 36116 25044 36168
rect 25096 36116 25102 36168
rect 20524 36091 20582 36097
rect 20524 36057 20536 36091
rect 20570 36088 20582 36091
rect 20622 36088 20628 36100
rect 20570 36060 20628 36088
rect 20570 36057 20582 36060
rect 20524 36051 20582 36057
rect 20622 36048 20628 36060
rect 20680 36048 20686 36100
rect 23008 36091 23066 36097
rect 23008 36057 23020 36091
rect 23054 36088 23066 36091
rect 25314 36088 25320 36100
rect 23054 36060 25320 36088
rect 23054 36057 23066 36060
rect 23008 36051 23066 36057
rect 25314 36048 25320 36060
rect 25372 36048 25378 36100
rect 25406 36048 25412 36100
rect 25464 36088 25470 36100
rect 25593 36091 25651 36097
rect 25593 36088 25605 36091
rect 25464 36060 25605 36088
rect 25464 36048 25470 36060
rect 25593 36057 25605 36060
rect 25639 36057 25651 36091
rect 25593 36051 25651 36057
rect 25685 36091 25743 36097
rect 25685 36057 25697 36091
rect 25731 36088 25743 36091
rect 26326 36088 26332 36100
rect 25731 36060 26332 36088
rect 25731 36057 25743 36060
rect 25685 36051 25743 36057
rect 26326 36048 26332 36060
rect 26384 36048 26390 36100
rect 26452 36088 26480 36264
rect 26694 36184 26700 36236
rect 26752 36184 26758 36236
rect 26896 36233 26924 36264
rect 26881 36227 26939 36233
rect 26881 36193 26893 36227
rect 26927 36193 26939 36227
rect 26881 36187 26939 36193
rect 26513 36159 26571 36165
rect 26513 36125 26525 36159
rect 26559 36156 26571 36159
rect 27540 36156 27568 36323
rect 28074 36320 28080 36332
rect 28132 36320 28138 36372
rect 28166 36320 28172 36372
rect 28224 36360 28230 36372
rect 28718 36360 28724 36372
rect 28224 36332 28724 36360
rect 28224 36320 28230 36332
rect 28718 36320 28724 36332
rect 28776 36360 28782 36372
rect 28776 36332 29224 36360
rect 28776 36320 28782 36332
rect 28810 36292 28816 36304
rect 26559 36128 27568 36156
rect 28368 36264 28816 36292
rect 26559 36125 26571 36128
rect 26513 36119 26571 36125
rect 26452 36060 26556 36088
rect 4982 35980 4988 36032
rect 5040 35980 5046 36032
rect 6546 35980 6552 36032
rect 6604 35980 6610 36032
rect 7282 35980 7288 36032
rect 7340 35980 7346 36032
rect 8754 35980 8760 36032
rect 8812 35980 8818 36032
rect 9490 35980 9496 36032
rect 9548 36020 9554 36032
rect 12802 36020 12808 36032
rect 9548 35992 12808 36020
rect 9548 35980 9554 35992
rect 12802 35980 12808 35992
rect 12860 35980 12866 36032
rect 13078 35980 13084 36032
rect 13136 35980 13142 36032
rect 13446 35980 13452 36032
rect 13504 35980 13510 36032
rect 13814 35980 13820 36032
rect 13872 35980 13878 36032
rect 14093 36023 14151 36029
rect 14093 35989 14105 36023
rect 14139 36020 14151 36023
rect 14274 36020 14280 36032
rect 14139 35992 14280 36020
rect 14139 35989 14151 35992
rect 14093 35983 14151 35989
rect 14274 35980 14280 35992
rect 14332 35980 14338 36032
rect 16206 35980 16212 36032
rect 16264 36020 16270 36032
rect 17313 36023 17371 36029
rect 17313 36020 17325 36023
rect 16264 35992 17325 36020
rect 16264 35980 16270 35992
rect 17313 35989 17325 35992
rect 17359 35989 17371 36023
rect 17313 35983 17371 35989
rect 17402 35980 17408 36032
rect 17460 35980 17466 36032
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 18233 36023 18291 36029
rect 18233 36020 18245 36023
rect 18196 35992 18245 36020
rect 18196 35980 18202 35992
rect 18233 35989 18245 35992
rect 18279 35989 18291 36023
rect 18233 35983 18291 35989
rect 19061 36023 19119 36029
rect 19061 35989 19073 36023
rect 19107 36020 19119 36023
rect 19613 36023 19671 36029
rect 19613 36020 19625 36023
rect 19107 35992 19625 36020
rect 19107 35989 19119 35992
rect 19061 35983 19119 35989
rect 19613 35989 19625 35992
rect 19659 35989 19671 36023
rect 19613 35983 19671 35989
rect 20162 35980 20168 36032
rect 20220 35980 20226 36032
rect 21637 36023 21695 36029
rect 21637 35989 21649 36023
rect 21683 36020 21695 36023
rect 21726 36020 21732 36032
rect 21683 35992 21732 36020
rect 21683 35989 21695 35992
rect 21637 35983 21695 35989
rect 21726 35980 21732 35992
rect 21784 35980 21790 36032
rect 25225 36023 25283 36029
rect 25225 35989 25237 36023
rect 25271 36020 25283 36023
rect 25498 36020 25504 36032
rect 25271 35992 25504 36020
rect 25271 35989 25283 35992
rect 25225 35983 25283 35989
rect 25498 35980 25504 35992
rect 25556 35980 25562 36032
rect 26050 35980 26056 36032
rect 26108 35980 26114 36032
rect 26418 35980 26424 36032
rect 26476 35980 26482 36032
rect 26528 36020 26556 36060
rect 26970 36048 26976 36100
rect 27028 36088 27034 36100
rect 28368 36088 28396 36264
rect 28810 36252 28816 36264
rect 28868 36252 28874 36304
rect 28442 36184 28448 36236
rect 28500 36184 28506 36236
rect 28534 36184 28540 36236
rect 28592 36184 28598 36236
rect 28626 36184 28632 36236
rect 28684 36224 28690 36236
rect 28902 36224 28908 36236
rect 28684 36196 28908 36224
rect 28684 36184 28690 36196
rect 28902 36184 28908 36196
rect 28960 36224 28966 36236
rect 29196 36233 29224 36332
rect 29454 36320 29460 36372
rect 29512 36320 29518 36372
rect 29730 36360 29736 36372
rect 29564 36332 29736 36360
rect 28997 36227 29055 36233
rect 28997 36224 29009 36227
rect 28960 36196 29009 36224
rect 28960 36184 28966 36196
rect 28997 36193 29009 36196
rect 29043 36193 29055 36227
rect 28997 36187 29055 36193
rect 29172 36227 29230 36233
rect 29172 36193 29184 36227
rect 29218 36193 29230 36227
rect 29172 36187 29230 36193
rect 29273 36227 29331 36233
rect 29273 36193 29285 36227
rect 29319 36224 29331 36227
rect 29472 36224 29500 36320
rect 29564 36233 29592 36332
rect 29730 36320 29736 36332
rect 29788 36320 29794 36372
rect 29319 36196 29500 36224
rect 29549 36227 29607 36233
rect 29319 36193 29331 36196
rect 29273 36187 29331 36193
rect 29549 36193 29561 36227
rect 29595 36193 29607 36227
rect 29549 36187 29607 36193
rect 32122 36184 32128 36236
rect 32180 36224 32186 36236
rect 33042 36224 33048 36236
rect 32180 36196 33048 36224
rect 32180 36184 32186 36196
rect 33042 36184 33048 36196
rect 33100 36224 33106 36236
rect 33137 36227 33195 36233
rect 33137 36224 33149 36227
rect 33100 36196 33149 36224
rect 33100 36184 33106 36196
rect 33137 36193 33149 36196
rect 33183 36193 33195 36227
rect 33137 36187 33195 36193
rect 29086 36116 29092 36168
rect 29144 36116 29150 36168
rect 30098 36156 30104 36168
rect 29564 36128 30104 36156
rect 27028 36060 28396 36088
rect 27028 36048 27034 36060
rect 27801 36023 27859 36029
rect 27801 36020 27813 36023
rect 26528 35992 27813 36020
rect 27801 35989 27813 35992
rect 27847 36020 27859 36023
rect 27890 36020 27896 36032
rect 27847 35992 27896 36020
rect 27847 35989 27859 35992
rect 27801 35983 27859 35989
rect 27890 35980 27896 35992
rect 27948 35980 27954 36032
rect 27982 35980 27988 36032
rect 28040 35980 28046 36032
rect 28350 35980 28356 36032
rect 28408 35980 28414 36032
rect 28534 35980 28540 36032
rect 28592 36020 28598 36032
rect 28718 36020 28724 36032
rect 28592 35992 28724 36020
rect 28592 35980 28598 35992
rect 28718 35980 28724 35992
rect 28776 35980 28782 36032
rect 28813 36023 28871 36029
rect 28813 35989 28825 36023
rect 28859 36020 28871 36023
rect 29564 36020 29592 36128
rect 30098 36116 30104 36128
rect 30156 36116 30162 36168
rect 30282 36116 30288 36168
rect 30340 36156 30346 36168
rect 31021 36159 31079 36165
rect 31021 36156 31033 36159
rect 30340 36128 31033 36156
rect 30340 36116 30346 36128
rect 31021 36125 31033 36128
rect 31067 36125 31079 36159
rect 31021 36119 31079 36125
rect 29816 36091 29874 36097
rect 29816 36057 29828 36091
rect 29862 36088 29874 36091
rect 31665 36091 31723 36097
rect 31665 36088 31677 36091
rect 29862 36060 30144 36088
rect 29862 36057 29874 36060
rect 29816 36051 29874 36057
rect 28859 35992 29592 36020
rect 30116 36020 30144 36060
rect 30291 36060 31677 36088
rect 30291 36020 30319 36060
rect 31665 36057 31677 36060
rect 31711 36057 31723 36091
rect 31665 36051 31723 36057
rect 32306 36048 32312 36100
rect 32364 36048 32370 36100
rect 30116 35992 30319 36020
rect 28859 35989 28871 35992
rect 28813 35983 28871 35989
rect 30374 35980 30380 36032
rect 30432 36020 30438 36032
rect 30929 36023 30987 36029
rect 30929 36020 30941 36023
rect 30432 35992 30941 36020
rect 30432 35980 30438 35992
rect 30929 35989 30941 35992
rect 30975 35989 30987 36023
rect 30929 35983 30987 35989
rect 31938 35980 31944 36032
rect 31996 35980 32002 36032
rect 32674 35980 32680 36032
rect 32732 35980 32738 36032
rect 1104 35930 43884 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 43884 35930
rect 1104 35856 43884 35878
rect 4430 35776 4436 35828
rect 4488 35816 4494 35828
rect 4617 35819 4675 35825
rect 4617 35816 4629 35819
rect 4488 35788 4629 35816
rect 4488 35776 4494 35788
rect 4617 35785 4629 35788
rect 4663 35785 4675 35819
rect 4617 35779 4675 35785
rect 5994 35776 6000 35828
rect 6052 35816 6058 35828
rect 6365 35819 6423 35825
rect 6365 35816 6377 35819
rect 6052 35788 6377 35816
rect 6052 35776 6058 35788
rect 6365 35785 6377 35788
rect 6411 35785 6423 35819
rect 6365 35779 6423 35785
rect 6733 35819 6791 35825
rect 6733 35785 6745 35819
rect 6779 35816 6791 35819
rect 7282 35816 7288 35828
rect 6779 35788 7288 35816
rect 6779 35785 6791 35788
rect 6733 35779 6791 35785
rect 7282 35776 7288 35788
rect 7340 35776 7346 35828
rect 7374 35776 7380 35828
rect 7432 35776 7438 35828
rect 7466 35776 7472 35828
rect 7524 35816 7530 35828
rect 8021 35819 8079 35825
rect 8021 35816 8033 35819
rect 7524 35788 8033 35816
rect 7524 35776 7530 35788
rect 8021 35785 8033 35788
rect 8067 35785 8079 35819
rect 8021 35779 8079 35785
rect 8110 35776 8116 35828
rect 8168 35776 8174 35828
rect 8389 35819 8447 35825
rect 8389 35785 8401 35819
rect 8435 35816 8447 35819
rect 8754 35816 8760 35828
rect 8435 35788 8760 35816
rect 8435 35785 8447 35788
rect 8389 35779 8447 35785
rect 8754 35776 8760 35788
rect 8812 35776 8818 35828
rect 8849 35819 8907 35825
rect 8849 35785 8861 35819
rect 8895 35816 8907 35819
rect 9398 35816 9404 35828
rect 8895 35788 9404 35816
rect 8895 35785 8907 35788
rect 8849 35779 8907 35785
rect 9398 35776 9404 35788
rect 9456 35776 9462 35828
rect 12526 35776 12532 35828
rect 12584 35776 12590 35828
rect 12618 35776 12624 35828
rect 12676 35776 12682 35828
rect 12989 35819 13047 35825
rect 12989 35785 13001 35819
rect 13035 35816 13047 35819
rect 13170 35816 13176 35828
rect 13035 35788 13176 35816
rect 13035 35785 13047 35788
rect 12989 35779 13047 35785
rect 13170 35776 13176 35788
rect 13228 35776 13234 35828
rect 13722 35776 13728 35828
rect 13780 35776 13786 35828
rect 13814 35776 13820 35828
rect 13872 35816 13878 35828
rect 16390 35816 16396 35828
rect 13872 35788 16396 35816
rect 13872 35776 13878 35788
rect 16390 35776 16396 35788
rect 16448 35776 16454 35828
rect 18322 35776 18328 35828
rect 18380 35776 18386 35828
rect 18506 35816 18512 35828
rect 18432 35788 18512 35816
rect 5626 35748 5632 35760
rect 3988 35720 5632 35748
rect 3988 35689 4016 35720
rect 5626 35708 5632 35720
rect 5684 35748 5690 35760
rect 5813 35751 5871 35757
rect 5813 35748 5825 35751
rect 5684 35720 5825 35748
rect 5684 35708 5690 35720
rect 5813 35717 5825 35720
rect 5859 35717 5871 35751
rect 7392 35748 7420 35776
rect 7561 35751 7619 35757
rect 7561 35748 7573 35751
rect 5813 35711 5871 35717
rect 6288 35720 6960 35748
rect 7392 35720 7573 35748
rect 3973 35683 4031 35689
rect 3973 35649 3985 35683
rect 4019 35649 4031 35683
rect 3973 35643 4031 35649
rect 4525 35683 4583 35689
rect 4525 35649 4537 35683
rect 4571 35680 4583 35683
rect 4985 35683 5043 35689
rect 4985 35680 4997 35683
rect 4571 35652 4997 35680
rect 4571 35649 4583 35652
rect 4525 35643 4583 35649
rect 4985 35649 4997 35652
rect 5031 35649 5043 35683
rect 4985 35643 5043 35649
rect 5077 35615 5135 35621
rect 5077 35581 5089 35615
rect 5123 35581 5135 35615
rect 5077 35575 5135 35581
rect 5092 35544 5120 35575
rect 5258 35572 5264 35624
rect 5316 35572 5322 35624
rect 5902 35572 5908 35624
rect 5960 35572 5966 35624
rect 6089 35615 6147 35621
rect 6089 35581 6101 35615
rect 6135 35612 6147 35615
rect 6288 35612 6316 35720
rect 6825 35683 6883 35689
rect 6825 35649 6837 35683
rect 6871 35649 6883 35683
rect 6932 35680 6960 35720
rect 7561 35717 7573 35720
rect 7607 35717 7619 35751
rect 7561 35711 7619 35717
rect 7653 35751 7711 35757
rect 7653 35717 7665 35751
rect 7699 35748 7711 35751
rect 7742 35748 7748 35760
rect 7699 35720 7748 35748
rect 7699 35717 7711 35720
rect 7653 35711 7711 35717
rect 7742 35708 7748 35720
rect 7800 35748 7806 35760
rect 8128 35748 8156 35776
rect 7800 35720 8156 35748
rect 7800 35708 7806 35720
rect 8294 35708 8300 35760
rect 8352 35748 8358 35760
rect 10134 35748 10140 35760
rect 8352 35720 9260 35748
rect 8352 35708 8358 35720
rect 8864 35692 8892 35720
rect 6932 35652 7880 35680
rect 6825 35643 6883 35649
rect 6135 35584 6316 35612
rect 6135 35581 6147 35584
rect 6089 35575 6147 35581
rect 6270 35544 6276 35556
rect 5092 35516 6276 35544
rect 6270 35504 6276 35516
rect 6328 35544 6334 35556
rect 6840 35544 6868 35643
rect 7006 35572 7012 35624
rect 7064 35572 7070 35624
rect 7852 35621 7880 35652
rect 8846 35640 8852 35692
rect 8904 35640 8910 35692
rect 9030 35640 9036 35692
rect 9088 35680 9094 35692
rect 9232 35689 9260 35720
rect 9416 35720 10140 35748
rect 9125 35683 9183 35689
rect 9125 35680 9137 35683
rect 9088 35652 9137 35680
rect 9088 35640 9094 35652
rect 9125 35649 9137 35652
rect 9171 35649 9183 35683
rect 9125 35643 9183 35649
rect 9217 35683 9275 35689
rect 9217 35649 9229 35683
rect 9263 35649 9275 35683
rect 9217 35643 9275 35649
rect 9314 35683 9372 35689
rect 9314 35649 9326 35683
rect 9360 35680 9372 35683
rect 9416 35680 9444 35720
rect 10134 35708 10140 35720
rect 10192 35708 10198 35760
rect 11330 35708 11336 35760
rect 11388 35748 11394 35760
rect 11793 35751 11851 35757
rect 11793 35748 11805 35751
rect 11388 35720 11805 35748
rect 11388 35708 11394 35720
rect 11793 35717 11805 35720
rect 11839 35748 11851 35751
rect 11839 35720 12680 35748
rect 11839 35717 11851 35720
rect 11793 35711 11851 35717
rect 9360 35652 9444 35680
rect 9493 35683 9551 35689
rect 9360 35649 9372 35652
rect 9314 35643 9372 35649
rect 9493 35649 9505 35683
rect 9539 35649 9551 35683
rect 9493 35643 9551 35649
rect 9585 35683 9643 35689
rect 9585 35649 9597 35683
rect 9631 35680 9643 35683
rect 9674 35680 9680 35692
rect 9631 35652 9680 35680
rect 9631 35649 9643 35652
rect 9585 35643 9643 35649
rect 7837 35615 7895 35621
rect 7837 35581 7849 35615
rect 7883 35612 7895 35615
rect 8018 35612 8024 35624
rect 7883 35584 8024 35612
rect 7883 35581 7895 35584
rect 7837 35575 7895 35581
rect 8018 35572 8024 35584
rect 8076 35572 8082 35624
rect 8481 35615 8539 35621
rect 8481 35581 8493 35615
rect 8527 35581 8539 35615
rect 8481 35575 8539 35581
rect 8665 35615 8723 35621
rect 8665 35581 8677 35615
rect 8711 35612 8723 35615
rect 9398 35612 9404 35624
rect 8711 35584 9404 35612
rect 8711 35581 8723 35584
rect 8665 35575 8723 35581
rect 8496 35544 8524 35575
rect 9398 35572 9404 35584
rect 9456 35572 9462 35624
rect 9508 35612 9536 35643
rect 9674 35640 9680 35652
rect 9732 35640 9738 35692
rect 9766 35640 9772 35692
rect 9824 35680 9830 35692
rect 9824 35652 10548 35680
rect 9824 35640 9830 35652
rect 9508 35584 9904 35612
rect 6328 35516 9628 35544
rect 6328 35504 6334 35516
rect 9600 35488 9628 35516
rect 9876 35488 9904 35584
rect 10520 35488 10548 35652
rect 11146 35640 11152 35692
rect 11204 35640 11210 35692
rect 11882 35640 11888 35692
rect 11940 35640 11946 35692
rect 12652 35680 12680 35720
rect 12710 35708 12716 35760
rect 12768 35748 12774 35760
rect 13081 35751 13139 35757
rect 13081 35748 13093 35751
rect 12768 35720 13093 35748
rect 12768 35708 12774 35720
rect 13081 35717 13093 35720
rect 13127 35748 13139 35751
rect 13740 35748 13768 35776
rect 13127 35720 13768 35748
rect 14553 35751 14611 35757
rect 13127 35717 13139 35720
rect 13081 35711 13139 35717
rect 14553 35717 14565 35751
rect 14599 35748 14611 35751
rect 14642 35748 14648 35760
rect 14599 35720 14648 35748
rect 14599 35717 14611 35720
rect 14553 35711 14611 35717
rect 14642 35708 14648 35720
rect 14700 35748 14706 35760
rect 15004 35751 15062 35757
rect 14700 35720 14780 35748
rect 14700 35708 14706 35720
rect 13725 35683 13783 35689
rect 13725 35680 13737 35683
rect 12652 35652 13737 35680
rect 13725 35649 13737 35652
rect 13771 35680 13783 35683
rect 13998 35680 14004 35692
rect 13771 35652 14004 35680
rect 13771 35649 13783 35652
rect 13725 35643 13783 35649
rect 13998 35640 14004 35652
rect 14056 35640 14062 35692
rect 14752 35689 14780 35720
rect 15004 35717 15016 35751
rect 15050 35748 15062 35751
rect 16206 35748 16212 35760
rect 15050 35720 16212 35748
rect 15050 35717 15062 35720
rect 15004 35711 15062 35717
rect 16206 35708 16212 35720
rect 16264 35708 16270 35760
rect 17681 35751 17739 35757
rect 17681 35717 17693 35751
rect 17727 35717 17739 35751
rect 18340 35748 18368 35776
rect 18432 35757 18460 35788
rect 18506 35776 18512 35788
rect 18564 35816 18570 35828
rect 19889 35819 19947 35825
rect 19889 35816 19901 35819
rect 18564 35788 19901 35816
rect 18564 35776 18570 35788
rect 19889 35785 19901 35788
rect 19935 35785 19947 35819
rect 19889 35779 19947 35785
rect 21545 35819 21603 35825
rect 21545 35785 21557 35819
rect 21591 35816 21603 35819
rect 21818 35816 21824 35828
rect 21591 35788 21824 35816
rect 21591 35785 21603 35788
rect 21545 35779 21603 35785
rect 21818 35776 21824 35788
rect 21876 35776 21882 35828
rect 23198 35776 23204 35828
rect 23256 35776 23262 35828
rect 23750 35776 23756 35828
rect 23808 35776 23814 35828
rect 25317 35819 25375 35825
rect 25317 35785 25329 35819
rect 25363 35816 25375 35819
rect 25406 35816 25412 35828
rect 25363 35788 25412 35816
rect 25363 35785 25375 35788
rect 25317 35779 25375 35785
rect 25406 35776 25412 35788
rect 25464 35776 25470 35828
rect 25685 35819 25743 35825
rect 25685 35785 25697 35819
rect 25731 35816 25743 35819
rect 25774 35816 25780 35828
rect 25731 35788 25780 35816
rect 25731 35785 25743 35788
rect 25685 35779 25743 35785
rect 25774 35776 25780 35788
rect 25832 35776 25838 35828
rect 26050 35776 26056 35828
rect 26108 35776 26114 35828
rect 26510 35776 26516 35828
rect 26568 35776 26574 35828
rect 26694 35776 26700 35828
rect 26752 35816 26758 35828
rect 28629 35819 28687 35825
rect 26752 35788 28580 35816
rect 26752 35776 26758 35788
rect 17681 35711 17739 35717
rect 18064 35720 18368 35748
rect 18417 35751 18475 35757
rect 14737 35683 14795 35689
rect 14737 35649 14749 35683
rect 14783 35649 14795 35683
rect 14737 35643 14795 35649
rect 14826 35640 14832 35692
rect 14884 35680 14890 35692
rect 17696 35680 17724 35711
rect 14884 35652 17724 35680
rect 17865 35683 17923 35689
rect 14884 35640 14890 35652
rect 17865 35649 17877 35683
rect 17911 35680 17923 35683
rect 18064 35680 18092 35720
rect 18417 35717 18429 35751
rect 18463 35717 18475 35751
rect 20432 35751 20490 35757
rect 18417 35711 18475 35717
rect 18524 35720 19840 35748
rect 17911 35652 18092 35680
rect 18141 35683 18199 35689
rect 17911 35649 17923 35652
rect 17865 35643 17923 35649
rect 18141 35649 18153 35683
rect 18187 35680 18199 35683
rect 18322 35680 18328 35692
rect 18187 35652 18328 35680
rect 18187 35649 18199 35652
rect 18141 35643 18199 35649
rect 18322 35640 18328 35652
rect 18380 35640 18386 35692
rect 10965 35615 11023 35621
rect 10965 35581 10977 35615
rect 11011 35612 11023 35615
rect 11422 35612 11428 35624
rect 11011 35584 11428 35612
rect 11011 35581 11023 35584
rect 10965 35575 11023 35581
rect 11422 35572 11428 35584
rect 11480 35572 11486 35624
rect 13262 35572 13268 35624
rect 13320 35572 13326 35624
rect 16942 35572 16948 35624
rect 17000 35572 17006 35624
rect 17497 35615 17555 35621
rect 17497 35581 17509 35615
rect 17543 35581 17555 35615
rect 17497 35575 17555 35581
rect 10873 35547 10931 35553
rect 10873 35513 10885 35547
rect 10919 35544 10931 35547
rect 11606 35544 11612 35556
rect 10919 35516 11612 35544
rect 10919 35513 10931 35516
rect 10873 35507 10931 35513
rect 11606 35504 11612 35516
rect 11664 35504 11670 35556
rect 12802 35504 12808 35556
rect 12860 35544 12866 35556
rect 13814 35544 13820 35556
rect 12860 35516 13820 35544
rect 12860 35504 12866 35516
rect 13814 35504 13820 35516
rect 13872 35544 13878 35556
rect 14182 35544 14188 35556
rect 13872 35516 14188 35544
rect 13872 35504 13878 35516
rect 14182 35504 14188 35516
rect 14240 35504 14246 35556
rect 16574 35504 16580 35556
rect 16632 35544 16638 35556
rect 17512 35544 17540 35575
rect 17678 35572 17684 35624
rect 17736 35612 17742 35624
rect 18524 35621 18552 35720
rect 18776 35683 18834 35689
rect 18776 35649 18788 35683
rect 18822 35680 18834 35683
rect 19334 35680 19340 35692
rect 18822 35652 19340 35680
rect 18822 35649 18834 35652
rect 18776 35643 18834 35649
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 19812 35680 19840 35720
rect 20432 35717 20444 35751
rect 20478 35748 20490 35751
rect 20530 35748 20536 35760
rect 20478 35720 20536 35748
rect 20478 35717 20490 35720
rect 20432 35711 20490 35717
rect 20530 35708 20536 35720
rect 20588 35708 20594 35760
rect 22088 35751 22146 35757
rect 22088 35717 22100 35751
rect 22134 35748 22146 35751
rect 23566 35748 23572 35760
rect 22134 35720 23572 35748
rect 22134 35717 22146 35720
rect 22088 35711 22146 35717
rect 23566 35708 23572 35720
rect 23624 35708 23630 35760
rect 24486 35708 24492 35760
rect 24544 35748 24550 35760
rect 24544 35720 25820 35748
rect 24544 35708 24550 35720
rect 20162 35680 20168 35692
rect 19812 35652 20168 35680
rect 20162 35640 20168 35652
rect 20220 35640 20226 35692
rect 21450 35640 21456 35692
rect 21508 35680 21514 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21508 35652 21833 35680
rect 21508 35640 21514 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 23661 35683 23719 35689
rect 23661 35680 23673 35683
rect 21821 35643 21879 35649
rect 23492 35652 23673 35680
rect 23492 35624 23520 35652
rect 23661 35649 23673 35652
rect 23707 35649 23719 35683
rect 24302 35680 24308 35692
rect 23661 35643 23719 35649
rect 23952 35652 24308 35680
rect 18509 35615 18567 35621
rect 18509 35612 18521 35615
rect 17736 35584 18521 35612
rect 17736 35572 17742 35584
rect 18509 35581 18521 35584
rect 18555 35581 18567 35615
rect 18509 35575 18567 35581
rect 23474 35572 23480 35624
rect 23532 35572 23538 35624
rect 23952 35621 23980 35652
rect 24302 35640 24308 35652
rect 24360 35640 24366 35692
rect 24394 35640 24400 35692
rect 24452 35680 24458 35692
rect 24452 35652 25084 35680
rect 24452 35640 24458 35652
rect 23937 35615 23995 35621
rect 23937 35581 23949 35615
rect 23983 35581 23995 35615
rect 23937 35575 23995 35581
rect 24670 35572 24676 35624
rect 24728 35612 24734 35624
rect 24949 35615 25007 35621
rect 24949 35612 24961 35615
rect 24728 35584 24961 35612
rect 24728 35572 24734 35584
rect 24949 35581 24961 35584
rect 24995 35581 25007 35615
rect 25056 35612 25084 35652
rect 25130 35640 25136 35692
rect 25188 35640 25194 35692
rect 25501 35683 25559 35689
rect 25501 35680 25513 35683
rect 25231 35652 25513 35680
rect 25231 35612 25259 35652
rect 25501 35649 25513 35652
rect 25547 35680 25559 35683
rect 25590 35680 25596 35692
rect 25547 35652 25596 35680
rect 25547 35649 25559 35652
rect 25501 35643 25559 35649
rect 25590 35640 25596 35652
rect 25648 35640 25654 35692
rect 25792 35689 25820 35720
rect 26068 35689 26096 35776
rect 26528 35748 26556 35776
rect 27433 35751 27491 35757
rect 27433 35748 27445 35751
rect 26528 35720 27445 35748
rect 27433 35717 27445 35720
rect 27479 35717 27491 35751
rect 27433 35711 27491 35717
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35649 25835 35683
rect 25777 35643 25835 35649
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35649 26111 35683
rect 26053 35643 26111 35649
rect 27249 35683 27307 35689
rect 27249 35649 27261 35683
rect 27295 35680 27307 35683
rect 27338 35680 27344 35692
rect 27295 35652 27344 35680
rect 27295 35649 27307 35652
rect 27249 35643 27307 35649
rect 27338 35640 27344 35652
rect 27396 35640 27402 35692
rect 27448 35680 27476 35711
rect 28258 35680 28264 35692
rect 27448 35652 28264 35680
rect 28258 35640 28264 35652
rect 28316 35640 28322 35692
rect 28445 35683 28503 35689
rect 28445 35649 28457 35683
rect 28491 35649 28503 35683
rect 28445 35643 28503 35649
rect 25056 35584 25259 35612
rect 24949 35575 25007 35581
rect 25314 35572 25320 35624
rect 25372 35572 25378 35624
rect 25869 35615 25927 35621
rect 25869 35581 25881 35615
rect 25915 35612 25927 35615
rect 26605 35615 26663 35621
rect 26605 35612 26617 35615
rect 25915 35584 26617 35612
rect 25915 35581 25927 35584
rect 25869 35575 25927 35581
rect 26605 35581 26617 35584
rect 26651 35612 26663 35615
rect 26786 35612 26792 35624
rect 26651 35584 26792 35612
rect 26651 35581 26663 35584
rect 26605 35575 26663 35581
rect 16632 35516 17540 35544
rect 17589 35547 17647 35553
rect 16632 35504 16638 35516
rect 17589 35513 17601 35547
rect 17635 35544 17647 35547
rect 17862 35544 17868 35556
rect 17635 35516 17868 35544
rect 17635 35513 17647 35516
rect 17589 35507 17647 35513
rect 17862 35504 17868 35516
rect 17920 35544 17926 35556
rect 23293 35547 23351 35553
rect 17920 35516 18258 35544
rect 17920 35504 17926 35516
rect 5445 35479 5503 35485
rect 5445 35445 5457 35479
rect 5491 35476 5503 35479
rect 6454 35476 6460 35488
rect 5491 35448 6460 35476
rect 5491 35445 5503 35448
rect 5445 35439 5503 35445
rect 6454 35436 6460 35448
rect 6512 35436 6518 35488
rect 7190 35436 7196 35488
rect 7248 35436 7254 35488
rect 9582 35436 9588 35488
rect 9640 35436 9646 35488
rect 9858 35436 9864 35488
rect 9916 35436 9922 35488
rect 9950 35436 9956 35488
rect 10008 35436 10014 35488
rect 10502 35436 10508 35488
rect 10560 35436 10566 35488
rect 11333 35479 11391 35485
rect 11333 35445 11345 35479
rect 11379 35476 11391 35479
rect 12342 35476 12348 35488
rect 11379 35448 12348 35476
rect 11379 35445 11391 35448
rect 11333 35439 11391 35445
rect 12342 35436 12348 35448
rect 12400 35476 12406 35488
rect 12986 35476 12992 35488
rect 12400 35448 12992 35476
rect 12400 35436 12406 35448
rect 12986 35436 12992 35448
rect 13044 35436 13050 35488
rect 16114 35436 16120 35488
rect 16172 35436 16178 35488
rect 16485 35479 16543 35485
rect 16485 35445 16497 35479
rect 16531 35476 16543 35479
rect 18138 35476 18144 35488
rect 16531 35448 18144 35476
rect 16531 35445 16543 35448
rect 16485 35439 16543 35445
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 18230 35476 18258 35516
rect 23293 35513 23305 35547
rect 23339 35544 23351 35547
rect 25130 35544 25136 35556
rect 23339 35516 25136 35544
rect 23339 35513 23351 35516
rect 23293 35507 23351 35513
rect 25130 35504 25136 35516
rect 25188 35504 25194 35556
rect 25332 35544 25360 35572
rect 25501 35547 25559 35553
rect 25501 35544 25513 35547
rect 25332 35516 25513 35544
rect 25501 35513 25513 35516
rect 25547 35513 25559 35547
rect 25501 35507 25559 35513
rect 19150 35476 19156 35488
rect 18230 35448 19156 35476
rect 19150 35436 19156 35448
rect 19208 35436 19214 35488
rect 24854 35436 24860 35488
rect 24912 35436 24918 35488
rect 25222 35436 25228 35488
rect 25280 35476 25286 35488
rect 25884 35476 25912 35575
rect 26786 35572 26792 35584
rect 26844 35572 26850 35624
rect 27065 35615 27123 35621
rect 27065 35581 27077 35615
rect 27111 35581 27123 35615
rect 27065 35575 27123 35581
rect 26142 35504 26148 35556
rect 26200 35544 26206 35556
rect 27080 35544 27108 35575
rect 27154 35572 27160 35624
rect 27212 35612 27218 35624
rect 27525 35615 27583 35621
rect 27525 35612 27537 35615
rect 27212 35584 27537 35612
rect 27212 35572 27218 35584
rect 27525 35581 27537 35584
rect 27571 35581 27583 35615
rect 27525 35575 27583 35581
rect 28166 35572 28172 35624
rect 28224 35572 28230 35624
rect 28184 35544 28212 35572
rect 26200 35516 28212 35544
rect 28460 35544 28488 35643
rect 28552 35612 28580 35788
rect 28629 35785 28641 35819
rect 28675 35816 28687 35819
rect 29178 35816 29184 35828
rect 28675 35788 29184 35816
rect 28675 35785 28687 35788
rect 28629 35779 28687 35785
rect 29178 35776 29184 35788
rect 29236 35776 29242 35828
rect 29270 35776 29276 35828
rect 29328 35776 29334 35828
rect 29730 35776 29736 35828
rect 29788 35776 29794 35828
rect 33042 35776 33048 35828
rect 33100 35776 33106 35828
rect 29086 35708 29092 35760
rect 29144 35708 29150 35760
rect 29748 35748 29776 35776
rect 29748 35720 30512 35748
rect 28994 35640 29000 35692
rect 29052 35680 29058 35692
rect 29641 35683 29699 35689
rect 29641 35680 29653 35683
rect 29052 35652 29653 35680
rect 29052 35640 29058 35652
rect 29641 35649 29653 35652
rect 29687 35649 29699 35683
rect 29641 35643 29699 35649
rect 30374 35640 30380 35692
rect 30432 35640 30438 35692
rect 30484 35689 30512 35720
rect 31018 35708 31024 35760
rect 31076 35748 31082 35760
rect 32769 35751 32827 35757
rect 32769 35748 32781 35751
rect 31076 35720 32781 35748
rect 31076 35708 31082 35720
rect 32769 35717 32781 35720
rect 32815 35717 32827 35751
rect 32769 35711 32827 35717
rect 30469 35683 30527 35689
rect 30469 35649 30481 35683
rect 30515 35649 30527 35683
rect 30469 35643 30527 35649
rect 30736 35683 30794 35689
rect 30736 35649 30748 35683
rect 30782 35680 30794 35683
rect 32214 35680 32220 35692
rect 30782 35652 32220 35680
rect 30782 35649 30794 35652
rect 30736 35643 30794 35649
rect 32214 35640 32220 35652
rect 32272 35640 32278 35692
rect 29365 35615 29423 35621
rect 29365 35612 29377 35615
rect 28552 35584 29377 35612
rect 29365 35581 29377 35584
rect 29411 35581 29423 35615
rect 29365 35575 29423 35581
rect 29549 35615 29607 35621
rect 29549 35581 29561 35615
rect 29595 35612 29607 35615
rect 29730 35612 29736 35624
rect 29595 35584 29736 35612
rect 29595 35581 29607 35584
rect 29549 35575 29607 35581
rect 29730 35572 29736 35584
rect 29788 35612 29794 35624
rect 30282 35612 30288 35624
rect 29788 35584 30288 35612
rect 29788 35572 29794 35584
rect 30282 35572 30288 35584
rect 30340 35572 30346 35624
rect 28902 35544 28908 35556
rect 28460 35516 28908 35544
rect 26200 35504 26206 35516
rect 28902 35504 28908 35516
rect 28960 35544 28966 35556
rect 30392 35544 30420 35640
rect 32125 35615 32183 35621
rect 32125 35612 32137 35615
rect 31864 35584 32137 35612
rect 31864 35553 31892 35584
rect 32125 35581 32137 35584
rect 32171 35581 32183 35615
rect 32125 35575 32183 35581
rect 28960 35516 30420 35544
rect 31849 35547 31907 35553
rect 28960 35504 28966 35516
rect 31849 35513 31861 35547
rect 31895 35513 31907 35547
rect 31849 35507 31907 35513
rect 25958 35476 25964 35488
rect 25280 35448 25964 35476
rect 25280 35436 25286 35448
rect 25958 35436 25964 35448
rect 26016 35436 26022 35488
rect 26234 35436 26240 35488
rect 26292 35436 26298 35488
rect 28166 35436 28172 35488
rect 28224 35436 28230 35488
rect 28810 35436 28816 35488
rect 28868 35436 28874 35488
rect 29086 35436 29092 35488
rect 29144 35476 29150 35488
rect 29825 35479 29883 35485
rect 29825 35476 29837 35479
rect 29144 35448 29837 35476
rect 29144 35436 29150 35448
rect 29825 35445 29837 35448
rect 29871 35445 29883 35479
rect 29825 35439 29883 35445
rect 30098 35436 30104 35488
rect 30156 35476 30162 35488
rect 31754 35476 31760 35488
rect 30156 35448 31760 35476
rect 30156 35436 30162 35448
rect 31754 35436 31760 35448
rect 31812 35436 31818 35488
rect 1104 35386 43884 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 43884 35386
rect 1104 35312 43884 35334
rect 3605 35275 3663 35281
rect 3605 35241 3617 35275
rect 3651 35272 3663 35275
rect 3651 35244 5580 35272
rect 3651 35241 3663 35244
rect 3605 35235 3663 35241
rect 5552 35204 5580 35244
rect 5626 35232 5632 35284
rect 5684 35232 5690 35284
rect 6086 35272 6092 35284
rect 5736 35244 6092 35272
rect 5736 35204 5764 35244
rect 6086 35232 6092 35244
rect 6144 35272 6150 35284
rect 7101 35275 7159 35281
rect 6144 35244 7052 35272
rect 6144 35232 6150 35244
rect 5552 35176 5764 35204
rect 7024 35204 7052 35244
rect 7101 35241 7113 35275
rect 7147 35272 7159 35275
rect 7374 35272 7380 35284
rect 7147 35244 7380 35272
rect 7147 35241 7159 35244
rect 7101 35235 7159 35241
rect 7374 35232 7380 35244
rect 7432 35232 7438 35284
rect 8662 35232 8668 35284
rect 8720 35272 8726 35284
rect 9585 35275 9643 35281
rect 9585 35272 9597 35275
rect 8720 35244 9597 35272
rect 8720 35232 8726 35244
rect 9585 35241 9597 35244
rect 9631 35241 9643 35275
rect 9585 35235 9643 35241
rect 9858 35232 9864 35284
rect 9916 35272 9922 35284
rect 10413 35275 10471 35281
rect 10413 35272 10425 35275
rect 9916 35244 10425 35272
rect 9916 35232 9922 35244
rect 10413 35241 10425 35244
rect 10459 35241 10471 35275
rect 10413 35235 10471 35241
rect 10597 35275 10655 35281
rect 10597 35241 10609 35275
rect 10643 35272 10655 35275
rect 11146 35272 11152 35284
rect 10643 35244 11152 35272
rect 10643 35241 10655 35244
rect 10597 35235 10655 35241
rect 11146 35232 11152 35244
rect 11204 35232 11210 35284
rect 11425 35275 11483 35281
rect 11425 35241 11437 35275
rect 11471 35272 11483 35275
rect 11698 35272 11704 35284
rect 11471 35244 11704 35272
rect 11471 35241 11483 35244
rect 11425 35235 11483 35241
rect 11698 35232 11704 35244
rect 11756 35232 11762 35284
rect 12710 35232 12716 35284
rect 12768 35232 12774 35284
rect 12802 35232 12808 35284
rect 12860 35272 12866 35284
rect 12897 35275 12955 35281
rect 12897 35272 12909 35275
rect 12860 35244 12909 35272
rect 12860 35232 12866 35244
rect 12897 35241 12909 35244
rect 12943 35241 12955 35275
rect 12897 35235 12955 35241
rect 12986 35232 12992 35284
rect 13044 35272 13050 35284
rect 13909 35275 13967 35281
rect 13044 35244 13584 35272
rect 13044 35232 13050 35244
rect 7469 35207 7527 35213
rect 7469 35204 7481 35207
rect 7024 35176 7481 35204
rect 7469 35173 7481 35176
rect 7515 35173 7527 35207
rect 7469 35167 7527 35173
rect 7484 35136 7512 35167
rect 7650 35164 7656 35216
rect 7708 35164 7714 35216
rect 9030 35204 9036 35216
rect 7760 35176 9036 35204
rect 7760 35136 7788 35176
rect 9030 35164 9036 35176
rect 9088 35164 9094 35216
rect 11330 35204 11336 35216
rect 9140 35176 11336 35204
rect 7484 35108 7788 35136
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1581 35071 1639 35077
rect 1581 35068 1593 35071
rect 992 35040 1593 35068
rect 992 35028 998 35040
rect 1581 35037 1593 35040
rect 1627 35037 1639 35071
rect 1581 35031 1639 35037
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35068 4307 35071
rect 5721 35071 5779 35077
rect 5721 35068 5733 35071
rect 4295 35040 5733 35068
rect 4295 35037 4307 35040
rect 4249 35031 4307 35037
rect 5721 35037 5733 35040
rect 5767 35068 5779 35071
rect 7006 35068 7012 35080
rect 5767 35040 7012 35068
rect 5767 35037 5779 35040
rect 5721 35031 5779 35037
rect 7006 35028 7012 35040
rect 7064 35028 7070 35080
rect 7558 35028 7564 35080
rect 7616 35028 7622 35080
rect 7668 35070 7696 35108
rect 8570 35096 8576 35148
rect 8628 35096 8634 35148
rect 8938 35096 8944 35148
rect 8996 35096 9002 35148
rect 7745 35071 7803 35077
rect 7745 35070 7757 35071
rect 7668 35042 7757 35070
rect 7745 35037 7757 35042
rect 7791 35037 7803 35071
rect 7745 35031 7803 35037
rect 4516 35003 4574 35009
rect 4516 34969 4528 35003
rect 4562 35000 4574 35003
rect 4982 35000 4988 35012
rect 4562 34972 4988 35000
rect 4562 34969 4574 34972
rect 4516 34963 4574 34969
rect 4982 34960 4988 34972
rect 5040 34960 5046 35012
rect 5988 35003 6046 35009
rect 5988 34969 6000 35003
rect 6034 35000 6046 35003
rect 6546 35000 6552 35012
rect 6034 34972 6552 35000
rect 6034 34969 6046 34972
rect 5988 34963 6046 34969
rect 6546 34960 6552 34972
rect 6604 34960 6610 35012
rect 6822 34960 6828 35012
rect 6880 35000 6886 35012
rect 7837 35003 7895 35009
rect 7837 35000 7849 35003
rect 6880 34972 7849 35000
rect 6880 34960 6886 34972
rect 7837 34969 7849 34972
rect 7883 35000 7895 35003
rect 9140 35000 9168 35176
rect 11330 35164 11336 35176
rect 11388 35164 11394 35216
rect 12618 35164 12624 35216
rect 12676 35164 12682 35216
rect 13354 35204 13360 35216
rect 12820 35176 13360 35204
rect 9766 35096 9772 35148
rect 9824 35096 9830 35148
rect 11241 35139 11299 35145
rect 11241 35105 11253 35139
rect 11287 35136 11299 35139
rect 11287 35108 11321 35136
rect 11287 35105 11299 35108
rect 11241 35099 11299 35105
rect 9214 35028 9220 35080
rect 9272 35068 9278 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9272 35040 9873 35068
rect 9272 35028 9278 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 10318 35028 10324 35080
rect 10376 35028 10382 35080
rect 10502 35028 10508 35080
rect 10560 35068 10566 35080
rect 10870 35068 10876 35080
rect 10560 35040 10876 35068
rect 10560 35028 10566 35040
rect 10870 35028 10876 35040
rect 10928 35068 10934 35080
rect 11256 35068 11284 35099
rect 11422 35096 11428 35148
rect 11480 35136 11486 35148
rect 12636 35136 12664 35164
rect 11480 35108 12664 35136
rect 11480 35096 11486 35108
rect 11701 35071 11759 35077
rect 11701 35068 11713 35071
rect 10928 35040 11713 35068
rect 10928 35028 10934 35040
rect 11701 35037 11713 35040
rect 11747 35037 11759 35071
rect 11701 35031 11759 35037
rect 11790 35028 11796 35080
rect 11848 35028 11854 35080
rect 11900 35077 11928 35108
rect 12820 35077 12848 35176
rect 13354 35164 13360 35176
rect 13412 35164 13418 35216
rect 13081 35139 13139 35145
rect 13081 35105 13093 35139
rect 13127 35136 13139 35139
rect 13446 35136 13452 35148
rect 13127 35108 13452 35136
rect 13127 35105 13139 35108
rect 13081 35099 13139 35105
rect 13446 35096 13452 35108
rect 13504 35096 13510 35148
rect 11885 35071 11943 35077
rect 11885 35037 11897 35071
rect 11931 35037 11943 35071
rect 11885 35031 11943 35037
rect 12069 35071 12127 35077
rect 12069 35037 12081 35071
rect 12115 35037 12127 35071
rect 12069 35031 12127 35037
rect 12805 35071 12863 35077
rect 12805 35037 12817 35071
rect 12851 35037 12863 35071
rect 12805 35031 12863 35037
rect 11057 35003 11115 35009
rect 11057 35000 11069 35003
rect 7883 34972 9168 35000
rect 10244 34972 11069 35000
rect 7883 34969 7895 34972
rect 7837 34963 7895 34969
rect 3237 34935 3295 34941
rect 3237 34901 3249 34935
rect 3283 34932 3295 34935
rect 3326 34932 3332 34944
rect 3283 34904 3332 34932
rect 3283 34901 3295 34904
rect 3237 34895 3295 34901
rect 3326 34892 3332 34904
rect 3384 34892 3390 34944
rect 4157 34935 4215 34941
rect 4157 34901 4169 34935
rect 4203 34932 4215 34935
rect 4614 34932 4620 34944
rect 4203 34904 4620 34932
rect 4203 34901 4215 34904
rect 4157 34895 4215 34901
rect 4614 34892 4620 34904
rect 4672 34892 4678 34944
rect 8202 34892 8208 34944
rect 8260 34932 8266 34944
rect 9858 34932 9864 34944
rect 8260 34904 9864 34932
rect 8260 34892 8266 34904
rect 9858 34892 9864 34904
rect 9916 34892 9922 34944
rect 10244 34941 10272 34972
rect 11057 34969 11069 34972
rect 11103 34969 11115 35003
rect 11057 34963 11115 34969
rect 11238 34960 11244 35012
rect 11296 35000 11302 35012
rect 12084 35000 12112 35031
rect 13170 35028 13176 35080
rect 13228 35028 13234 35080
rect 13556 35077 13584 35244
rect 13909 35241 13921 35275
rect 13955 35272 13967 35275
rect 14366 35272 14372 35284
rect 13955 35244 14372 35272
rect 13955 35241 13967 35244
rect 13909 35235 13967 35241
rect 14366 35232 14372 35244
rect 14424 35232 14430 35284
rect 15378 35232 15384 35284
rect 15436 35272 15442 35284
rect 16209 35275 16267 35281
rect 16209 35272 16221 35275
rect 15436 35244 16221 35272
rect 15436 35232 15442 35244
rect 16209 35241 16221 35244
rect 16255 35241 16267 35275
rect 18322 35272 18328 35284
rect 16209 35235 16267 35241
rect 17420 35244 18328 35272
rect 15562 35164 15568 35216
rect 15620 35204 15626 35216
rect 16758 35204 16764 35216
rect 15620 35176 16764 35204
rect 15620 35164 15626 35176
rect 16758 35164 16764 35176
rect 16816 35164 16822 35216
rect 17034 35204 17040 35216
rect 16868 35176 17040 35204
rect 15746 35096 15752 35148
rect 15804 35136 15810 35148
rect 16868 35136 16896 35176
rect 17034 35164 17040 35176
rect 17092 35204 17098 35216
rect 17218 35204 17224 35216
rect 17092 35176 17224 35204
rect 17092 35164 17098 35176
rect 17218 35164 17224 35176
rect 17276 35204 17282 35216
rect 17420 35213 17448 35244
rect 18322 35232 18328 35244
rect 18380 35232 18386 35284
rect 19061 35275 19119 35281
rect 19061 35241 19073 35275
rect 19107 35272 19119 35275
rect 23201 35275 23259 35281
rect 19107 35244 21036 35272
rect 19107 35241 19119 35244
rect 19061 35235 19119 35241
rect 21008 35216 21036 35244
rect 23201 35241 23213 35275
rect 23247 35272 23259 35275
rect 24486 35272 24492 35284
rect 23247 35244 24492 35272
rect 23247 35241 23259 35244
rect 23201 35235 23259 35241
rect 24486 35232 24492 35244
rect 24544 35232 24550 35284
rect 24670 35232 24676 35284
rect 24728 35272 24734 35284
rect 24857 35275 24915 35281
rect 24857 35272 24869 35275
rect 24728 35244 24869 35272
rect 24728 35232 24734 35244
rect 24857 35241 24869 35244
rect 24903 35272 24915 35275
rect 25222 35272 25228 35284
rect 24903 35244 25228 35272
rect 24903 35241 24915 35244
rect 24857 35235 24915 35241
rect 25222 35232 25228 35244
rect 25280 35232 25286 35284
rect 26694 35272 26700 35284
rect 25700 35244 26700 35272
rect 17405 35207 17463 35213
rect 17405 35204 17417 35207
rect 17276 35176 17417 35204
rect 17276 35164 17282 35176
rect 17405 35173 17417 35176
rect 17451 35173 17463 35207
rect 18690 35204 18696 35216
rect 17405 35167 17463 35173
rect 17788 35176 18696 35204
rect 15804 35108 16896 35136
rect 15804 35096 15810 35108
rect 17126 35096 17132 35148
rect 17184 35096 17190 35148
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35037 13415 35071
rect 13357 35031 13415 35037
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35037 13599 35071
rect 13541 35031 13599 35037
rect 11296 34972 12112 35000
rect 11296 34960 11302 34972
rect 12250 34960 12256 35012
rect 12308 34960 12314 35012
rect 10229 34935 10287 34941
rect 10229 34901 10241 34935
rect 10275 34901 10287 34935
rect 10229 34895 10287 34901
rect 10962 34892 10968 34944
rect 11020 34892 11026 34944
rect 12802 34892 12808 34944
rect 12860 34932 12866 34944
rect 13173 34935 13231 34941
rect 13173 34932 13185 34935
rect 12860 34904 13185 34932
rect 12860 34892 12866 34904
rect 13173 34901 13185 34904
rect 13219 34901 13231 34935
rect 13372 34932 13400 35031
rect 13630 35028 13636 35080
rect 13688 35028 13694 35080
rect 13725 35071 13783 35077
rect 13725 35037 13737 35071
rect 13771 35068 13783 35071
rect 13906 35068 13912 35080
rect 13771 35040 13912 35068
rect 13771 35037 13783 35040
rect 13725 35031 13783 35037
rect 13906 35028 13912 35040
rect 13964 35028 13970 35080
rect 14093 35071 14151 35077
rect 14093 35037 14105 35071
rect 14139 35068 14151 35071
rect 14642 35068 14648 35080
rect 14139 35040 14648 35068
rect 14139 35037 14151 35040
rect 14093 35031 14151 35037
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 15565 35071 15623 35077
rect 15565 35068 15577 35071
rect 15488 35040 15577 35068
rect 14360 35003 14418 35009
rect 14360 34969 14372 35003
rect 14406 35000 14418 35003
rect 14918 35000 14924 35012
rect 14406 34972 14924 35000
rect 14406 34969 14418 34972
rect 14360 34963 14418 34969
rect 14918 34960 14924 34972
rect 14976 34960 14982 35012
rect 14090 34932 14096 34944
rect 13372 34904 14096 34932
rect 13173 34895 13231 34901
rect 14090 34892 14096 34904
rect 14148 34892 14154 34944
rect 14182 34892 14188 34944
rect 14240 34932 14246 34944
rect 15488 34941 15516 35040
rect 15565 35037 15577 35040
rect 15611 35037 15623 35071
rect 15565 35031 15623 35037
rect 16482 35028 16488 35080
rect 16540 35068 16546 35080
rect 17788 35077 17816 35176
rect 18690 35164 18696 35176
rect 18748 35204 18754 35216
rect 19426 35204 19432 35216
rect 18748 35176 19432 35204
rect 18748 35164 18754 35176
rect 19426 35164 19432 35176
rect 19484 35164 19490 35216
rect 20070 35164 20076 35216
rect 20128 35164 20134 35216
rect 20990 35164 20996 35216
rect 21048 35164 21054 35216
rect 23569 35207 23627 35213
rect 23569 35204 23581 35207
rect 22480 35176 23581 35204
rect 20088 35136 20116 35164
rect 22186 35136 22192 35148
rect 18524 35108 20116 35136
rect 21192 35108 22192 35136
rect 18524 35080 18552 35108
rect 17773 35071 17831 35077
rect 17773 35068 17785 35071
rect 16540 35040 17785 35068
rect 16540 35028 16546 35040
rect 17773 35037 17785 35040
rect 17819 35037 17831 35071
rect 17773 35031 17831 35037
rect 18506 35028 18512 35080
rect 18564 35028 18570 35080
rect 19245 35071 19303 35077
rect 19245 35037 19257 35071
rect 19291 35037 19303 35071
rect 19245 35031 19303 35037
rect 19260 35000 19288 35031
rect 20070 35028 20076 35080
rect 20128 35028 20134 35080
rect 20993 35071 21051 35077
rect 20993 35037 21005 35071
rect 21039 35037 21051 35071
rect 20993 35031 21051 35037
rect 16500 34972 19288 35000
rect 20625 35003 20683 35009
rect 16500 34941 16528 34972
rect 20625 34969 20637 35003
rect 20671 35000 20683 35003
rect 20898 35000 20904 35012
rect 20671 34972 20904 35000
rect 20671 34969 20683 34972
rect 20625 34963 20683 34969
rect 20898 34960 20904 34972
rect 20956 34960 20962 35012
rect 15473 34935 15531 34941
rect 15473 34932 15485 34935
rect 14240 34904 15485 34932
rect 14240 34892 14246 34904
rect 15473 34901 15485 34904
rect 15519 34901 15531 34935
rect 15473 34895 15531 34901
rect 16485 34935 16543 34941
rect 16485 34901 16497 34935
rect 16531 34901 16543 34935
rect 16485 34895 16543 34901
rect 16574 34892 16580 34944
rect 16632 34932 16638 34944
rect 16853 34935 16911 34941
rect 16853 34932 16865 34935
rect 16632 34904 16865 34932
rect 16632 34892 16638 34904
rect 16853 34901 16865 34904
rect 16899 34901 16911 34935
rect 16853 34895 16911 34901
rect 16945 34935 17003 34941
rect 16945 34901 16957 34935
rect 16991 34932 17003 34935
rect 17126 34932 17132 34944
rect 16991 34904 17132 34932
rect 16991 34901 17003 34904
rect 16945 34895 17003 34901
rect 17126 34892 17132 34904
rect 17184 34932 17190 34944
rect 18598 34932 18604 34944
rect 17184 34904 18604 34932
rect 17184 34892 17190 34904
rect 18598 34892 18604 34904
rect 18656 34892 18662 34944
rect 19058 34892 19064 34944
rect 19116 34932 19122 34944
rect 19889 34935 19947 34941
rect 19889 34932 19901 34935
rect 19116 34904 19901 34932
rect 19116 34892 19122 34904
rect 19889 34901 19901 34904
rect 19935 34901 19947 34935
rect 19889 34895 19947 34901
rect 20714 34892 20720 34944
rect 20772 34892 20778 34944
rect 21008 34932 21036 35031
rect 21082 35028 21088 35080
rect 21140 35028 21146 35080
rect 21192 35077 21220 35108
rect 22186 35096 22192 35108
rect 22244 35096 22250 35148
rect 21177 35071 21235 35077
rect 21177 35037 21189 35071
rect 21223 35037 21235 35071
rect 21177 35031 21235 35037
rect 21358 35028 21364 35080
rect 21416 35028 21422 35080
rect 22480 35077 22508 35176
rect 23569 35173 23581 35176
rect 23615 35204 23627 35207
rect 24394 35204 24400 35216
rect 23615 35176 24400 35204
rect 23615 35173 23627 35176
rect 23569 35167 23627 35173
rect 24394 35164 24400 35176
rect 24452 35164 24458 35216
rect 24581 35207 24639 35213
rect 24581 35173 24593 35207
rect 24627 35204 24639 35207
rect 25700 35204 25728 35244
rect 26694 35232 26700 35244
rect 26752 35232 26758 35284
rect 27614 35232 27620 35284
rect 27672 35272 27678 35284
rect 28626 35272 28632 35284
rect 27672 35244 28632 35272
rect 27672 35232 27678 35244
rect 28626 35232 28632 35244
rect 28684 35232 28690 35284
rect 30377 35275 30435 35281
rect 30377 35241 30389 35275
rect 30423 35272 30435 35275
rect 30926 35272 30932 35284
rect 30423 35244 30932 35272
rect 30423 35241 30435 35244
rect 30377 35235 30435 35241
rect 30926 35232 30932 35244
rect 30984 35232 30990 35284
rect 32214 35232 32220 35284
rect 32272 35232 32278 35284
rect 24627 35176 25728 35204
rect 24627 35173 24639 35176
rect 24581 35167 24639 35173
rect 23474 35096 23480 35148
rect 23532 35136 23538 35148
rect 24596 35136 24624 35167
rect 25866 35164 25872 35216
rect 25924 35204 25930 35216
rect 25961 35207 26019 35213
rect 25961 35204 25973 35207
rect 25924 35176 25973 35204
rect 25924 35164 25930 35176
rect 25961 35173 25973 35176
rect 26007 35173 26019 35207
rect 25961 35167 26019 35173
rect 27890 35164 27896 35216
rect 27948 35164 27954 35216
rect 28258 35164 28264 35216
rect 28316 35204 28322 35216
rect 30006 35204 30012 35216
rect 28316 35176 30012 35204
rect 28316 35164 28322 35176
rect 30006 35164 30012 35176
rect 30064 35164 30070 35216
rect 32493 35207 32551 35213
rect 32493 35204 32505 35207
rect 30668 35176 32505 35204
rect 23532 35108 24164 35136
rect 23532 35096 23538 35108
rect 24136 35077 24164 35108
rect 24320 35108 24624 35136
rect 22465 35071 22523 35077
rect 22465 35068 22477 35071
rect 22020 35040 22477 35068
rect 22020 35012 22048 35040
rect 22465 35037 22477 35040
rect 22511 35037 22523 35071
rect 22465 35031 22523 35037
rect 22741 35071 22799 35077
rect 22741 35037 22753 35071
rect 22787 35068 22799 35071
rect 23109 35071 23167 35077
rect 23109 35068 23121 35071
rect 22787 35040 23121 35068
rect 22787 35037 22799 35040
rect 22741 35031 22799 35037
rect 23109 35037 23121 35040
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 23293 35071 23351 35077
rect 23293 35037 23305 35071
rect 23339 35037 23351 35071
rect 23293 35031 23351 35037
rect 24121 35071 24179 35077
rect 24121 35037 24133 35071
rect 24167 35037 24179 35071
rect 24121 35031 24179 35037
rect 21818 34960 21824 35012
rect 21876 34960 21882 35012
rect 22002 34960 22008 35012
rect 22060 34960 22066 35012
rect 22189 35003 22247 35009
rect 22189 34969 22201 35003
rect 22235 35000 22247 35003
rect 22756 35000 22784 35031
rect 22235 34972 22784 35000
rect 22235 34969 22247 34972
rect 22189 34963 22247 34969
rect 21082 34932 21088 34944
rect 21008 34904 21088 34932
rect 21082 34892 21088 34904
rect 21140 34932 21146 34944
rect 22204 34932 22232 34963
rect 21140 34904 22232 34932
rect 21140 34892 21146 34904
rect 22278 34892 22284 34944
rect 22336 34892 22342 34944
rect 22646 34892 22652 34944
rect 22704 34892 22710 34944
rect 23124 34932 23152 35031
rect 23308 35000 23336 35031
rect 24320 35000 24348 35108
rect 24854 35096 24860 35148
rect 24912 35096 24918 35148
rect 24946 35096 24952 35148
rect 25004 35136 25010 35148
rect 28350 35136 28356 35148
rect 25004 35108 26648 35136
rect 25004 35096 25010 35108
rect 24397 35071 24455 35077
rect 24397 35037 24409 35071
rect 24443 35068 24455 35071
rect 24872 35068 24900 35096
rect 24443 35040 24900 35068
rect 24443 35037 24455 35040
rect 24397 35031 24455 35037
rect 25222 35028 25228 35080
rect 25280 35068 25286 35080
rect 25409 35071 25467 35077
rect 25409 35068 25421 35071
rect 25280 35040 25421 35068
rect 25280 35028 25286 35040
rect 25409 35037 25421 35040
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 25498 35028 25504 35080
rect 25556 35068 25562 35080
rect 25593 35071 25651 35077
rect 25593 35068 25605 35071
rect 25556 35040 25605 35068
rect 25556 35028 25562 35040
rect 25593 35037 25605 35040
rect 25639 35068 25651 35071
rect 25869 35071 25927 35077
rect 25869 35068 25881 35071
rect 25639 35040 25881 35068
rect 25639 35037 25651 35040
rect 25593 35031 25651 35037
rect 25869 35037 25881 35040
rect 25915 35037 25927 35071
rect 25869 35031 25927 35037
rect 25958 35028 25964 35080
rect 26016 35068 26022 35080
rect 26620 35077 26648 35108
rect 27080 35108 28356 35136
rect 26053 35071 26111 35077
rect 26053 35068 26065 35071
rect 26016 35040 26065 35068
rect 26016 35028 26022 35040
rect 26053 35037 26065 35040
rect 26099 35037 26111 35071
rect 26053 35031 26111 35037
rect 26605 35071 26663 35077
rect 26605 35037 26617 35071
rect 26651 35037 26663 35071
rect 26605 35031 26663 35037
rect 26878 35028 26884 35080
rect 26936 35068 26942 35080
rect 27080 35077 27108 35108
rect 28350 35096 28356 35108
rect 28408 35096 28414 35148
rect 28902 35096 28908 35148
rect 28960 35096 28966 35148
rect 28997 35139 29055 35145
rect 28997 35105 29009 35139
rect 29043 35105 29055 35139
rect 28997 35099 29055 35105
rect 29549 35139 29607 35145
rect 29549 35105 29561 35139
rect 29595 35136 29607 35139
rect 29822 35136 29828 35148
rect 29595 35108 29828 35136
rect 29595 35105 29607 35108
rect 29549 35099 29607 35105
rect 27065 35071 27123 35077
rect 27065 35068 27077 35071
rect 26936 35040 27077 35068
rect 26936 35028 26942 35040
rect 27065 35037 27077 35040
rect 27111 35037 27123 35071
rect 27065 35031 27123 35037
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35037 27951 35071
rect 27893 35031 27951 35037
rect 23308 34972 24348 35000
rect 25774 34960 25780 35012
rect 25832 34960 25838 35012
rect 26789 35003 26847 35009
rect 26789 34969 26801 35003
rect 26835 35000 26847 35003
rect 27709 35003 27767 35009
rect 27709 35000 27721 35003
rect 26835 34972 27721 35000
rect 26835 34969 26847 34972
rect 26789 34963 26847 34969
rect 27709 34969 27721 34972
rect 27755 34969 27767 35003
rect 27709 34963 27767 34969
rect 26050 34932 26056 34944
rect 23124 34904 26056 34932
rect 26050 34892 26056 34904
rect 26108 34892 26114 34944
rect 26694 34892 26700 34944
rect 26752 34932 26758 34944
rect 26973 34935 27031 34941
rect 26973 34932 26985 34935
rect 26752 34904 26985 34932
rect 26752 34892 26758 34904
rect 26973 34901 26985 34904
rect 27019 34901 27031 34935
rect 27908 34932 27936 35031
rect 28074 35028 28080 35080
rect 28132 35028 28138 35080
rect 28718 35028 28724 35080
rect 28776 35068 28782 35080
rect 29012 35068 29040 35099
rect 29822 35096 29828 35108
rect 29880 35096 29886 35148
rect 28776 35040 29040 35068
rect 29733 35071 29791 35077
rect 28776 35028 28782 35040
rect 29733 35037 29745 35071
rect 29779 35068 29791 35071
rect 29779 35040 30144 35068
rect 29779 35037 29791 35040
rect 29733 35031 29791 35037
rect 28442 34932 28448 34944
rect 27908 34904 28448 34932
rect 26973 34895 27031 34901
rect 28442 34892 28448 34904
rect 28500 34892 28506 34944
rect 28534 34892 28540 34944
rect 28592 34932 28598 34944
rect 28813 34935 28871 34941
rect 28813 34932 28825 34935
rect 28592 34904 28825 34932
rect 28592 34892 28598 34904
rect 28813 34901 28825 34904
rect 28859 34932 28871 34935
rect 29748 34932 29776 35031
rect 30006 34960 30012 35012
rect 30064 34960 30070 35012
rect 30116 35000 30144 35040
rect 30190 35028 30196 35080
rect 30248 35028 30254 35080
rect 30668 35012 30696 35176
rect 32493 35173 32505 35176
rect 32539 35173 32551 35207
rect 32493 35167 32551 35173
rect 32674 35164 32680 35216
rect 32732 35164 32738 35216
rect 31018 35096 31024 35148
rect 31076 35096 31082 35148
rect 31754 35096 31760 35148
rect 31812 35136 31818 35148
rect 31812 35108 32076 35136
rect 31812 35096 31818 35108
rect 30834 35028 30840 35080
rect 30892 35068 30898 35080
rect 32048 35077 32076 35108
rect 31113 35071 31171 35077
rect 31113 35068 31125 35071
rect 30892 35040 31125 35068
rect 30892 35028 30898 35040
rect 31113 35037 31125 35040
rect 31159 35037 31171 35071
rect 31113 35031 31171 35037
rect 31297 35071 31355 35077
rect 31297 35037 31309 35071
rect 31343 35068 31355 35071
rect 31941 35071 31999 35077
rect 31343 35040 31432 35068
rect 31343 35037 31355 35040
rect 31297 35031 31355 35037
rect 30650 35000 30656 35012
rect 30116 34972 30656 35000
rect 30650 34960 30656 34972
rect 30708 34960 30714 35012
rect 31404 34944 31432 35040
rect 31941 35037 31953 35071
rect 31987 35037 31999 35071
rect 31941 35031 31999 35037
rect 32033 35071 32091 35077
rect 32033 35037 32045 35071
rect 32079 35068 32091 35071
rect 32306 35068 32312 35080
rect 32079 35040 32312 35068
rect 32079 35037 32091 35040
rect 32033 35031 32091 35037
rect 31956 35000 31984 35031
rect 32306 35028 32312 35040
rect 32364 35068 32370 35080
rect 32692 35068 32720 35164
rect 32364 35040 32720 35068
rect 32364 35028 32370 35040
rect 32122 35000 32128 35012
rect 31956 34972 32128 35000
rect 32122 34960 32128 34972
rect 32180 34960 32186 35012
rect 28859 34904 29776 34932
rect 28859 34901 28871 34904
rect 28813 34895 28871 34901
rect 29914 34892 29920 34944
rect 29972 34892 29978 34944
rect 31386 34892 31392 34944
rect 31444 34932 31450 34944
rect 32861 34935 32919 34941
rect 32861 34932 32873 34935
rect 31444 34904 32873 34932
rect 31444 34892 31450 34904
rect 32861 34901 32873 34904
rect 32907 34901 32919 34935
rect 32861 34895 32919 34901
rect 1104 34842 43884 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 43884 34842
rect 1104 34768 43884 34790
rect 4157 34731 4215 34737
rect 4157 34697 4169 34731
rect 4203 34728 4215 34731
rect 4706 34728 4712 34740
rect 4203 34700 4712 34728
rect 4203 34697 4215 34700
rect 4157 34691 4215 34697
rect 4706 34688 4712 34700
rect 4764 34688 4770 34740
rect 7742 34688 7748 34740
rect 7800 34688 7806 34740
rect 8113 34731 8171 34737
rect 8113 34697 8125 34731
rect 8159 34728 8171 34731
rect 8159 34700 9812 34728
rect 8159 34697 8171 34700
rect 8113 34691 8171 34697
rect 9398 34660 9404 34672
rect 4264 34632 7052 34660
rect 4264 34601 4292 34632
rect 4249 34595 4307 34601
rect 4249 34561 4261 34595
rect 4295 34561 4307 34595
rect 4249 34555 4307 34561
rect 4516 34595 4574 34601
rect 4516 34561 4528 34595
rect 4562 34592 4574 34595
rect 4982 34592 4988 34604
rect 4562 34564 4988 34592
rect 4562 34561 4574 34564
rect 4516 34555 4574 34561
rect 4982 34552 4988 34564
rect 5040 34552 5046 34604
rect 6380 34601 6408 34632
rect 7024 34604 7052 34632
rect 8312 34632 9404 34660
rect 6365 34595 6423 34601
rect 6365 34561 6377 34595
rect 6411 34561 6423 34595
rect 6365 34555 6423 34561
rect 6632 34595 6690 34601
rect 6632 34561 6644 34595
rect 6678 34592 6690 34595
rect 6914 34592 6920 34604
rect 6678 34564 6920 34592
rect 6678 34561 6690 34564
rect 6632 34555 6690 34561
rect 6914 34552 6920 34564
rect 6972 34552 6978 34604
rect 7006 34552 7012 34604
rect 7064 34552 7070 34604
rect 1762 34484 1768 34536
rect 1820 34484 1826 34536
rect 2130 34484 2136 34536
rect 2188 34484 2194 34536
rect 2222 34484 2228 34536
rect 2280 34524 2286 34536
rect 2685 34527 2743 34533
rect 2685 34524 2697 34527
rect 2280 34496 2697 34524
rect 2280 34484 2286 34496
rect 2685 34493 2697 34496
rect 2731 34493 2743 34527
rect 2685 34487 2743 34493
rect 2866 34484 2872 34536
rect 2924 34484 2930 34536
rect 3510 34484 3516 34536
rect 3568 34484 3574 34536
rect 8312 34533 8340 34632
rect 9398 34620 9404 34632
rect 9456 34620 9462 34672
rect 9582 34620 9588 34672
rect 9640 34620 9646 34672
rect 8389 34595 8447 34601
rect 8389 34561 8401 34595
rect 8435 34592 8447 34595
rect 9493 34595 9551 34601
rect 9493 34592 9505 34595
rect 8435 34564 9505 34592
rect 8435 34561 8447 34564
rect 8389 34555 8447 34561
rect 9493 34561 9505 34564
rect 9539 34561 9551 34595
rect 9493 34555 9551 34561
rect 8297 34527 8355 34533
rect 8297 34493 8309 34527
rect 8343 34493 8355 34527
rect 8297 34487 8355 34493
rect 8662 34484 8668 34536
rect 8720 34524 8726 34536
rect 8849 34527 8907 34533
rect 8849 34524 8861 34527
rect 8720 34496 8861 34524
rect 8720 34484 8726 34496
rect 8849 34493 8861 34496
rect 8895 34493 8907 34527
rect 8849 34487 8907 34493
rect 9214 34484 9220 34536
rect 9272 34484 9278 34536
rect 9309 34527 9367 34533
rect 9309 34493 9321 34527
rect 9355 34524 9367 34527
rect 9582 34524 9588 34536
rect 9355 34496 9588 34524
rect 9355 34493 9367 34496
rect 9309 34487 9367 34493
rect 9582 34484 9588 34496
rect 9640 34484 9646 34536
rect 9784 34524 9812 34700
rect 9950 34688 9956 34740
rect 10008 34688 10014 34740
rect 10134 34688 10140 34740
rect 10192 34728 10198 34740
rect 11422 34728 11428 34740
rect 10192 34700 11428 34728
rect 10192 34688 10198 34700
rect 11422 34688 11428 34700
rect 11480 34688 11486 34740
rect 11793 34731 11851 34737
rect 11793 34697 11805 34731
rect 11839 34728 11851 34731
rect 11974 34728 11980 34740
rect 11839 34700 11980 34728
rect 11839 34697 11851 34700
rect 11793 34691 11851 34697
rect 11974 34688 11980 34700
rect 12032 34688 12038 34740
rect 12805 34731 12863 34737
rect 12805 34728 12817 34731
rect 12084 34700 12817 34728
rect 9968 34660 9996 34688
rect 9968 34632 10272 34660
rect 9858 34552 9864 34604
rect 9916 34552 9922 34604
rect 9950 34552 9956 34604
rect 10008 34552 10014 34604
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34592 10103 34595
rect 10134 34592 10140 34604
rect 10091 34564 10140 34592
rect 10091 34561 10103 34564
rect 10045 34555 10103 34561
rect 10134 34552 10140 34564
rect 10192 34552 10198 34604
rect 10244 34601 10272 34632
rect 12084 34601 12112 34700
rect 12805 34697 12817 34700
rect 12851 34728 12863 34731
rect 13078 34728 13084 34740
rect 12851 34700 13084 34728
rect 12851 34697 12863 34700
rect 12805 34691 12863 34697
rect 13078 34688 13084 34700
rect 13136 34688 13142 34740
rect 13173 34731 13231 34737
rect 13173 34697 13185 34731
rect 13219 34728 13231 34731
rect 13906 34728 13912 34740
rect 13219 34700 13912 34728
rect 13219 34697 13231 34700
rect 13173 34691 13231 34697
rect 13906 34688 13912 34700
rect 13964 34688 13970 34740
rect 14090 34688 14096 34740
rect 14148 34728 14154 34740
rect 14148 34700 14504 34728
rect 14148 34688 14154 34700
rect 14476 34672 14504 34700
rect 14918 34688 14924 34740
rect 14976 34688 14982 34740
rect 15102 34688 15108 34740
rect 15160 34688 15166 34740
rect 15289 34731 15347 34737
rect 15289 34697 15301 34731
rect 15335 34728 15347 34731
rect 15470 34728 15476 34740
rect 15335 34700 15476 34728
rect 15335 34697 15347 34700
rect 15289 34691 15347 34697
rect 15470 34688 15476 34700
rect 15528 34688 15534 34740
rect 16206 34688 16212 34740
rect 16264 34728 16270 34740
rect 16390 34728 16396 34740
rect 16264 34700 16396 34728
rect 16264 34688 16270 34700
rect 16390 34688 16396 34700
rect 16448 34728 16454 34740
rect 16448 34700 16804 34728
rect 16448 34688 16454 34700
rect 12989 34663 13047 34669
rect 12989 34660 13001 34663
rect 12636 34632 13001 34660
rect 10229 34595 10287 34601
rect 10229 34561 10241 34595
rect 10275 34561 10287 34595
rect 10229 34555 10287 34561
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34561 11943 34595
rect 11885 34555 11943 34561
rect 12069 34595 12127 34601
rect 12069 34561 12081 34595
rect 12115 34561 12127 34595
rect 12069 34555 12127 34561
rect 9968 34524 9996 34552
rect 9784 34496 9996 34524
rect 11790 34484 11796 34536
rect 11848 34484 11854 34536
rect 11900 34524 11928 34555
rect 12158 34552 12164 34604
rect 12216 34552 12222 34604
rect 12636 34601 12664 34632
rect 12989 34629 13001 34632
rect 13035 34629 13047 34663
rect 12989 34623 13047 34629
rect 13280 34632 14136 34660
rect 12253 34595 12311 34601
rect 12253 34561 12265 34595
rect 12299 34592 12311 34595
rect 12621 34595 12679 34601
rect 12621 34592 12633 34595
rect 12299 34564 12633 34592
rect 12299 34561 12311 34564
rect 12253 34555 12311 34561
rect 12621 34561 12633 34564
rect 12667 34561 12679 34595
rect 12621 34555 12679 34561
rect 12802 34552 12808 34604
rect 12860 34592 12866 34604
rect 13280 34601 13308 34632
rect 14108 34604 14136 34632
rect 14182 34620 14188 34672
rect 14240 34620 14246 34672
rect 14458 34620 14464 34672
rect 14516 34660 14522 34672
rect 15013 34663 15071 34669
rect 15013 34660 15025 34663
rect 14516 34632 15025 34660
rect 14516 34620 14522 34632
rect 15013 34629 15025 34632
rect 15059 34629 15071 34663
rect 15013 34623 15071 34629
rect 12897 34595 12955 34601
rect 12897 34592 12909 34595
rect 12860 34564 12909 34592
rect 12860 34552 12866 34564
rect 12897 34561 12909 34564
rect 12943 34561 12955 34595
rect 12897 34555 12955 34561
rect 13265 34595 13323 34601
rect 13265 34561 13277 34595
rect 13311 34561 13323 34595
rect 13265 34555 13323 34561
rect 13633 34595 13691 34601
rect 13633 34561 13645 34595
rect 13679 34561 13691 34595
rect 13633 34555 13691 34561
rect 12820 34524 12848 34552
rect 11900 34496 12848 34524
rect 13078 34484 13084 34536
rect 13136 34524 13142 34536
rect 13449 34527 13507 34533
rect 13449 34524 13461 34527
rect 13136 34496 13461 34524
rect 13136 34484 13142 34496
rect 13449 34493 13461 34496
rect 13495 34493 13507 34527
rect 13648 34524 13676 34555
rect 13814 34552 13820 34604
rect 13872 34552 13878 34604
rect 14090 34552 14096 34604
rect 14148 34552 14154 34604
rect 15120 34592 15148 34688
rect 16776 34672 16804 34700
rect 16942 34688 16948 34740
rect 17000 34728 17006 34740
rect 17494 34728 17500 34740
rect 17000 34700 17500 34728
rect 17000 34688 17006 34700
rect 17494 34688 17500 34700
rect 17552 34728 17558 34740
rect 18233 34731 18291 34737
rect 18233 34728 18245 34731
rect 17552 34700 18245 34728
rect 17552 34688 17558 34700
rect 18233 34697 18245 34700
rect 18279 34697 18291 34731
rect 18233 34691 18291 34697
rect 20070 34688 20076 34740
rect 20128 34688 20134 34740
rect 20714 34688 20720 34740
rect 20772 34688 20778 34740
rect 20898 34688 20904 34740
rect 20956 34688 20962 34740
rect 21637 34731 21695 34737
rect 21637 34697 21649 34731
rect 21683 34728 21695 34731
rect 21818 34728 21824 34740
rect 21683 34700 21824 34728
rect 21683 34697 21695 34700
rect 21637 34691 21695 34697
rect 21818 34688 21824 34700
rect 21876 34688 21882 34740
rect 22186 34688 22192 34740
rect 22244 34688 22250 34740
rect 22646 34688 22652 34740
rect 22704 34728 22710 34740
rect 22925 34731 22983 34737
rect 22925 34728 22937 34731
rect 22704 34700 22937 34728
rect 22704 34688 22710 34700
rect 22925 34697 22937 34700
rect 22971 34697 22983 34731
rect 22925 34691 22983 34697
rect 23014 34688 23020 34740
rect 23072 34728 23078 34740
rect 25869 34731 25927 34737
rect 25869 34728 25881 34731
rect 23072 34700 25881 34728
rect 23072 34688 23078 34700
rect 25869 34697 25881 34700
rect 25915 34697 25927 34731
rect 25869 34691 25927 34697
rect 26694 34688 26700 34740
rect 26752 34688 26758 34740
rect 27706 34728 27712 34740
rect 26896 34700 27712 34728
rect 16666 34660 16672 34672
rect 16224 34632 16672 34660
rect 15197 34595 15255 34601
rect 15197 34592 15209 34595
rect 14200 34564 14964 34592
rect 15120 34564 15209 34592
rect 14200 34524 14228 34564
rect 13648 34496 14228 34524
rect 13449 34487 13507 34493
rect 14274 34484 14280 34536
rect 14332 34484 14338 34536
rect 14550 34484 14556 34536
rect 14608 34484 14614 34536
rect 14936 34524 14964 34564
rect 15197 34561 15209 34564
rect 15243 34592 15255 34595
rect 15838 34592 15844 34604
rect 15243 34564 15844 34592
rect 15243 34561 15255 34564
rect 15197 34555 15255 34561
rect 15838 34552 15844 34564
rect 15896 34552 15902 34604
rect 16224 34601 16252 34632
rect 16666 34620 16672 34632
rect 16724 34620 16730 34672
rect 16758 34620 16764 34672
rect 16816 34620 16822 34672
rect 19426 34660 19432 34672
rect 16868 34632 19432 34660
rect 16209 34595 16267 34601
rect 16209 34561 16221 34595
rect 16255 34561 16267 34595
rect 16209 34555 16267 34561
rect 16482 34552 16488 34604
rect 16540 34552 16546 34604
rect 16868 34601 16896 34632
rect 19426 34620 19432 34632
rect 19484 34660 19490 34672
rect 19484 34632 20024 34660
rect 19484 34620 19490 34632
rect 16853 34595 16911 34601
rect 16853 34561 16865 34595
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17120 34595 17178 34601
rect 17120 34561 17132 34595
rect 17166 34592 17178 34595
rect 19058 34592 19064 34604
rect 17166 34564 19064 34592
rect 17166 34561 17178 34564
rect 17120 34555 17178 34561
rect 19058 34552 19064 34564
rect 19116 34552 19122 34604
rect 19245 34595 19303 34601
rect 19245 34561 19257 34595
rect 19291 34561 19303 34595
rect 19245 34555 19303 34561
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34592 19671 34595
rect 19886 34592 19892 34604
rect 19659 34564 19892 34592
rect 19659 34561 19671 34564
rect 19613 34555 19671 34561
rect 15286 34524 15292 34536
rect 14936 34496 15292 34524
rect 15286 34484 15292 34496
rect 15344 34484 15350 34536
rect 16025 34527 16083 34533
rect 16025 34493 16037 34527
rect 16071 34524 16083 34527
rect 16574 34524 16580 34536
rect 16071 34496 16580 34524
rect 16071 34493 16083 34496
rect 16025 34487 16083 34493
rect 16574 34484 16580 34496
rect 16632 34484 16638 34536
rect 18601 34527 18659 34533
rect 18601 34493 18613 34527
rect 18647 34524 18659 34527
rect 18690 34524 18696 34536
rect 18647 34496 18696 34524
rect 18647 34493 18659 34496
rect 18601 34487 18659 34493
rect 18690 34484 18696 34496
rect 18748 34484 18754 34536
rect 19150 34484 19156 34536
rect 19208 34484 19214 34536
rect 19260 34524 19288 34555
rect 19886 34552 19892 34564
rect 19944 34552 19950 34604
rect 19996 34601 20024 34632
rect 19981 34595 20039 34601
rect 19981 34561 19993 34595
rect 20027 34561 20039 34595
rect 20088 34592 20116 34688
rect 20248 34663 20306 34669
rect 20248 34629 20260 34663
rect 20294 34660 20306 34663
rect 20732 34660 20760 34688
rect 20294 34632 20760 34660
rect 20916 34660 20944 34688
rect 22005 34663 22063 34669
rect 22005 34660 22017 34663
rect 20916 34632 22017 34660
rect 20294 34629 20306 34632
rect 20248 34623 20306 34629
rect 22005 34629 22017 34632
rect 22051 34629 22063 34663
rect 23750 34660 23756 34672
rect 22005 34623 22063 34629
rect 22204 34632 23756 34660
rect 20622 34592 20628 34604
rect 20088 34564 20628 34592
rect 19981 34555 20039 34561
rect 20622 34552 20628 34564
rect 20680 34592 20686 34604
rect 20680 34564 21036 34592
rect 20680 34552 20686 34564
rect 19260 34496 19656 34524
rect 6178 34456 6184 34468
rect 5368 34428 6184 34456
rect 5368 34400 5396 34428
rect 6178 34416 6184 34428
rect 6236 34416 6242 34468
rect 8757 34459 8815 34465
rect 8757 34425 8769 34459
rect 8803 34456 8815 34459
rect 10318 34456 10324 34468
rect 8803 34428 10324 34456
rect 8803 34425 8815 34428
rect 8757 34419 8815 34425
rect 10318 34416 10324 34428
rect 10376 34416 10382 34468
rect 11808 34456 11836 34484
rect 11977 34459 12035 34465
rect 11977 34456 11989 34459
rect 11808 34428 11989 34456
rect 11977 34425 11989 34428
rect 12023 34425 12035 34459
rect 12802 34456 12808 34468
rect 11977 34419 12035 34425
rect 12360 34428 12808 34456
rect 3418 34348 3424 34400
rect 3476 34348 3482 34400
rect 5350 34348 5356 34400
rect 5408 34348 5414 34400
rect 5629 34391 5687 34397
rect 5629 34357 5641 34391
rect 5675 34388 5687 34391
rect 5994 34388 6000 34400
rect 5675 34360 6000 34388
rect 5675 34357 5687 34360
rect 5629 34351 5687 34357
rect 5994 34348 6000 34360
rect 6052 34348 6058 34400
rect 6546 34348 6552 34400
rect 6604 34388 6610 34400
rect 7098 34388 7104 34400
rect 6604 34360 7104 34388
rect 6604 34348 6610 34360
rect 7098 34348 7104 34360
rect 7156 34348 7162 34400
rect 10505 34391 10563 34397
rect 10505 34357 10517 34391
rect 10551 34388 10563 34391
rect 10870 34388 10876 34400
rect 10551 34360 10876 34388
rect 10551 34357 10563 34360
rect 10505 34351 10563 34357
rect 10870 34348 10876 34360
rect 10928 34348 10934 34400
rect 10962 34348 10968 34400
rect 11020 34388 11026 34400
rect 11333 34391 11391 34397
rect 11333 34388 11345 34391
rect 11020 34360 11345 34388
rect 11020 34348 11026 34360
rect 11333 34357 11345 34360
rect 11379 34388 11391 34391
rect 12360 34388 12388 34428
rect 12802 34416 12808 34428
rect 12860 34456 12866 34468
rect 13357 34459 13415 34465
rect 12860 34428 13124 34456
rect 12860 34416 12866 34428
rect 11379 34360 12388 34388
rect 11379 34357 11391 34360
rect 11333 34351 11391 34357
rect 12434 34348 12440 34400
rect 12492 34348 12498 34400
rect 12986 34348 12992 34400
rect 13044 34348 13050 34400
rect 13096 34388 13124 34428
rect 13357 34425 13369 34459
rect 13403 34456 13415 34459
rect 14568 34456 14596 34484
rect 13403 34428 14596 34456
rect 13403 34425 13415 34428
rect 13357 34419 13415 34425
rect 15102 34416 15108 34468
rect 15160 34456 15166 34468
rect 15470 34456 15476 34468
rect 15160 34428 15476 34456
rect 15160 34416 15166 34428
rect 15470 34416 15476 34428
rect 15528 34416 15534 34468
rect 15933 34391 15991 34397
rect 15933 34388 15945 34391
rect 13096 34360 15945 34388
rect 15933 34357 15945 34360
rect 15979 34388 15991 34391
rect 17034 34388 17040 34400
rect 15979 34360 17040 34388
rect 15979 34357 15991 34360
rect 15933 34351 15991 34357
rect 17034 34348 17040 34360
rect 17092 34348 17098 34400
rect 19628 34388 19656 34496
rect 19702 34484 19708 34536
rect 19760 34484 19766 34536
rect 21008 34524 21036 34564
rect 21266 34552 21272 34604
rect 21324 34592 21330 34604
rect 21453 34595 21511 34601
rect 21453 34592 21465 34595
rect 21324 34564 21465 34592
rect 21324 34552 21330 34564
rect 21453 34561 21465 34564
rect 21499 34561 21511 34595
rect 21453 34555 21511 34561
rect 21637 34595 21695 34601
rect 21637 34561 21649 34595
rect 21683 34561 21695 34595
rect 21637 34555 21695 34561
rect 21008 34496 21404 34524
rect 21376 34465 21404 34496
rect 21361 34459 21419 34465
rect 21361 34425 21373 34459
rect 21407 34425 21419 34459
rect 21361 34419 21419 34425
rect 20714 34388 20720 34400
rect 19628 34360 20720 34388
rect 20714 34348 20720 34360
rect 20772 34348 20778 34400
rect 20990 34348 20996 34400
rect 21048 34388 21054 34400
rect 21266 34388 21272 34400
rect 21048 34360 21272 34388
rect 21048 34348 21054 34360
rect 21266 34348 21272 34360
rect 21324 34388 21330 34400
rect 21652 34388 21680 34555
rect 21818 34552 21824 34604
rect 21876 34592 21882 34604
rect 22204 34592 22232 34632
rect 21876 34564 22232 34592
rect 21876 34552 21882 34564
rect 22278 34552 22284 34604
rect 22336 34592 22342 34604
rect 23477 34595 23535 34601
rect 23477 34592 23489 34595
rect 22336 34564 23489 34592
rect 22336 34552 22342 34564
rect 23477 34561 23489 34564
rect 23523 34561 23535 34595
rect 23477 34555 23535 34561
rect 22370 34484 22376 34536
rect 22428 34484 22434 34536
rect 23201 34527 23259 34533
rect 23201 34493 23213 34527
rect 23247 34493 23259 34527
rect 23201 34487 23259 34493
rect 23216 34456 23244 34487
rect 23290 34484 23296 34536
rect 23348 34484 23354 34536
rect 23385 34527 23443 34533
rect 23385 34493 23397 34527
rect 23431 34524 23443 34527
rect 23584 34524 23612 34632
rect 23750 34620 23756 34632
rect 23808 34660 23814 34672
rect 24670 34660 24676 34672
rect 23808 34632 24676 34660
rect 23808 34620 23814 34632
rect 24670 34620 24676 34632
rect 24728 34620 24734 34672
rect 24762 34620 24768 34672
rect 24820 34620 24826 34672
rect 24995 34629 25053 34635
rect 24486 34552 24492 34604
rect 24544 34592 24550 34604
rect 24995 34595 25007 34629
rect 25041 34595 25053 34629
rect 25332 34632 25535 34660
rect 25332 34601 25360 34632
rect 24995 34592 25053 34595
rect 24544 34589 25053 34592
rect 25317 34595 25375 34601
rect 24544 34564 25024 34589
rect 24544 34552 24550 34564
rect 25317 34561 25329 34595
rect 25363 34561 25375 34595
rect 25317 34555 25375 34561
rect 25406 34552 25412 34604
rect 25464 34552 25470 34604
rect 25507 34592 25535 34632
rect 25682 34620 25688 34672
rect 25740 34660 25746 34672
rect 26418 34660 26424 34672
rect 25740 34632 26424 34660
rect 25740 34620 25746 34632
rect 26418 34620 26424 34632
rect 26476 34620 26482 34672
rect 25866 34592 25872 34604
rect 25507 34564 25872 34592
rect 25866 34552 25872 34564
rect 25924 34552 25930 34604
rect 26050 34552 26056 34604
rect 26108 34592 26114 34604
rect 26329 34595 26387 34601
rect 26329 34592 26341 34595
rect 26108 34564 26341 34592
rect 26108 34552 26114 34564
rect 26329 34561 26341 34564
rect 26375 34561 26387 34595
rect 26329 34555 26387 34561
rect 26605 34595 26663 34601
rect 26605 34561 26617 34595
rect 26651 34592 26663 34595
rect 26712 34592 26740 34688
rect 26651 34564 26740 34592
rect 26789 34595 26847 34601
rect 26651 34561 26663 34564
rect 26605 34555 26663 34561
rect 26789 34561 26801 34595
rect 26835 34592 26847 34595
rect 26896 34592 26924 34700
rect 27706 34688 27712 34700
rect 27764 34688 27770 34740
rect 28166 34688 28172 34740
rect 28224 34688 28230 34740
rect 28350 34688 28356 34740
rect 28408 34688 28414 34740
rect 28442 34688 28448 34740
rect 28500 34688 28506 34740
rect 29273 34731 29331 34737
rect 29273 34697 29285 34731
rect 29319 34728 29331 34731
rect 29546 34728 29552 34740
rect 29319 34700 29552 34728
rect 29319 34697 29331 34700
rect 29273 34691 29331 34697
rect 29546 34688 29552 34700
rect 29604 34688 29610 34740
rect 29914 34688 29920 34740
rect 29972 34688 29978 34740
rect 30282 34688 30288 34740
rect 30340 34728 30346 34740
rect 31757 34731 31815 34737
rect 31757 34728 31769 34731
rect 30340 34700 31769 34728
rect 30340 34688 30346 34700
rect 31757 34697 31769 34700
rect 31803 34697 31815 34731
rect 31757 34691 31815 34697
rect 32306 34688 32312 34740
rect 32364 34688 32370 34740
rect 27240 34663 27298 34669
rect 27240 34629 27252 34663
rect 27286 34660 27298 34663
rect 28184 34660 28212 34688
rect 27286 34632 28212 34660
rect 27286 34629 27298 34632
rect 27240 34623 27298 34629
rect 26835 34564 26924 34592
rect 26835 34561 26847 34564
rect 26789 34555 26847 34561
rect 26896 34536 26924 34564
rect 26970 34552 26976 34604
rect 27028 34552 27034 34604
rect 27522 34552 27528 34604
rect 27580 34592 27586 34604
rect 28460 34592 28488 34688
rect 29632 34663 29690 34669
rect 29632 34629 29644 34663
rect 29678 34660 29690 34663
rect 29932 34660 29960 34688
rect 29678 34632 29960 34660
rect 29678 34629 29690 34632
rect 29632 34623 29690 34629
rect 28629 34595 28687 34601
rect 28629 34592 28641 34595
rect 27580 34564 28028 34592
rect 28460 34564 28641 34592
rect 27580 34552 27586 34564
rect 23431 34496 23612 34524
rect 23937 34527 23995 34533
rect 23431 34493 23443 34496
rect 23385 34487 23443 34493
rect 23937 34493 23949 34527
rect 23983 34524 23995 34527
rect 24854 34524 24860 34536
rect 23983 34496 24860 34524
rect 23983 34493 23995 34496
rect 23937 34487 23995 34493
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 25038 34484 25044 34536
rect 25096 34524 25102 34536
rect 26142 34524 26148 34536
rect 25096 34496 26148 34524
rect 25096 34484 25102 34496
rect 26142 34484 26148 34496
rect 26200 34484 26206 34536
rect 26878 34484 26884 34536
rect 26936 34484 26942 34536
rect 24394 34456 24400 34468
rect 23216 34428 24400 34456
rect 24394 34416 24400 34428
rect 24452 34416 24458 34468
rect 25501 34459 25559 34465
rect 25501 34456 25513 34459
rect 24964 34428 25513 34456
rect 21324 34360 21680 34388
rect 21324 34348 21330 34360
rect 23014 34348 23020 34400
rect 23072 34348 23078 34400
rect 23842 34348 23848 34400
rect 23900 34388 23906 34400
rect 24964 34397 24992 34428
rect 25501 34425 25513 34428
rect 25547 34425 25559 34459
rect 25501 34419 25559 34425
rect 24489 34391 24547 34397
rect 24489 34388 24501 34391
rect 23900 34360 24501 34388
rect 23900 34348 23906 34360
rect 24489 34357 24501 34360
rect 24535 34357 24547 34391
rect 24489 34351 24547 34357
rect 24949 34391 25007 34397
rect 24949 34357 24961 34391
rect 24995 34357 25007 34391
rect 24949 34351 25007 34357
rect 25130 34348 25136 34400
rect 25188 34348 25194 34400
rect 25516 34388 25544 34419
rect 26418 34416 26424 34468
rect 26476 34416 26482 34468
rect 26510 34416 26516 34468
rect 26568 34416 26574 34468
rect 28000 34456 28028 34564
rect 28629 34561 28641 34564
rect 28675 34561 28687 34595
rect 30837 34595 30895 34601
rect 30837 34592 30849 34595
rect 28629 34555 28687 34561
rect 30760 34564 30849 34592
rect 28074 34484 28080 34536
rect 28132 34524 28138 34536
rect 28445 34527 28503 34533
rect 28445 34524 28457 34527
rect 28132 34496 28457 34524
rect 28132 34484 28138 34496
rect 28445 34493 28457 34496
rect 28491 34524 28503 34527
rect 28902 34524 28908 34536
rect 28491 34496 28908 34524
rect 28491 34493 28503 34496
rect 28445 34487 28503 34493
rect 28902 34484 28908 34496
rect 28960 34484 28966 34536
rect 29362 34484 29368 34536
rect 29420 34484 29426 34536
rect 30760 34465 30788 34564
rect 30837 34561 30849 34564
rect 30883 34561 30895 34595
rect 30837 34555 30895 34561
rect 28813 34459 28871 34465
rect 28813 34456 28825 34459
rect 28000 34428 28825 34456
rect 28813 34425 28825 34428
rect 28859 34425 28871 34459
rect 28813 34419 28871 34425
rect 30745 34459 30803 34465
rect 30745 34425 30757 34459
rect 30791 34425 30803 34459
rect 30745 34419 30803 34425
rect 25590 34388 25596 34400
rect 25516 34360 25596 34388
rect 25590 34348 25596 34360
rect 25648 34348 25654 34400
rect 26145 34391 26203 34397
rect 26145 34357 26157 34391
rect 26191 34388 26203 34391
rect 27154 34388 27160 34400
rect 26191 34360 27160 34388
rect 26191 34357 26203 34360
rect 26145 34351 26203 34357
rect 27154 34348 27160 34360
rect 27212 34348 27218 34400
rect 27338 34348 27344 34400
rect 27396 34388 27402 34400
rect 28534 34388 28540 34400
rect 27396 34360 28540 34388
rect 27396 34348 27402 34360
rect 28534 34348 28540 34360
rect 28592 34348 28598 34400
rect 30558 34348 30564 34400
rect 30616 34388 30622 34400
rect 31481 34391 31539 34397
rect 31481 34388 31493 34391
rect 30616 34360 31493 34388
rect 30616 34348 30622 34360
rect 31481 34357 31493 34360
rect 31527 34357 31539 34391
rect 31481 34351 31539 34357
rect 1104 34298 43884 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 43884 34298
rect 1104 34224 43884 34246
rect 2130 34144 2136 34196
rect 2188 34184 2194 34196
rect 2685 34187 2743 34193
rect 2685 34184 2697 34187
rect 2188 34156 2697 34184
rect 2188 34144 2194 34156
rect 2685 34153 2697 34156
rect 2731 34153 2743 34187
rect 2685 34147 2743 34153
rect 4249 34187 4307 34193
rect 4249 34153 4261 34187
rect 4295 34184 4307 34187
rect 4614 34184 4620 34196
rect 4295 34156 4620 34184
rect 4295 34153 4307 34156
rect 4249 34147 4307 34153
rect 4614 34144 4620 34156
rect 4672 34184 4678 34196
rect 6822 34184 6828 34196
rect 4672 34156 6828 34184
rect 4672 34144 4678 34156
rect 6822 34144 6828 34156
rect 6880 34144 6886 34196
rect 7558 34144 7564 34196
rect 7616 34184 7622 34196
rect 8389 34187 8447 34193
rect 8389 34184 8401 34187
rect 7616 34156 8401 34184
rect 7616 34144 7622 34156
rect 8389 34153 8401 34156
rect 8435 34153 8447 34187
rect 8389 34147 8447 34153
rect 8570 34144 8576 34196
rect 8628 34184 8634 34196
rect 8665 34187 8723 34193
rect 8665 34184 8677 34187
rect 8628 34156 8677 34184
rect 8628 34144 8634 34156
rect 8665 34153 8677 34156
rect 8711 34184 8723 34187
rect 9122 34184 9128 34196
rect 8711 34156 9128 34184
rect 8711 34153 8723 34156
rect 8665 34147 8723 34153
rect 9122 34144 9128 34156
rect 9180 34144 9186 34196
rect 9306 34144 9312 34196
rect 9364 34184 9370 34196
rect 9401 34187 9459 34193
rect 9401 34184 9413 34187
rect 9364 34156 9413 34184
rect 9364 34144 9370 34156
rect 9401 34153 9413 34156
rect 9447 34153 9459 34187
rect 9401 34147 9459 34153
rect 9585 34187 9643 34193
rect 9585 34153 9597 34187
rect 9631 34184 9643 34187
rect 9766 34184 9772 34196
rect 9631 34156 9772 34184
rect 9631 34153 9643 34156
rect 9585 34147 9643 34153
rect 9766 34144 9772 34156
rect 9824 34144 9830 34196
rect 9950 34144 9956 34196
rect 10008 34184 10014 34196
rect 10137 34187 10195 34193
rect 10137 34184 10149 34187
rect 10008 34156 10149 34184
rect 10008 34144 10014 34156
rect 10137 34153 10149 34156
rect 10183 34184 10195 34187
rect 10962 34184 10968 34196
rect 10183 34156 10968 34184
rect 10183 34153 10195 34156
rect 10137 34147 10195 34153
rect 10962 34144 10968 34156
rect 11020 34144 11026 34196
rect 11149 34187 11207 34193
rect 11149 34153 11161 34187
rect 11195 34184 11207 34187
rect 11238 34184 11244 34196
rect 11195 34156 11244 34184
rect 11195 34153 11207 34156
rect 11149 34147 11207 34153
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 11793 34187 11851 34193
rect 11793 34153 11805 34187
rect 11839 34184 11851 34187
rect 12250 34184 12256 34196
rect 11839 34156 12256 34184
rect 11839 34153 11851 34156
rect 11793 34147 11851 34153
rect 12250 34144 12256 34156
rect 12308 34144 12314 34196
rect 13538 34144 13544 34196
rect 13596 34144 13602 34196
rect 15194 34144 15200 34196
rect 15252 34144 15258 34196
rect 17402 34184 17408 34196
rect 15304 34156 17408 34184
rect 4982 34076 4988 34128
rect 5040 34076 5046 34128
rect 5077 34119 5135 34125
rect 5077 34085 5089 34119
rect 5123 34085 5135 34119
rect 5077 34079 5135 34085
rect 1946 34008 1952 34060
rect 2004 34048 2010 34060
rect 3326 34048 3332 34060
rect 2004 34020 3332 34048
rect 2004 34008 2010 34020
rect 3326 34008 3332 34020
rect 3384 34048 3390 34060
rect 4062 34048 4068 34060
rect 3384 34020 4068 34048
rect 3384 34008 3390 34020
rect 4062 34008 4068 34020
rect 4120 34008 4126 34060
rect 4433 34051 4491 34057
rect 4433 34017 4445 34051
rect 4479 34048 4491 34051
rect 5092 34048 5120 34079
rect 5534 34076 5540 34128
rect 5592 34116 5598 34128
rect 5592 34088 5672 34116
rect 5592 34076 5598 34088
rect 5644 34057 5672 34088
rect 4479 34020 5120 34048
rect 5629 34051 5687 34057
rect 4479 34017 4491 34020
rect 4433 34011 4491 34017
rect 5629 34017 5641 34051
rect 5675 34017 5687 34051
rect 5629 34011 5687 34017
rect 6270 34008 6276 34060
rect 6328 34008 6334 34060
rect 6454 34008 6460 34060
rect 6512 34008 6518 34060
rect 6638 34008 6644 34060
rect 6696 34008 6702 34060
rect 934 33940 940 33992
rect 992 33980 998 33992
rect 1581 33983 1639 33989
rect 1581 33980 1593 33983
rect 992 33952 1593 33980
rect 992 33940 998 33952
rect 1581 33949 1593 33952
rect 1627 33949 1639 33983
rect 1581 33943 1639 33949
rect 2038 33940 2044 33992
rect 2096 33940 2102 33992
rect 5537 33983 5595 33989
rect 5537 33949 5549 33983
rect 5583 33980 5595 33983
rect 6288 33980 6316 34008
rect 6840 33989 6868 34144
rect 9217 34119 9275 34125
rect 9217 34116 9229 34119
rect 8036 34088 9229 34116
rect 5583 33952 6316 33980
rect 6825 33983 6883 33989
rect 5583 33949 5595 33952
rect 5537 33943 5595 33949
rect 6825 33949 6837 33983
rect 6871 33949 6883 33983
rect 7190 33980 7196 33992
rect 6825 33943 6883 33949
rect 6932 33952 7196 33980
rect 3053 33915 3111 33921
rect 3053 33881 3065 33915
rect 3099 33912 3111 33915
rect 3418 33912 3424 33924
rect 3099 33884 3424 33912
rect 3099 33881 3111 33884
rect 3053 33875 3111 33881
rect 3418 33872 3424 33884
rect 3476 33912 3482 33924
rect 6365 33915 6423 33921
rect 3476 33884 3924 33912
rect 3476 33872 3482 33884
rect 3896 33856 3924 33884
rect 6365 33881 6377 33915
rect 6411 33912 6423 33915
rect 6932 33912 6960 33952
rect 7190 33940 7196 33952
rect 7248 33940 7254 33992
rect 7466 33940 7472 33992
rect 7524 33980 7530 33992
rect 8036 33989 8064 34088
rect 9217 34085 9229 34088
rect 9263 34085 9275 34119
rect 9217 34079 9275 34085
rect 12618 34076 12624 34128
rect 12676 34116 12682 34128
rect 13556 34116 13584 34144
rect 12676 34088 13584 34116
rect 13633 34119 13691 34125
rect 12676 34076 12682 34088
rect 8113 34051 8171 34057
rect 8113 34017 8125 34051
rect 8159 34017 8171 34051
rect 8113 34011 8171 34017
rect 8021 33983 8079 33989
rect 8021 33980 8033 33983
rect 7524 33952 8033 33980
rect 7524 33940 7530 33952
rect 8021 33949 8033 33952
rect 8067 33949 8079 33983
rect 8128 33980 8156 34011
rect 8662 34008 8668 34060
rect 8720 34048 8726 34060
rect 8720 34020 9720 34048
rect 8720 34008 8726 34020
rect 8754 33980 8760 33992
rect 8128 33952 8760 33980
rect 8021 33943 8079 33949
rect 8754 33940 8760 33952
rect 8812 33980 8818 33992
rect 9692 33989 9720 34020
rect 10870 34008 10876 34060
rect 10928 34048 10934 34060
rect 11241 34051 11299 34057
rect 11241 34048 11253 34051
rect 10928 34020 11253 34048
rect 10928 34008 10934 34020
rect 11241 34017 11253 34020
rect 11287 34048 11299 34051
rect 11287 34020 11658 34048
rect 11287 34017 11299 34020
rect 11241 34011 11299 34017
rect 8941 33983 8999 33989
rect 8941 33980 8953 33983
rect 8812 33952 8953 33980
rect 8812 33940 8818 33952
rect 8941 33949 8953 33952
rect 8987 33949 8999 33983
rect 8941 33943 8999 33949
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33980 9551 33983
rect 9677 33983 9735 33989
rect 9539 33952 9628 33980
rect 9539 33949 9551 33952
rect 9493 33943 9551 33949
rect 9600 33924 9628 33952
rect 9677 33949 9689 33983
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33949 11023 33983
rect 10965 33943 11023 33949
rect 6411 33884 6960 33912
rect 6411 33881 6423 33884
rect 6365 33875 6423 33881
rect 7006 33872 7012 33924
rect 7064 33912 7070 33924
rect 7561 33915 7619 33921
rect 7561 33912 7573 33915
rect 7064 33884 7573 33912
rect 7064 33872 7070 33884
rect 7561 33881 7573 33884
rect 7607 33881 7619 33915
rect 7561 33875 7619 33881
rect 9582 33872 9588 33924
rect 9640 33872 9646 33924
rect 10502 33872 10508 33924
rect 10560 33872 10566 33924
rect 2590 33804 2596 33856
rect 2648 33804 2654 33856
rect 3145 33847 3203 33853
rect 3145 33813 3157 33847
rect 3191 33844 3203 33847
rect 3602 33844 3608 33856
rect 3191 33816 3608 33844
rect 3191 33813 3203 33816
rect 3145 33807 3203 33813
rect 3602 33804 3608 33816
rect 3660 33804 3666 33856
rect 3878 33804 3884 33856
rect 3936 33804 3942 33856
rect 5442 33804 5448 33856
rect 5500 33804 5506 33856
rect 5997 33847 6055 33853
rect 5997 33813 6009 33847
rect 6043 33844 6055 33847
rect 7282 33844 7288 33856
rect 6043 33816 7288 33844
rect 6043 33813 6055 33816
rect 5997 33807 6055 33813
rect 7282 33804 7288 33816
rect 7340 33804 7346 33856
rect 10980 33844 11008 33943
rect 11054 33940 11060 33992
rect 11112 33940 11118 33992
rect 11238 33844 11244 33856
rect 10980 33816 11244 33844
rect 11238 33804 11244 33816
rect 11296 33804 11302 33856
rect 11630 33844 11658 34020
rect 11698 34008 11704 34060
rect 11756 34008 11762 34060
rect 11992 34020 12664 34048
rect 11992 33989 12020 34020
rect 11977 33983 12035 33989
rect 11977 33949 11989 33983
rect 12023 33949 12035 33983
rect 11977 33943 12035 33949
rect 12066 33940 12072 33992
rect 12124 33940 12130 33992
rect 12158 33940 12164 33992
rect 12216 33940 12222 33992
rect 12253 33983 12311 33989
rect 12253 33949 12265 33983
rect 12299 33949 12311 33983
rect 12253 33943 12311 33949
rect 12268 33912 12296 33943
rect 12434 33940 12440 33992
rect 12492 33940 12498 33992
rect 12636 33989 12664 34020
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33980 12679 33983
rect 12802 33980 12808 33992
rect 12667 33952 12808 33980
rect 12667 33949 12679 33952
rect 12621 33943 12679 33949
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 12912 33989 12940 34088
rect 13633 34085 13645 34119
rect 13679 34116 13691 34119
rect 15102 34116 15108 34128
rect 13679 34088 15108 34116
rect 13679 34085 13691 34088
rect 13633 34079 13691 34085
rect 15102 34076 15108 34088
rect 15160 34076 15166 34128
rect 13262 34008 13268 34060
rect 13320 34008 13326 34060
rect 13906 34008 13912 34060
rect 13964 34048 13970 34060
rect 14826 34048 14832 34060
rect 13964 34020 14832 34048
rect 13964 34008 13970 34020
rect 12897 33983 12955 33989
rect 12897 33949 12909 33983
rect 12943 33949 12955 33983
rect 12897 33943 12955 33949
rect 13078 33940 13084 33992
rect 13136 33940 13142 33992
rect 13173 33983 13231 33989
rect 13173 33949 13185 33983
rect 13219 33949 13231 33983
rect 13173 33943 13231 33949
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33980 13507 33983
rect 13538 33980 13544 33992
rect 13495 33952 13544 33980
rect 13495 33949 13507 33952
rect 13449 33943 13507 33949
rect 12529 33915 12587 33921
rect 12529 33912 12541 33915
rect 12268 33884 12541 33912
rect 12529 33881 12541 33884
rect 12575 33881 12587 33915
rect 12529 33875 12587 33881
rect 12710 33872 12716 33924
rect 12768 33912 12774 33924
rect 13188 33912 13216 33943
rect 12768 33884 13216 33912
rect 12768 33872 12774 33884
rect 13464 33844 13492 33943
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 14090 33940 14096 33992
rect 14148 33940 14154 33992
rect 14292 33989 14320 34020
rect 14826 34008 14832 34020
rect 14884 34008 14890 34060
rect 15212 34048 15240 34144
rect 15304 34057 15332 34156
rect 17402 34144 17408 34156
rect 17460 34144 17466 34196
rect 19610 34144 19616 34196
rect 19668 34184 19674 34196
rect 22370 34184 22376 34196
rect 19668 34156 22376 34184
rect 19668 34144 19674 34156
rect 22370 34144 22376 34156
rect 22428 34144 22434 34196
rect 23198 34144 23204 34196
rect 23256 34184 23262 34196
rect 24578 34184 24584 34196
rect 23256 34156 24584 34184
rect 23256 34144 23262 34156
rect 24578 34144 24584 34156
rect 24636 34144 24642 34196
rect 24859 34144 24865 34196
rect 24917 34184 24923 34196
rect 25133 34187 25191 34193
rect 25133 34184 25145 34187
rect 24917 34156 25145 34184
rect 24917 34144 24923 34156
rect 25133 34153 25145 34156
rect 25179 34153 25191 34187
rect 25133 34147 25191 34153
rect 26418 34144 26424 34196
rect 26476 34144 26482 34196
rect 26510 34144 26516 34196
rect 26568 34184 26574 34196
rect 26697 34187 26755 34193
rect 26697 34184 26709 34187
rect 26568 34156 26709 34184
rect 26568 34144 26574 34156
rect 26697 34153 26709 34156
rect 26743 34153 26755 34187
rect 26697 34147 26755 34153
rect 27062 34144 27068 34196
rect 27120 34184 27126 34196
rect 29178 34184 29184 34196
rect 27120 34156 29184 34184
rect 27120 34144 27126 34156
rect 29178 34144 29184 34156
rect 29236 34184 29242 34196
rect 29273 34187 29331 34193
rect 29273 34184 29285 34187
rect 29236 34156 29285 34184
rect 29236 34144 29242 34156
rect 29273 34153 29285 34156
rect 29319 34153 29331 34187
rect 29273 34147 29331 34153
rect 31386 34144 31392 34196
rect 31444 34144 31450 34196
rect 16022 34116 16028 34128
rect 15488 34088 16028 34116
rect 14936 34020 15240 34048
rect 15289 34051 15347 34057
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33949 14335 33983
rect 14277 33943 14335 33949
rect 14550 33940 14556 33992
rect 14608 33940 14614 33992
rect 14936 33989 14964 34020
rect 15289 34017 15301 34051
rect 15335 34017 15347 34051
rect 15289 34011 15347 34017
rect 14921 33983 14979 33989
rect 14921 33949 14933 33983
rect 14967 33949 14979 33983
rect 14921 33943 14979 33949
rect 15010 33940 15016 33992
rect 15068 33940 15074 33992
rect 15102 33940 15108 33992
rect 15160 33980 15166 33992
rect 15304 33980 15332 34011
rect 15160 33952 15332 33980
rect 15160 33940 15166 33952
rect 15378 33940 15384 33992
rect 15436 33980 15442 33992
rect 15488 33989 15516 34088
rect 16022 34076 16028 34088
rect 16080 34076 16086 34128
rect 17126 34076 17132 34128
rect 17184 34076 17190 34128
rect 18616 34088 20024 34116
rect 18616 34060 18644 34088
rect 15838 34008 15844 34060
rect 15896 34008 15902 34060
rect 15948 34020 18092 34048
rect 15948 33992 15976 34020
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 15436 33952 15485 33980
rect 15436 33940 15442 33952
rect 15473 33949 15485 33952
rect 15519 33949 15531 33983
rect 15473 33943 15531 33949
rect 15930 33940 15936 33992
rect 15988 33940 15994 33992
rect 17405 33983 17463 33989
rect 17405 33980 17417 33983
rect 16316 33952 17417 33980
rect 14108 33912 14136 33940
rect 14734 33912 14740 33924
rect 14108 33884 14740 33912
rect 14734 33872 14740 33884
rect 14792 33872 14798 33924
rect 15028 33912 15056 33940
rect 16316 33912 16344 33952
rect 17405 33949 17417 33952
rect 17451 33949 17463 33983
rect 17405 33943 17463 33949
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33949 17555 33983
rect 17497 33943 17555 33949
rect 15028 33884 16344 33912
rect 16390 33872 16396 33924
rect 16448 33912 16454 33924
rect 16669 33915 16727 33921
rect 16669 33912 16681 33915
rect 16448 33884 16681 33912
rect 16448 33872 16454 33884
rect 16669 33881 16681 33884
rect 16715 33881 16727 33915
rect 16669 33875 16727 33881
rect 17034 33872 17040 33924
rect 17092 33912 17098 33924
rect 17512 33912 17540 33943
rect 17586 33940 17592 33992
rect 17644 33940 17650 33992
rect 17770 33940 17776 33992
rect 17828 33940 17834 33992
rect 17092 33884 17540 33912
rect 17865 33915 17923 33921
rect 17092 33872 17098 33884
rect 17420 33856 17448 33884
rect 17865 33881 17877 33915
rect 17911 33912 17923 33915
rect 17954 33912 17960 33924
rect 17911 33884 17960 33912
rect 17911 33881 17923 33884
rect 17865 33875 17923 33881
rect 17954 33872 17960 33884
rect 18012 33872 18018 33924
rect 18064 33912 18092 34020
rect 18598 34008 18604 34060
rect 18656 34008 18662 34060
rect 18892 34020 19656 34048
rect 19996 34034 20024 34088
rect 20346 34076 20352 34128
rect 20404 34116 20410 34128
rect 20625 34119 20683 34125
rect 20625 34116 20637 34119
rect 20404 34088 20637 34116
rect 20404 34076 20410 34088
rect 20625 34085 20637 34088
rect 20671 34085 20683 34119
rect 20625 34079 20683 34085
rect 22646 34076 22652 34128
rect 22704 34076 22710 34128
rect 25038 34076 25044 34128
rect 25096 34076 25102 34128
rect 26234 34076 26240 34128
rect 26292 34076 26298 34128
rect 26436 34116 26464 34144
rect 27614 34116 27620 34128
rect 26436 34088 27620 34116
rect 27614 34076 27620 34088
rect 27672 34076 27678 34128
rect 27706 34076 27712 34128
rect 27764 34076 27770 34128
rect 20809 34051 20867 34057
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 18782 33980 18788 33992
rect 18555 33952 18788 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 18782 33940 18788 33952
rect 18840 33940 18846 33992
rect 18892 33989 18920 34020
rect 19628 33992 19656 34020
rect 20809 34017 20821 34051
rect 20855 34048 20867 34051
rect 22186 34048 22192 34060
rect 20855 34020 22192 34048
rect 20855 34017 20867 34020
rect 20809 34011 20867 34017
rect 22186 34008 22192 34020
rect 22244 34008 22250 34060
rect 22664 34048 22692 34076
rect 24673 34051 24731 34057
rect 22664 34020 22876 34048
rect 18877 33983 18935 33989
rect 18877 33949 18889 33983
rect 18923 33949 18935 33983
rect 18877 33943 18935 33949
rect 18966 33940 18972 33992
rect 19024 33980 19030 33992
rect 19245 33983 19303 33989
rect 19245 33980 19257 33983
rect 19024 33952 19257 33980
rect 19024 33940 19030 33952
rect 19245 33949 19257 33952
rect 19291 33949 19303 33983
rect 19245 33943 19303 33949
rect 19610 33940 19616 33992
rect 19668 33940 19674 33992
rect 19886 33940 19892 33992
rect 19944 33980 19950 33992
rect 20257 33983 20315 33989
rect 20257 33980 20269 33983
rect 19944 33952 20269 33980
rect 19944 33940 19950 33952
rect 20257 33949 20269 33952
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 20346 33940 20352 33992
rect 20404 33980 20410 33992
rect 21358 33980 21364 33992
rect 20404 33952 21364 33980
rect 20404 33940 20410 33952
rect 21358 33940 21364 33952
rect 21416 33940 21422 33992
rect 21453 33983 21511 33989
rect 21453 33949 21465 33983
rect 21499 33980 21511 33983
rect 21634 33980 21640 33992
rect 21499 33952 21640 33980
rect 21499 33949 21511 33952
rect 21453 33943 21511 33949
rect 21468 33912 21496 33943
rect 21634 33940 21640 33952
rect 21692 33980 21698 33992
rect 22649 33983 22707 33989
rect 22649 33980 22661 33983
rect 21692 33952 22661 33980
rect 21692 33940 21698 33952
rect 22649 33949 22661 33952
rect 22695 33980 22707 33983
rect 22738 33980 22744 33992
rect 22695 33952 22744 33980
rect 22695 33949 22707 33952
rect 22649 33943 22707 33949
rect 22738 33940 22744 33952
rect 22796 33940 22802 33992
rect 22848 33989 22876 34020
rect 24673 34017 24685 34051
rect 24719 34048 24731 34051
rect 25056 34048 25084 34076
rect 24719 34020 25084 34048
rect 26252 34048 26280 34076
rect 26510 34048 26516 34060
rect 26252 34020 26516 34048
rect 24719 34017 24731 34020
rect 24673 34011 24731 34017
rect 26510 34008 26516 34020
rect 26568 34048 26574 34060
rect 27724 34048 27752 34076
rect 26568 34020 27016 34048
rect 26568 34008 26574 34020
rect 22833 33983 22891 33989
rect 22833 33949 22845 33983
rect 22879 33949 22891 33983
rect 22833 33943 22891 33949
rect 23100 33983 23158 33989
rect 23100 33949 23112 33983
rect 23146 33980 23158 33983
rect 23842 33980 23848 33992
rect 23146 33952 23848 33980
rect 23146 33949 23158 33952
rect 23100 33943 23158 33949
rect 23842 33940 23848 33952
rect 23900 33940 23906 33992
rect 24397 33983 24455 33989
rect 24397 33980 24409 33983
rect 24320 33952 24409 33980
rect 24320 33924 24348 33952
rect 24397 33949 24409 33952
rect 24443 33949 24455 33983
rect 24397 33943 24455 33949
rect 24569 33983 24627 33989
rect 24569 33949 24581 33983
rect 24615 33949 24627 33983
rect 24569 33943 24627 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 24949 33983 25007 33989
rect 24949 33949 24961 33983
rect 24995 33982 25007 33983
rect 25317 33983 25375 33989
rect 24995 33954 25176 33982
rect 24995 33949 25007 33954
rect 24949 33943 25007 33949
rect 18064 33884 21496 33912
rect 21910 33872 21916 33924
rect 21968 33912 21974 33924
rect 22189 33915 22247 33921
rect 22189 33912 22201 33915
rect 21968 33884 22201 33912
rect 21968 33872 21974 33884
rect 22189 33881 22201 33884
rect 22235 33881 22247 33915
rect 22189 33875 22247 33881
rect 11630 33816 13492 33844
rect 13814 33804 13820 33856
rect 13872 33844 13878 33856
rect 14185 33847 14243 33853
rect 14185 33844 14197 33847
rect 13872 33816 14197 33844
rect 13872 33804 13878 33816
rect 14185 33813 14197 33816
rect 14231 33813 14243 33847
rect 14185 33807 14243 33813
rect 17402 33804 17408 33856
rect 17460 33804 17466 33856
rect 18782 33804 18788 33856
rect 18840 33844 18846 33856
rect 19702 33844 19708 33856
rect 18840 33816 19708 33844
rect 18840 33804 18846 33816
rect 19702 33804 19708 33816
rect 19760 33804 19766 33856
rect 21358 33804 21364 33856
rect 21416 33804 21422 33856
rect 22204 33844 22232 33875
rect 22922 33872 22928 33924
rect 22980 33912 22986 33924
rect 24026 33912 24032 33924
rect 22980 33884 24032 33912
rect 22980 33872 22986 33884
rect 24026 33872 24032 33884
rect 24084 33912 24090 33924
rect 24084 33884 24256 33912
rect 24084 33872 24090 33884
rect 22646 33844 22652 33856
rect 22204 33816 22652 33844
rect 22646 33804 22652 33816
rect 22704 33804 22710 33856
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 23382 33844 23388 33856
rect 22796 33816 23388 33844
rect 22796 33804 22802 33816
rect 23382 33804 23388 33816
rect 23440 33804 23446 33856
rect 24228 33853 24256 33884
rect 24302 33872 24308 33924
rect 24360 33872 24366 33924
rect 24213 33847 24271 33853
rect 24213 33813 24225 33847
rect 24259 33813 24271 33847
rect 24596 33844 24624 33943
rect 24780 33912 24808 33943
rect 24780 33884 24992 33912
rect 24964 33856 24992 33884
rect 24670 33844 24676 33856
rect 24596 33816 24676 33844
rect 24213 33807 24271 33813
rect 24670 33804 24676 33816
rect 24728 33804 24734 33856
rect 24946 33804 24952 33856
rect 25004 33804 25010 33856
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 25148 33844 25176 33954
rect 25317 33949 25329 33983
rect 25363 33980 25375 33983
rect 25498 33980 25504 33992
rect 25363 33952 25504 33980
rect 25363 33949 25375 33952
rect 25317 33943 25375 33949
rect 25498 33940 25504 33952
rect 25556 33940 25562 33992
rect 25866 33940 25872 33992
rect 25924 33940 25930 33992
rect 26142 33940 26148 33992
rect 26200 33940 26206 33992
rect 26237 33983 26295 33989
rect 26237 33949 26249 33983
rect 26283 33980 26295 33983
rect 26605 33983 26663 33989
rect 26283 33952 26464 33980
rect 26283 33949 26295 33952
rect 26237 33943 26295 33949
rect 25682 33872 25688 33924
rect 25740 33912 25746 33924
rect 25884 33912 25912 33940
rect 25740 33884 26372 33912
rect 25740 33872 25746 33884
rect 26068 33856 26096 33884
rect 25869 33847 25927 33853
rect 25869 33844 25881 33847
rect 25096 33816 25881 33844
rect 25096 33804 25102 33816
rect 25869 33813 25881 33816
rect 25915 33813 25927 33847
rect 25869 33807 25927 33813
rect 25958 33804 25964 33856
rect 26016 33804 26022 33856
rect 26050 33804 26056 33856
rect 26108 33804 26114 33856
rect 26344 33853 26372 33884
rect 26329 33847 26387 33853
rect 26329 33813 26341 33847
rect 26375 33813 26387 33847
rect 26436 33844 26464 33952
rect 26605 33949 26617 33983
rect 26651 33980 26663 33983
rect 26694 33980 26700 33992
rect 26651 33952 26700 33980
rect 26651 33949 26663 33952
rect 26605 33943 26663 33949
rect 26694 33940 26700 33952
rect 26752 33940 26758 33992
rect 26988 33989 27016 34020
rect 27264 34020 27752 34048
rect 26973 33983 27031 33989
rect 26973 33949 26985 33983
rect 27019 33949 27031 33983
rect 26973 33943 27031 33949
rect 27062 33940 27068 33992
rect 27120 33940 27126 33992
rect 27154 33940 27160 33992
rect 27212 33940 27218 33992
rect 26513 33915 26571 33921
rect 26513 33881 26525 33915
rect 26559 33912 26571 33915
rect 27264 33912 27292 34020
rect 27982 34008 27988 34060
rect 28040 34008 28046 34060
rect 28350 34008 28356 34060
rect 28408 34048 28414 34060
rect 28810 34048 28816 34060
rect 28408 34020 28816 34048
rect 28408 34008 28414 34020
rect 28810 34008 28816 34020
rect 28868 34048 28874 34060
rect 29917 34051 29975 34057
rect 28868 34020 29132 34048
rect 28868 34008 28874 34020
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33980 27399 33983
rect 27522 33980 27528 33992
rect 27387 33952 27528 33980
rect 27387 33949 27399 33952
rect 27341 33943 27399 33949
rect 27522 33940 27528 33952
rect 27580 33980 27586 33992
rect 27580 33952 27660 33980
rect 27580 33940 27586 33952
rect 26559 33884 27292 33912
rect 26559 33881 26571 33884
rect 26513 33875 26571 33881
rect 27430 33872 27436 33924
rect 27488 33872 27494 33924
rect 27632 33912 27660 33952
rect 27890 33940 27896 33992
rect 27948 33940 27954 33992
rect 28074 33940 28080 33992
rect 28132 33940 28138 33992
rect 28258 33940 28264 33992
rect 28316 33980 28322 33992
rect 28445 33983 28503 33989
rect 28445 33980 28457 33983
rect 28316 33952 28457 33980
rect 28316 33940 28322 33952
rect 28445 33949 28457 33952
rect 28491 33949 28503 33983
rect 28445 33943 28503 33949
rect 28721 33983 28779 33989
rect 28721 33949 28733 33983
rect 28767 33980 28779 33983
rect 28902 33980 28908 33992
rect 28767 33952 28908 33980
rect 28767 33949 28779 33952
rect 28721 33943 28779 33949
rect 28902 33940 28908 33952
rect 28960 33940 28966 33992
rect 29104 33989 29132 34020
rect 29917 34017 29929 34051
rect 29963 34048 29975 34051
rect 30558 34048 30564 34060
rect 29963 34020 30564 34048
rect 29963 34017 29975 34020
rect 29917 34011 29975 34017
rect 30558 34008 30564 34020
rect 30616 34008 30622 34060
rect 30650 34008 30656 34060
rect 30708 34048 30714 34060
rect 30929 34051 30987 34057
rect 30929 34048 30941 34051
rect 30708 34020 30941 34048
rect 30708 34008 30714 34020
rect 30929 34017 30941 34020
rect 30975 34017 30987 34051
rect 30929 34011 30987 34017
rect 29089 33983 29147 33989
rect 29089 33949 29101 33983
rect 29135 33949 29147 33983
rect 29089 33943 29147 33949
rect 29454 33940 29460 33992
rect 29512 33980 29518 33992
rect 30009 33983 30067 33989
rect 30009 33980 30021 33983
rect 29512 33952 30021 33980
rect 29512 33940 29518 33952
rect 30009 33949 30021 33952
rect 30055 33949 30067 33983
rect 30009 33943 30067 33949
rect 30193 33983 30251 33989
rect 30193 33949 30205 33983
rect 30239 33980 30251 33983
rect 31404 33980 31432 34144
rect 30239 33952 31432 33980
rect 30239 33949 30251 33952
rect 30193 33943 30251 33949
rect 27908 33912 27936 33940
rect 27632 33884 27936 33912
rect 27154 33844 27160 33856
rect 26436 33816 27160 33844
rect 26329 33807 26387 33813
rect 27154 33804 27160 33816
rect 27212 33844 27218 33856
rect 27448 33844 27476 33872
rect 27212 33816 27476 33844
rect 27212 33804 27218 33816
rect 27614 33804 27620 33856
rect 27672 33804 27678 33856
rect 27706 33804 27712 33856
rect 27764 33804 27770 33856
rect 27801 33847 27859 33853
rect 27801 33813 27813 33847
rect 27847 33844 27859 33847
rect 28074 33844 28080 33856
rect 27847 33816 28080 33844
rect 27847 33813 27859 33816
rect 27801 33807 27859 33813
rect 28074 33804 28080 33816
rect 28132 33804 28138 33856
rect 1104 33754 43884 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 43884 33754
rect 1104 33680 43884 33702
rect 1946 33600 1952 33652
rect 2004 33600 2010 33652
rect 2038 33600 2044 33652
rect 2096 33600 2102 33652
rect 2590 33600 2596 33652
rect 2648 33600 2654 33652
rect 3421 33643 3479 33649
rect 3421 33609 3433 33643
rect 3467 33640 3479 33643
rect 3510 33640 3516 33652
rect 3467 33612 3516 33640
rect 3467 33609 3479 33612
rect 3421 33603 3479 33609
rect 3510 33600 3516 33612
rect 3568 33600 3574 33652
rect 5442 33600 5448 33652
rect 5500 33640 5506 33652
rect 7009 33643 7067 33649
rect 7009 33640 7021 33643
rect 5500 33612 7021 33640
rect 5500 33600 5506 33612
rect 7009 33609 7021 33612
rect 7055 33609 7067 33643
rect 7009 33603 7067 33609
rect 8662 33600 8668 33652
rect 8720 33600 8726 33652
rect 8754 33600 8760 33652
rect 8812 33600 8818 33652
rect 9582 33600 9588 33652
rect 9640 33640 9646 33652
rect 9861 33643 9919 33649
rect 9861 33640 9873 33643
rect 9640 33612 9873 33640
rect 9640 33600 9646 33612
rect 9861 33609 9873 33612
rect 9907 33609 9919 33643
rect 9861 33603 9919 33609
rect 10597 33643 10655 33649
rect 10597 33609 10609 33643
rect 10643 33640 10655 33643
rect 11054 33640 11060 33652
rect 10643 33612 11060 33640
rect 10643 33609 10655 33612
rect 10597 33603 10655 33609
rect 11054 33600 11060 33612
rect 11112 33600 11118 33652
rect 11514 33640 11520 33652
rect 11256 33612 11520 33640
rect 2056 33504 2084 33600
rect 2308 33575 2366 33581
rect 2308 33541 2320 33575
rect 2354 33572 2366 33575
rect 2608 33572 2636 33600
rect 9493 33575 9551 33581
rect 9493 33572 9505 33575
rect 2354 33544 2636 33572
rect 8496 33544 9505 33572
rect 2354 33541 2366 33544
rect 2308 33535 2366 33541
rect 3881 33507 3939 33513
rect 2056 33476 3556 33504
rect 1854 33396 1860 33448
rect 1912 33436 1918 33448
rect 2041 33439 2099 33445
rect 2041 33436 2053 33439
rect 1912 33408 2053 33436
rect 1912 33396 1918 33408
rect 2041 33405 2053 33408
rect 2087 33405 2099 33439
rect 2041 33399 2099 33405
rect 3528 33377 3556 33476
rect 3881 33473 3893 33507
rect 3927 33504 3939 33507
rect 4706 33504 4712 33516
rect 3927 33476 4712 33504
rect 3927 33473 3939 33476
rect 3881 33467 3939 33473
rect 4706 33464 4712 33476
rect 4764 33504 4770 33516
rect 5813 33507 5871 33513
rect 5813 33504 5825 33507
rect 4764 33476 5825 33504
rect 4764 33464 4770 33476
rect 5813 33473 5825 33476
rect 5859 33473 5871 33507
rect 5813 33467 5871 33473
rect 5994 33464 6000 33516
rect 6052 33504 6058 33516
rect 6365 33507 6423 33513
rect 6365 33504 6377 33507
rect 6052 33476 6377 33504
rect 6052 33464 6058 33476
rect 6365 33473 6377 33476
rect 6411 33473 6423 33507
rect 6365 33467 6423 33473
rect 6638 33464 6644 33516
rect 6696 33504 6702 33516
rect 8496 33513 8524 33544
rect 9140 33516 9168 33544
rect 9493 33541 9505 33544
rect 9539 33541 9551 33575
rect 9493 33535 9551 33541
rect 10965 33575 11023 33581
rect 10965 33541 10977 33575
rect 11011 33572 11023 33575
rect 11256 33572 11284 33612
rect 11514 33600 11520 33612
rect 11572 33600 11578 33652
rect 11615 33643 11673 33649
rect 11615 33609 11627 33643
rect 11661 33640 11673 33643
rect 12158 33640 12164 33652
rect 11661 33612 12164 33640
rect 11661 33609 11673 33612
rect 11615 33603 11673 33609
rect 12158 33600 12164 33612
rect 12216 33600 12222 33652
rect 12437 33643 12495 33649
rect 12437 33609 12449 33643
rect 12483 33640 12495 33643
rect 12526 33640 12532 33652
rect 12483 33612 12532 33640
rect 12483 33609 12495 33612
rect 12437 33603 12495 33609
rect 12526 33600 12532 33612
rect 12584 33600 12590 33652
rect 13078 33600 13084 33652
rect 13136 33600 13142 33652
rect 13170 33600 13176 33652
rect 13228 33640 13234 33652
rect 13228 33612 13492 33640
rect 13228 33600 13234 33612
rect 11011 33544 11284 33572
rect 11885 33575 11943 33581
rect 11011 33541 11023 33544
rect 10965 33535 11023 33541
rect 11885 33541 11897 33575
rect 11931 33572 11943 33575
rect 12805 33575 12863 33581
rect 12805 33572 12817 33575
rect 11931 33544 12817 33572
rect 11931 33541 11943 33544
rect 11885 33535 11943 33541
rect 12805 33541 12817 33544
rect 12851 33572 12863 33575
rect 12851 33544 13216 33572
rect 12851 33541 12863 33544
rect 12805 33535 12863 33541
rect 8481 33507 8539 33513
rect 6696 33476 7512 33504
rect 6696 33464 6702 33476
rect 3970 33396 3976 33448
rect 4028 33396 4034 33448
rect 4062 33396 4068 33448
rect 4120 33396 4126 33448
rect 4890 33396 4896 33448
rect 4948 33396 4954 33448
rect 5721 33439 5779 33445
rect 5721 33405 5733 33439
rect 5767 33405 5779 33439
rect 5721 33399 5779 33405
rect 3513 33371 3571 33377
rect 3513 33337 3525 33371
rect 3559 33337 3571 33371
rect 3513 33331 3571 33337
rect 3878 33328 3884 33380
rect 3936 33368 3942 33380
rect 5736 33368 5764 33399
rect 7374 33396 7380 33448
rect 7432 33396 7438 33448
rect 7484 33436 7512 33476
rect 8481 33473 8493 33507
rect 8527 33473 8539 33507
rect 8481 33467 8539 33473
rect 8665 33507 8723 33513
rect 8665 33473 8677 33507
rect 8711 33473 8723 33507
rect 8665 33467 8723 33473
rect 8941 33507 8999 33513
rect 8941 33473 8953 33507
rect 8987 33504 8999 33507
rect 9122 33504 9128 33516
rect 8987 33476 9128 33504
rect 8987 33473 8999 33476
rect 8941 33467 8999 33473
rect 8680 33436 8708 33467
rect 9122 33464 9128 33476
rect 9180 33464 9186 33516
rect 9214 33464 9220 33516
rect 9272 33464 9278 33516
rect 9306 33464 9312 33516
rect 9364 33504 9370 33516
rect 9401 33507 9459 33513
rect 9401 33504 9413 33507
rect 9364 33476 9413 33504
rect 9364 33464 9370 33476
rect 9401 33473 9413 33476
rect 9447 33473 9459 33507
rect 9401 33467 9459 33473
rect 9677 33507 9735 33513
rect 9677 33473 9689 33507
rect 9723 33473 9735 33507
rect 9677 33467 9735 33473
rect 9692 33436 9720 33467
rect 10594 33464 10600 33516
rect 10652 33464 10658 33516
rect 10686 33464 10692 33516
rect 10744 33504 10750 33516
rect 10980 33504 11008 33535
rect 10744 33476 11008 33504
rect 11149 33507 11207 33513
rect 10744 33464 10750 33476
rect 11149 33473 11161 33507
rect 11195 33473 11207 33507
rect 11149 33467 11207 33473
rect 7484 33408 9720 33436
rect 10873 33439 10931 33445
rect 10873 33405 10885 33439
rect 10919 33436 10931 33439
rect 11054 33436 11060 33448
rect 10919 33408 11060 33436
rect 10919 33405 10931 33408
rect 10873 33399 10931 33405
rect 11054 33396 11060 33408
rect 11112 33396 11118 33448
rect 11164 33436 11192 33467
rect 11238 33464 11244 33516
rect 11296 33504 11302 33516
rect 11517 33507 11575 33513
rect 11517 33504 11529 33507
rect 11296 33476 11529 33504
rect 11296 33464 11302 33476
rect 11517 33473 11529 33476
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 11698 33464 11704 33516
rect 11756 33464 11762 33516
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 12069 33507 12127 33513
rect 12069 33473 12081 33507
rect 12115 33504 12127 33507
rect 12158 33504 12164 33516
rect 12115 33476 12164 33504
rect 12115 33473 12127 33476
rect 12069 33467 12127 33473
rect 11330 33436 11336 33448
rect 11164 33408 11336 33436
rect 3936 33340 5764 33368
rect 6181 33371 6239 33377
rect 3936 33328 3942 33340
rect 6181 33337 6193 33371
rect 6227 33368 6239 33371
rect 10962 33368 10968 33380
rect 6227 33340 10968 33368
rect 6227 33337 6239 33340
rect 6181 33331 6239 33337
rect 10962 33328 10968 33340
rect 11020 33328 11026 33380
rect 3418 33260 3424 33312
rect 3476 33300 3482 33312
rect 4525 33303 4583 33309
rect 4525 33300 4537 33303
rect 3476 33272 4537 33300
rect 3476 33260 3482 33272
rect 4525 33269 4537 33272
rect 4571 33300 4583 33303
rect 5350 33300 5356 33312
rect 4571 33272 5356 33300
rect 4571 33269 4583 33272
rect 4525 33263 4583 33269
rect 5350 33260 5356 33272
rect 5408 33260 5414 33312
rect 5537 33303 5595 33309
rect 5537 33269 5549 33303
rect 5583 33300 5595 33303
rect 5626 33300 5632 33312
rect 5583 33272 5632 33300
rect 5583 33269 5595 33272
rect 5537 33263 5595 33269
rect 5626 33260 5632 33272
rect 5684 33260 5690 33312
rect 7926 33260 7932 33312
rect 7984 33260 7990 33312
rect 8386 33260 8392 33312
rect 8444 33260 8450 33312
rect 10505 33303 10563 33309
rect 10505 33269 10517 33303
rect 10551 33300 10563 33303
rect 10870 33300 10876 33312
rect 10551 33272 10876 33300
rect 10551 33269 10563 33272
rect 10505 33263 10563 33269
rect 10870 33260 10876 33272
rect 10928 33300 10934 33312
rect 11164 33300 11192 33408
rect 11330 33396 11336 33408
rect 11388 33396 11394 33448
rect 11808 33368 11836 33467
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 12250 33464 12256 33516
rect 12308 33464 12314 33516
rect 12342 33464 12348 33516
rect 12400 33504 12406 33516
rect 12621 33507 12679 33513
rect 12400 33476 12572 33504
rect 12400 33464 12406 33476
rect 12544 33436 12572 33476
rect 12621 33473 12633 33507
rect 12667 33504 12679 33507
rect 12710 33504 12716 33516
rect 12667 33476 12716 33504
rect 12667 33473 12679 33476
rect 12621 33467 12679 33473
rect 12710 33464 12716 33476
rect 12768 33464 12774 33516
rect 12894 33464 12900 33516
rect 12952 33504 12958 33516
rect 13188 33513 13216 33544
rect 13464 33513 13492 33612
rect 13998 33600 14004 33652
rect 14056 33640 14062 33652
rect 15930 33640 15936 33652
rect 14056 33612 15936 33640
rect 14056 33600 14062 33612
rect 15930 33600 15936 33612
rect 15988 33600 15994 33652
rect 16206 33600 16212 33652
rect 16264 33600 16270 33652
rect 16298 33600 16304 33652
rect 16356 33600 16362 33652
rect 16758 33600 16764 33652
rect 16816 33640 16822 33652
rect 18046 33640 18052 33652
rect 16816 33612 18052 33640
rect 16816 33600 16822 33612
rect 18046 33600 18052 33612
rect 18104 33600 18110 33652
rect 18138 33600 18144 33652
rect 18196 33640 18202 33652
rect 18966 33640 18972 33652
rect 18196 33612 18972 33640
rect 18196 33600 18202 33612
rect 18966 33600 18972 33612
rect 19024 33640 19030 33652
rect 20806 33640 20812 33652
rect 19024 33612 20812 33640
rect 19024 33600 19030 33612
rect 20806 33600 20812 33612
rect 20864 33600 20870 33652
rect 21358 33640 21364 33652
rect 21284 33612 21364 33640
rect 14185 33575 14243 33581
rect 14185 33541 14197 33575
rect 14231 33572 14243 33575
rect 14458 33572 14464 33584
rect 14231 33544 14464 33572
rect 14231 33541 14243 33544
rect 14185 33535 14243 33541
rect 14458 33532 14464 33544
rect 14516 33532 14522 33584
rect 15102 33572 15108 33584
rect 14568 33544 15108 33572
rect 12989 33507 13047 33513
rect 12989 33504 13001 33507
rect 12952 33476 13001 33504
rect 12952 33464 12958 33476
rect 12989 33473 13001 33476
rect 13035 33473 13047 33507
rect 12989 33467 13047 33473
rect 13173 33507 13231 33513
rect 13173 33473 13185 33507
rect 13219 33473 13231 33507
rect 13173 33467 13231 33473
rect 13265 33507 13323 33513
rect 13265 33473 13277 33507
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 13449 33507 13507 33513
rect 13449 33473 13461 33507
rect 13495 33473 13507 33507
rect 13449 33467 13507 33473
rect 13280 33436 13308 33467
rect 13630 33464 13636 33516
rect 13688 33504 13694 33516
rect 14568 33513 14596 33544
rect 15102 33532 15108 33544
rect 15160 33532 15166 33584
rect 15286 33532 15292 33584
rect 15344 33572 15350 33584
rect 15344 33544 15976 33572
rect 15344 33532 15350 33544
rect 14093 33507 14151 33513
rect 14093 33504 14105 33507
rect 13688 33476 14105 33504
rect 13688 33464 13694 33476
rect 14093 33473 14105 33476
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 14277 33507 14335 33513
rect 14277 33473 14289 33507
rect 14323 33473 14335 33507
rect 14277 33467 14335 33473
rect 14553 33507 14611 33513
rect 14553 33473 14565 33507
rect 14599 33473 14611 33507
rect 14553 33467 14611 33473
rect 14182 33436 14188 33448
rect 12544 33408 13308 33436
rect 13740 33408 14188 33436
rect 12526 33368 12532 33380
rect 11348 33340 12532 33368
rect 11348 33309 11376 33340
rect 12526 33328 12532 33340
rect 12584 33328 12590 33380
rect 12802 33328 12808 33380
rect 12860 33328 12866 33380
rect 10928 33272 11192 33300
rect 11333 33303 11391 33309
rect 10928 33260 10934 33272
rect 11333 33269 11345 33303
rect 11379 33269 11391 33303
rect 11333 33263 11391 33269
rect 12158 33260 12164 33312
rect 12216 33300 12222 33312
rect 12820 33300 12848 33328
rect 13740 33312 13768 33408
rect 14182 33396 14188 33408
rect 14240 33436 14246 33448
rect 14292 33436 14320 33467
rect 14642 33464 14648 33516
rect 14700 33464 14706 33516
rect 14737 33507 14795 33513
rect 14737 33473 14749 33507
rect 14783 33504 14795 33507
rect 15194 33504 15200 33516
rect 14783 33476 15200 33504
rect 14783 33473 14795 33476
rect 14737 33467 14795 33473
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 15473 33507 15531 33513
rect 15473 33473 15485 33507
rect 15519 33504 15531 33507
rect 15654 33504 15660 33516
rect 15519 33476 15660 33504
rect 15519 33473 15531 33476
rect 15473 33467 15531 33473
rect 15654 33464 15660 33476
rect 15712 33464 15718 33516
rect 15948 33513 15976 33544
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 16224 33504 16252 33600
rect 16316 33572 16344 33600
rect 16316 33544 16436 33572
rect 16408 33513 16436 33544
rect 17494 33532 17500 33584
rect 17552 33532 17558 33584
rect 21284 33572 21312 33612
rect 21358 33600 21364 33612
rect 21416 33640 21422 33652
rect 21416 33612 21496 33640
rect 21416 33600 21422 33612
rect 17696 33544 21312 33572
rect 16301 33507 16359 33513
rect 16301 33504 16313 33507
rect 16224 33476 16313 33504
rect 16301 33473 16313 33476
rect 16347 33473 16359 33507
rect 16301 33467 16359 33473
rect 16393 33507 16451 33513
rect 16393 33473 16405 33507
rect 16439 33473 16451 33507
rect 16393 33467 16451 33473
rect 16574 33464 16580 33516
rect 16632 33504 16638 33516
rect 16853 33507 16911 33513
rect 16853 33504 16865 33507
rect 16632 33476 16865 33504
rect 16632 33464 16638 33476
rect 16853 33473 16865 33476
rect 16899 33473 16911 33507
rect 16853 33467 16911 33473
rect 17218 33464 17224 33516
rect 17276 33464 17282 33516
rect 17696 33513 17724 33544
rect 17681 33507 17739 33513
rect 17681 33473 17693 33507
rect 17727 33473 17739 33507
rect 17681 33467 17739 33473
rect 17862 33464 17868 33516
rect 17920 33504 17926 33516
rect 18233 33507 18291 33513
rect 18233 33504 18245 33507
rect 17920 33476 18245 33504
rect 17920 33464 17926 33476
rect 18233 33473 18245 33476
rect 18279 33473 18291 33507
rect 18233 33467 18291 33473
rect 18877 33507 18935 33513
rect 18877 33473 18889 33507
rect 18923 33473 18935 33507
rect 18877 33467 18935 33473
rect 14240 33408 14320 33436
rect 14660 33436 14688 33464
rect 14829 33439 14887 33445
rect 14829 33436 14841 33439
rect 14660 33408 14841 33436
rect 14240 33396 14246 33408
rect 14829 33405 14841 33408
rect 14875 33405 14887 33439
rect 14829 33399 14887 33405
rect 14918 33396 14924 33448
rect 14976 33436 14982 33448
rect 15565 33439 15623 33445
rect 15565 33436 15577 33439
rect 14976 33408 15577 33436
rect 14976 33396 14982 33408
rect 15565 33405 15577 33408
rect 15611 33405 15623 33439
rect 15565 33399 15623 33405
rect 15749 33439 15807 33445
rect 15749 33405 15761 33439
rect 15795 33436 15807 33439
rect 16206 33436 16212 33448
rect 15795 33408 16212 33436
rect 15795 33405 15807 33408
rect 15749 33399 15807 33405
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 16669 33439 16727 33445
rect 16669 33405 16681 33439
rect 16715 33436 16727 33439
rect 17954 33436 17960 33448
rect 16715 33408 17960 33436
rect 16715 33405 16727 33408
rect 16669 33399 16727 33405
rect 17954 33396 17960 33408
rect 18012 33396 18018 33448
rect 18506 33396 18512 33448
rect 18564 33396 18570 33448
rect 18892 33436 18920 33467
rect 19058 33464 19064 33516
rect 19116 33464 19122 33516
rect 19150 33464 19156 33516
rect 19208 33464 19214 33516
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19484 33476 19625 33504
rect 19484 33464 19490 33476
rect 19613 33473 19625 33476
rect 19659 33473 19671 33507
rect 19613 33467 19671 33473
rect 19880 33507 19938 33513
rect 19880 33473 19892 33507
rect 19926 33504 19938 33507
rect 20438 33504 20444 33516
rect 19926 33476 20444 33504
rect 19926 33473 19938 33476
rect 19880 33467 19938 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 21082 33464 21088 33516
rect 21140 33504 21146 33516
rect 21468 33513 21496 33612
rect 22370 33600 22376 33652
rect 22428 33640 22434 33652
rect 23385 33643 23443 33649
rect 23385 33640 23397 33643
rect 22428 33612 23397 33640
rect 22428 33600 22434 33612
rect 23385 33609 23397 33612
rect 23431 33609 23443 33643
rect 23385 33603 23443 33609
rect 24394 33600 24400 33652
rect 24452 33600 24458 33652
rect 25501 33643 25559 33649
rect 25501 33640 25513 33643
rect 24688 33612 25513 33640
rect 22002 33532 22008 33584
rect 22060 33532 22066 33584
rect 23014 33532 23020 33584
rect 23072 33532 23078 33584
rect 24210 33532 24216 33584
rect 24268 33572 24274 33584
rect 24688 33581 24716 33612
rect 25501 33609 25513 33612
rect 25547 33640 25559 33643
rect 27706 33640 27712 33652
rect 25547 33612 27712 33640
rect 25547 33609 25559 33612
rect 25501 33603 25559 33609
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 28074 33600 28080 33652
rect 28132 33640 28138 33652
rect 28132 33612 29960 33640
rect 28132 33600 28138 33612
rect 24673 33575 24731 33581
rect 24673 33572 24685 33575
rect 24268 33544 24685 33572
rect 24268 33532 24274 33544
rect 24673 33541 24685 33544
rect 24719 33541 24731 33575
rect 24673 33535 24731 33541
rect 24854 33532 24860 33584
rect 24912 33572 24918 33584
rect 26145 33575 26203 33581
rect 26145 33572 26157 33575
rect 24912 33544 26157 33572
rect 24912 33532 24918 33544
rect 26145 33541 26157 33544
rect 26191 33541 26203 33575
rect 26145 33535 26203 33541
rect 26513 33575 26571 33581
rect 26513 33541 26525 33575
rect 26559 33572 26571 33575
rect 26786 33572 26792 33584
rect 26559 33544 26792 33572
rect 26559 33541 26571 33544
rect 26513 33535 26571 33541
rect 26786 33532 26792 33544
rect 26844 33532 26850 33584
rect 27246 33532 27252 33584
rect 27304 33572 27310 33584
rect 27304 33544 27614 33572
rect 27304 33532 27310 33544
rect 21269 33507 21327 33513
rect 21269 33504 21281 33507
rect 21140 33476 21281 33504
rect 21140 33464 21146 33476
rect 21269 33473 21281 33476
rect 21315 33473 21327 33507
rect 21269 33467 21327 33473
rect 21434 33507 21496 33513
rect 21434 33473 21446 33507
rect 21480 33476 21496 33507
rect 21480 33473 21492 33476
rect 21434 33467 21492 33473
rect 21542 33464 21548 33516
rect 21600 33464 21606 33516
rect 21637 33507 21695 33513
rect 21637 33473 21649 33507
rect 21683 33504 21695 33507
rect 22020 33504 22048 33532
rect 21683 33476 22048 33504
rect 22272 33507 22330 33513
rect 21683 33473 21695 33476
rect 21637 33467 21695 33473
rect 22272 33473 22284 33507
rect 22318 33504 22330 33507
rect 23032 33504 23060 33532
rect 22318 33476 23060 33504
rect 22318 33473 22330 33476
rect 22272 33467 22330 33473
rect 23198 33464 23204 33516
rect 23256 33464 23262 33516
rect 23658 33464 23664 33516
rect 23716 33464 23722 33516
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 19168 33436 19196 33464
rect 18892 33408 19196 33436
rect 20898 33396 20904 33448
rect 20956 33436 20962 33448
rect 21910 33436 21916 33448
rect 20956 33408 21916 33436
rect 20956 33396 20962 33408
rect 21910 33396 21916 33408
rect 21968 33436 21974 33448
rect 22005 33439 22063 33445
rect 22005 33436 22017 33439
rect 21968 33408 22017 33436
rect 21968 33396 21974 33408
rect 22005 33405 22017 33408
rect 22051 33405 22063 33439
rect 23216 33436 23244 33464
rect 24044 33436 24072 33467
rect 24578 33464 24584 33516
rect 24636 33464 24642 33516
rect 24765 33507 24823 33513
rect 24765 33473 24777 33507
rect 24811 33473 24823 33507
rect 24872 33504 24900 33532
rect 24949 33507 25007 33513
rect 24949 33504 24961 33507
rect 24872 33476 24961 33504
rect 24765 33467 24823 33473
rect 24949 33473 24961 33476
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33504 25099 33507
rect 25222 33504 25228 33516
rect 25087 33476 25228 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 23216 33408 24072 33436
rect 24780 33436 24808 33467
rect 25222 33464 25228 33476
rect 25280 33464 25286 33516
rect 25317 33507 25375 33513
rect 25317 33473 25329 33507
rect 25363 33504 25375 33507
rect 25406 33504 25412 33516
rect 25363 33476 25412 33504
rect 25363 33473 25375 33476
rect 25317 33467 25375 33473
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 25777 33507 25835 33513
rect 25777 33504 25789 33507
rect 25648 33476 25789 33504
rect 25648 33464 25654 33476
rect 25777 33473 25789 33476
rect 25823 33473 25835 33507
rect 25777 33467 25835 33473
rect 26053 33507 26111 33513
rect 26053 33473 26065 33507
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 24854 33436 24860 33448
rect 24780 33408 24860 33436
rect 22005 33399 22063 33405
rect 24854 33396 24860 33408
rect 24912 33396 24918 33448
rect 25133 33439 25191 33445
rect 25133 33405 25145 33439
rect 25179 33436 25191 33439
rect 25682 33436 25688 33448
rect 25179 33408 25688 33436
rect 25179 33405 25191 33408
rect 25133 33399 25191 33405
rect 25682 33396 25688 33408
rect 25740 33396 25746 33448
rect 25866 33396 25872 33448
rect 25924 33396 25930 33448
rect 26068 33436 26096 33467
rect 26234 33464 26240 33516
rect 26292 33464 26298 33516
rect 26510 33436 26516 33448
rect 26068 33408 26516 33436
rect 26510 33396 26516 33408
rect 26568 33396 26574 33448
rect 26804 33436 26832 33532
rect 27586 33504 27614 33544
rect 28902 33532 28908 33584
rect 28960 33572 28966 33584
rect 29365 33575 29423 33581
rect 29365 33572 29377 33575
rect 28960 33544 29377 33572
rect 28960 33532 28966 33544
rect 29365 33541 29377 33544
rect 29411 33572 29423 33575
rect 29730 33572 29736 33584
rect 29411 33544 29736 33572
rect 29411 33541 29423 33544
rect 29365 33535 29423 33541
rect 29730 33532 29736 33544
rect 29788 33532 29794 33584
rect 27798 33504 27804 33516
rect 27586 33476 27804 33504
rect 27798 33464 27804 33476
rect 27856 33464 27862 33516
rect 28166 33464 28172 33516
rect 28224 33464 28230 33516
rect 28920 33504 28948 33532
rect 28828 33476 28948 33504
rect 27525 33439 27583 33445
rect 27525 33436 27537 33439
rect 26804 33408 27537 33436
rect 27525 33405 27537 33408
rect 27571 33405 27583 33439
rect 27525 33399 27583 33405
rect 28077 33439 28135 33445
rect 28077 33405 28089 33439
rect 28123 33436 28135 33439
rect 28534 33436 28540 33448
rect 28123 33408 28540 33436
rect 28123 33405 28135 33408
rect 28077 33399 28135 33405
rect 14734 33328 14740 33380
rect 14792 33368 14798 33380
rect 26234 33368 26240 33380
rect 14792 33340 15700 33368
rect 14792 33328 14798 33340
rect 12216 33272 12848 33300
rect 12216 33260 12222 33272
rect 13354 33260 13360 33312
rect 13412 33260 13418 33312
rect 13722 33260 13728 33312
rect 13780 33260 13786 33312
rect 14369 33303 14427 33309
rect 14369 33269 14381 33303
rect 14415 33300 14427 33303
rect 14642 33300 14648 33312
rect 14415 33272 14648 33300
rect 14415 33269 14427 33272
rect 14369 33263 14427 33269
rect 14642 33260 14648 33272
rect 14700 33260 14706 33312
rect 15105 33303 15163 33309
rect 15105 33269 15117 33303
rect 15151 33300 15163 33303
rect 15562 33300 15568 33312
rect 15151 33272 15568 33300
rect 15151 33269 15163 33272
rect 15105 33263 15163 33269
rect 15562 33260 15568 33272
rect 15620 33260 15626 33312
rect 15672 33300 15700 33340
rect 23584 33340 26240 33368
rect 23584 33312 23612 33340
rect 26234 33328 26240 33340
rect 26292 33328 26298 33380
rect 26326 33328 26332 33380
rect 26384 33368 26390 33380
rect 27338 33368 27344 33380
rect 26384 33340 27344 33368
rect 26384 33328 26390 33340
rect 27338 33328 27344 33340
rect 27396 33328 27402 33380
rect 27540 33368 27568 33399
rect 27985 33371 28043 33377
rect 27985 33368 27997 33371
rect 27540 33340 27997 33368
rect 27985 33337 27997 33340
rect 28031 33368 28043 33371
rect 28092 33368 28120 33399
rect 28534 33396 28540 33408
rect 28592 33436 28598 33448
rect 28828 33436 28856 33476
rect 28994 33464 29000 33516
rect 29052 33504 29058 33516
rect 29932 33513 29960 33612
rect 29641 33507 29699 33513
rect 29641 33504 29653 33507
rect 29052 33476 29653 33504
rect 29052 33464 29058 33476
rect 29641 33473 29653 33476
rect 29687 33473 29699 33507
rect 29641 33467 29699 33473
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 29825 33467 29883 33473
rect 29917 33507 29975 33513
rect 29917 33473 29929 33507
rect 29963 33473 29975 33507
rect 29917 33467 29975 33473
rect 28592 33408 28856 33436
rect 28592 33396 28598 33408
rect 28626 33368 28632 33380
rect 28031 33340 28120 33368
rect 28368 33340 28632 33368
rect 28031 33337 28043 33340
rect 27985 33331 28043 33337
rect 16761 33303 16819 33309
rect 16761 33300 16773 33303
rect 15672 33272 16773 33300
rect 16761 33269 16773 33272
rect 16807 33269 16819 33303
rect 16761 33263 16819 33269
rect 16850 33260 16856 33312
rect 16908 33300 16914 33312
rect 18874 33300 18880 33312
rect 16908 33272 18880 33300
rect 16908 33260 16914 33272
rect 18874 33260 18880 33272
rect 18932 33260 18938 33312
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20530 33300 20536 33312
rect 20036 33272 20536 33300
rect 20036 33260 20042 33272
rect 20530 33260 20536 33272
rect 20588 33300 20594 33312
rect 20993 33303 21051 33309
rect 20993 33300 21005 33303
rect 20588 33272 21005 33300
rect 20588 33260 20594 33272
rect 20993 33269 21005 33272
rect 21039 33269 21051 33303
rect 20993 33263 21051 33269
rect 21085 33303 21143 33309
rect 21085 33269 21097 33303
rect 21131 33300 21143 33303
rect 22370 33300 22376 33312
rect 21131 33272 22376 33300
rect 21131 33269 21143 33272
rect 21085 33263 21143 33269
rect 22370 33260 22376 33272
rect 22428 33260 22434 33312
rect 23566 33260 23572 33312
rect 23624 33260 23630 33312
rect 25682 33260 25688 33312
rect 25740 33300 25746 33312
rect 26878 33300 26884 33312
rect 25740 33272 26884 33300
rect 25740 33260 25746 33272
rect 26878 33260 26884 33272
rect 26936 33300 26942 33312
rect 27157 33303 27215 33309
rect 27157 33300 27169 33303
rect 26936 33272 27169 33300
rect 26936 33260 26942 33272
rect 27157 33269 27169 33272
rect 27203 33269 27215 33303
rect 27157 33263 27215 33269
rect 27706 33260 27712 33312
rect 27764 33300 27770 33312
rect 28258 33300 28264 33312
rect 27764 33272 28264 33300
rect 27764 33260 27770 33272
rect 28258 33260 28264 33272
rect 28316 33260 28322 33312
rect 28368 33309 28396 33340
rect 28626 33328 28632 33340
rect 28684 33368 28690 33380
rect 29840 33368 29868 33467
rect 30009 33439 30067 33445
rect 30009 33436 30021 33439
rect 28684 33340 29868 33368
rect 29932 33408 30021 33436
rect 28684 33328 28690 33340
rect 29932 33312 29960 33408
rect 30009 33405 30021 33408
rect 30055 33405 30067 33439
rect 30009 33399 30067 33405
rect 28353 33303 28411 33309
rect 28353 33269 28365 33303
rect 28399 33269 28411 33303
rect 28353 33263 28411 33269
rect 29454 33260 29460 33312
rect 29512 33260 29518 33312
rect 29914 33260 29920 33312
rect 29972 33260 29978 33312
rect 30466 33260 30472 33312
rect 30524 33300 30530 33312
rect 30653 33303 30711 33309
rect 30653 33300 30665 33303
rect 30524 33272 30665 33300
rect 30524 33260 30530 33272
rect 30653 33269 30665 33272
rect 30699 33269 30711 33303
rect 30653 33263 30711 33269
rect 1104 33210 43884 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 43884 33210
rect 1104 33136 43884 33158
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 3237 33099 3295 33105
rect 3237 33096 3249 33099
rect 2924 33068 3249 33096
rect 2924 33056 2930 33068
rect 3237 33065 3249 33068
rect 3283 33065 3295 33099
rect 3237 33059 3295 33065
rect 3513 33099 3571 33105
rect 3513 33065 3525 33099
rect 3559 33096 3571 33099
rect 3970 33096 3976 33108
rect 3559 33068 3976 33096
rect 3559 33065 3571 33068
rect 3513 33059 3571 33065
rect 3970 33056 3976 33068
rect 4028 33056 4034 33108
rect 5997 33099 6055 33105
rect 5997 33065 6009 33099
rect 6043 33096 6055 33099
rect 6270 33096 6276 33108
rect 6043 33068 6276 33096
rect 6043 33065 6055 33068
rect 5997 33059 6055 33065
rect 6270 33056 6276 33068
rect 6328 33096 6334 33108
rect 6638 33096 6644 33108
rect 6328 33068 6644 33096
rect 6328 33056 6334 33068
rect 6638 33056 6644 33068
rect 6696 33056 6702 33108
rect 9125 33099 9183 33105
rect 9125 33065 9137 33099
rect 9171 33096 9183 33099
rect 9214 33096 9220 33108
rect 9171 33068 9220 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 9214 33056 9220 33068
rect 9272 33056 9278 33108
rect 9398 33056 9404 33108
rect 9456 33056 9462 33108
rect 10413 33099 10471 33105
rect 10413 33065 10425 33099
rect 10459 33096 10471 33099
rect 10502 33096 10508 33108
rect 10459 33068 10508 33096
rect 10459 33065 10471 33068
rect 10413 33059 10471 33065
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 10594 33056 10600 33108
rect 10652 33096 10658 33108
rect 10689 33099 10747 33105
rect 10689 33096 10701 33099
rect 10652 33068 10701 33096
rect 10652 33056 10658 33068
rect 10689 33065 10701 33068
rect 10735 33096 10747 33099
rect 11609 33099 11667 33105
rect 11609 33096 11621 33099
rect 10735 33068 11621 33096
rect 10735 33065 10747 33068
rect 10689 33059 10747 33065
rect 1762 32960 1768 32972
rect 1412 32932 1768 32960
rect 1412 32901 1440 32932
rect 1762 32920 1768 32932
rect 1820 32960 1826 32972
rect 1820 32932 1992 32960
rect 1820 32920 1826 32932
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1854 32852 1860 32904
rect 1912 32852 1918 32904
rect 1964 32892 1992 32932
rect 8662 32920 8668 32972
rect 8720 32960 8726 32972
rect 9232 32960 9260 33056
rect 10045 32963 10103 32969
rect 10045 32960 10057 32963
rect 8720 32932 8984 32960
rect 9232 32932 10057 32960
rect 8720 32920 8726 32932
rect 2682 32892 2688 32904
rect 1964 32864 2688 32892
rect 2682 32852 2688 32864
rect 2740 32852 2746 32904
rect 3421 32895 3479 32901
rect 3421 32861 3433 32895
rect 3467 32892 3479 32895
rect 4522 32892 4528 32904
rect 3467 32864 4528 32892
rect 3467 32861 3479 32864
rect 3421 32855 3479 32861
rect 4522 32852 4528 32864
rect 4580 32852 4586 32904
rect 4617 32895 4675 32901
rect 4617 32861 4629 32895
rect 4663 32892 4675 32895
rect 6365 32895 6423 32901
rect 6365 32892 6377 32895
rect 4663 32864 6377 32892
rect 4663 32861 4675 32864
rect 4617 32855 4675 32861
rect 6365 32861 6377 32864
rect 6411 32892 6423 32895
rect 7006 32892 7012 32904
rect 6411 32864 7012 32892
rect 6411 32861 6423 32864
rect 6365 32855 6423 32861
rect 934 32716 940 32768
rect 992 32756 998 32768
rect 1581 32759 1639 32765
rect 1581 32756 1593 32759
rect 992 32728 1593 32756
rect 992 32716 998 32728
rect 1581 32725 1593 32728
rect 1627 32725 1639 32759
rect 1872 32756 1900 32852
rect 2130 32833 2136 32836
rect 2124 32824 2136 32833
rect 2091 32796 2136 32824
rect 2124 32787 2136 32796
rect 2130 32784 2136 32787
rect 2188 32784 2194 32836
rect 4632 32824 4660 32855
rect 7006 32852 7012 32864
rect 7064 32852 7070 32904
rect 7926 32852 7932 32904
rect 7984 32852 7990 32904
rect 8205 32895 8263 32901
rect 8205 32861 8217 32895
rect 8251 32861 8263 32895
rect 8205 32855 8263 32861
rect 2240 32796 4660 32824
rect 2240 32756 2268 32796
rect 4706 32784 4712 32836
rect 4764 32824 4770 32836
rect 4862 32827 4920 32833
rect 4862 32824 4874 32827
rect 4764 32796 4874 32824
rect 4764 32784 4770 32796
rect 4862 32793 4874 32796
rect 4908 32793 4920 32827
rect 4862 32787 4920 32793
rect 6632 32827 6690 32833
rect 6632 32793 6644 32827
rect 6678 32824 6690 32827
rect 7944 32824 7972 32852
rect 6678 32796 7972 32824
rect 8220 32824 8248 32855
rect 8386 32852 8392 32904
rect 8444 32892 8450 32904
rect 8846 32892 8852 32904
rect 8444 32864 8852 32892
rect 8444 32852 8450 32864
rect 8846 32852 8852 32864
rect 8904 32852 8910 32904
rect 8956 32901 8984 32932
rect 10045 32929 10057 32932
rect 10091 32960 10103 32963
rect 11164 32960 11192 33068
rect 11609 33065 11621 33068
rect 11655 33065 11667 33099
rect 11609 33059 11667 33065
rect 11698 33056 11704 33108
rect 11756 33096 11762 33108
rect 12621 33099 12679 33105
rect 11756 33068 12572 33096
rect 11756 33056 11762 33068
rect 11238 32988 11244 33040
rect 11296 33028 11302 33040
rect 12345 33031 12403 33037
rect 11296 33000 12204 33028
rect 11296 32988 11302 33000
rect 11885 32963 11943 32969
rect 11885 32960 11897 32963
rect 10091 32932 10732 32960
rect 11164 32932 11897 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 8941 32895 8999 32901
rect 8941 32861 8953 32895
rect 8987 32861 8999 32895
rect 8941 32855 8999 32861
rect 9034 32895 9092 32901
rect 9034 32861 9046 32895
rect 9080 32892 9092 32895
rect 9214 32894 9220 32904
rect 9140 32892 9220 32894
rect 9080 32866 9220 32892
rect 9080 32864 9168 32866
rect 9201 32864 9220 32866
rect 9080 32861 9092 32864
rect 9034 32855 9092 32861
rect 9214 32852 9220 32864
rect 9272 32852 9278 32904
rect 9766 32852 9772 32904
rect 9824 32852 9830 32904
rect 10704 32901 10732 32932
rect 11885 32929 11897 32932
rect 11931 32929 11943 32963
rect 11885 32923 11943 32929
rect 12176 32904 12204 33000
rect 12345 32997 12357 33031
rect 12391 32997 12403 33031
rect 12544 33028 12572 33068
rect 12621 33065 12633 33099
rect 12667 33096 12679 33099
rect 12710 33096 12716 33108
rect 12667 33068 12716 33096
rect 12667 33065 12679 33068
rect 12621 33059 12679 33065
rect 12710 33056 12716 33068
rect 12768 33096 12774 33108
rect 13354 33096 13360 33108
rect 12768 33068 13360 33096
rect 12768 33056 12774 33068
rect 13354 33056 13360 33068
rect 13412 33056 13418 33108
rect 13630 33056 13636 33108
rect 13688 33096 13694 33108
rect 13817 33099 13875 33105
rect 13817 33096 13829 33099
rect 13688 33068 13829 33096
rect 13688 33056 13694 33068
rect 13817 33065 13829 33068
rect 13863 33065 13875 33099
rect 16209 33099 16267 33105
rect 16209 33096 16221 33099
rect 13817 33059 13875 33065
rect 14108 33068 16221 33096
rect 12544 33000 13492 33028
rect 12345 32991 12403 32997
rect 12250 32920 12256 32972
rect 12308 32920 12314 32972
rect 12360 32960 12388 32991
rect 12894 32960 12900 32972
rect 12360 32932 12900 32960
rect 12894 32920 12900 32932
rect 12952 32920 12958 32972
rect 13262 32920 13268 32972
rect 13320 32920 13326 32972
rect 13464 32969 13492 33000
rect 13449 32963 13507 32969
rect 13449 32929 13461 32963
rect 13495 32929 13507 32963
rect 13449 32923 13507 32929
rect 10689 32895 10747 32901
rect 10689 32861 10701 32895
rect 10735 32861 10747 32895
rect 10689 32855 10747 32861
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32861 10931 32895
rect 10873 32855 10931 32861
rect 10229 32827 10287 32833
rect 8220 32796 9996 32824
rect 6678 32793 6690 32796
rect 6632 32787 6690 32793
rect 1872 32728 2268 32756
rect 1581 32719 1639 32725
rect 3970 32716 3976 32768
rect 4028 32716 4034 32768
rect 4062 32716 4068 32768
rect 4120 32756 4126 32768
rect 4525 32759 4583 32765
rect 4525 32756 4537 32759
rect 4120 32728 4537 32756
rect 4120 32716 4126 32728
rect 4525 32725 4537 32728
rect 4571 32756 4583 32759
rect 5350 32756 5356 32768
rect 4571 32728 5356 32756
rect 4571 32725 4583 32728
rect 4525 32719 4583 32725
rect 5350 32716 5356 32728
rect 5408 32716 5414 32768
rect 5902 32716 5908 32768
rect 5960 32756 5966 32768
rect 7466 32756 7472 32768
rect 5960 32728 7472 32756
rect 5960 32716 5966 32728
rect 7466 32716 7472 32728
rect 7524 32716 7530 32768
rect 7745 32759 7803 32765
rect 7745 32725 7757 32759
rect 7791 32756 7803 32759
rect 8220 32756 8248 32796
rect 7791 32728 8248 32756
rect 7791 32725 7803 32728
rect 7745 32719 7803 32725
rect 8294 32716 8300 32768
rect 8352 32756 8358 32768
rect 8757 32759 8815 32765
rect 8757 32756 8769 32759
rect 8352 32728 8769 32756
rect 8352 32716 8358 32728
rect 8757 32725 8769 32728
rect 8803 32725 8815 32759
rect 8757 32719 8815 32725
rect 8846 32716 8852 32768
rect 8904 32756 8910 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 8904 32728 9873 32756
rect 8904 32716 8910 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9968 32756 9996 32796
rect 10229 32793 10241 32827
rect 10275 32824 10287 32827
rect 10318 32824 10324 32836
rect 10275 32796 10324 32824
rect 10275 32793 10287 32796
rect 10229 32787 10287 32793
rect 10318 32784 10324 32796
rect 10376 32784 10382 32836
rect 10888 32824 10916 32855
rect 11054 32852 11060 32904
rect 11112 32892 11118 32904
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 11112 32864 11437 32892
rect 11112 32852 11118 32864
rect 11425 32861 11437 32864
rect 11471 32892 11483 32895
rect 11606 32892 11612 32904
rect 11471 32864 11612 32892
rect 11471 32861 11483 32864
rect 11425 32855 11483 32861
rect 11606 32852 11612 32864
rect 11664 32852 11670 32904
rect 11701 32895 11759 32901
rect 11701 32861 11713 32895
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 10520 32796 10916 32824
rect 10429 32759 10487 32765
rect 10429 32756 10441 32759
rect 9968 32728 10441 32756
rect 9861 32719 9919 32725
rect 10429 32725 10441 32728
rect 10475 32756 10487 32759
rect 10520 32756 10548 32796
rect 11514 32784 11520 32836
rect 11572 32824 11578 32836
rect 11716 32824 11744 32855
rect 11790 32852 11796 32904
rect 11848 32892 11854 32904
rect 11977 32895 12035 32901
rect 11977 32892 11989 32895
rect 11848 32864 11989 32892
rect 11848 32852 11854 32864
rect 11977 32861 11989 32864
rect 12023 32861 12035 32895
rect 11977 32855 12035 32861
rect 12158 32852 12164 32904
rect 12216 32852 12222 32904
rect 12268 32824 12296 32920
rect 14108 32904 14136 33068
rect 16209 33065 16221 33068
rect 16255 33065 16267 33099
rect 16209 33059 16267 33065
rect 16298 33056 16304 33108
rect 16356 33096 16362 33108
rect 16850 33096 16856 33108
rect 16356 33068 16856 33096
rect 16356 33056 16362 33068
rect 16850 33056 16856 33068
rect 16908 33056 16914 33108
rect 19978 33096 19984 33108
rect 17696 33068 19984 33096
rect 16390 33028 16396 33040
rect 15861 33000 16396 33028
rect 13541 32895 13599 32901
rect 13541 32861 13553 32895
rect 13587 32892 13599 32895
rect 13906 32892 13912 32904
rect 13587 32864 13912 32892
rect 13587 32861 13599 32864
rect 13541 32855 13599 32861
rect 13906 32852 13912 32864
rect 13964 32852 13970 32904
rect 14090 32894 14096 32904
rect 14016 32866 14096 32894
rect 11572 32796 12296 32824
rect 11572 32784 11578 32796
rect 12342 32784 12348 32836
rect 12400 32824 12406 32836
rect 12437 32827 12495 32833
rect 12437 32824 12449 32827
rect 12400 32796 12449 32824
rect 12400 32784 12406 32796
rect 12437 32793 12449 32796
rect 12483 32793 12495 32827
rect 12437 32787 12495 32793
rect 12526 32784 12532 32836
rect 12584 32824 12590 32836
rect 12637 32827 12695 32833
rect 12637 32824 12649 32827
rect 12584 32796 12649 32824
rect 12584 32784 12590 32796
rect 12637 32793 12649 32796
rect 12683 32793 12695 32827
rect 14016 32824 14044 32866
rect 14090 32852 14096 32866
rect 14148 32852 14154 32904
rect 14829 32895 14887 32901
rect 14829 32861 14841 32895
rect 14875 32892 14887 32895
rect 15654 32892 15660 32904
rect 14875 32864 15660 32892
rect 14875 32861 14887 32864
rect 14829 32855 14887 32861
rect 15654 32852 15660 32864
rect 15712 32892 15718 32904
rect 15861 32892 15889 33000
rect 16390 32988 16396 33000
rect 16448 32988 16454 33040
rect 17696 33037 17724 33068
rect 19978 33056 19984 33068
rect 20036 33056 20042 33108
rect 20070 33056 20076 33108
rect 20128 33096 20134 33108
rect 21818 33096 21824 33108
rect 20128 33068 21824 33096
rect 20128 33056 20134 33068
rect 21818 33056 21824 33068
rect 21876 33056 21882 33108
rect 22186 33056 22192 33108
rect 22244 33096 22250 33108
rect 22281 33099 22339 33105
rect 22281 33096 22293 33099
rect 22244 33068 22293 33096
rect 22244 33056 22250 33068
rect 22281 33065 22293 33068
rect 22327 33065 22339 33099
rect 22281 33059 22339 33065
rect 24670 33056 24676 33108
rect 24728 33096 24734 33108
rect 25501 33099 25559 33105
rect 25501 33096 25513 33099
rect 24728 33068 25513 33096
rect 24728 33056 24734 33068
rect 25501 33065 25513 33068
rect 25547 33096 25559 33099
rect 25958 33096 25964 33108
rect 25547 33068 25964 33096
rect 25547 33065 25559 33068
rect 25501 33059 25559 33065
rect 25958 33056 25964 33068
rect 26016 33056 26022 33108
rect 26142 33056 26148 33108
rect 26200 33096 26206 33108
rect 26418 33096 26424 33108
rect 26200 33068 26424 33096
rect 26200 33056 26206 33068
rect 26418 33056 26424 33068
rect 26476 33096 26482 33108
rect 26786 33096 26792 33108
rect 26476 33068 26792 33096
rect 26476 33056 26482 33068
rect 26786 33056 26792 33068
rect 26844 33056 26850 33108
rect 27890 33056 27896 33108
rect 27948 33056 27954 33108
rect 28534 33056 28540 33108
rect 28592 33056 28598 33108
rect 29270 33056 29276 33108
rect 29328 33096 29334 33108
rect 29546 33096 29552 33108
rect 29328 33068 29552 33096
rect 29328 33056 29334 33068
rect 29546 33056 29552 33068
rect 29604 33056 29610 33108
rect 17681 33031 17739 33037
rect 17681 32997 17693 33031
rect 17727 32997 17739 33031
rect 18138 33028 18144 33040
rect 17681 32991 17739 32997
rect 17880 33000 18144 33028
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 17497 32963 17555 32969
rect 17497 32960 17509 32963
rect 16264 32932 17509 32960
rect 16264 32920 16270 32932
rect 17497 32929 17509 32932
rect 17543 32960 17555 32963
rect 17880 32960 17908 33000
rect 18138 32988 18144 33000
rect 18196 32988 18202 33040
rect 18233 33031 18291 33037
rect 18233 32997 18245 33031
rect 18279 33028 18291 33031
rect 18598 33028 18604 33040
rect 18279 33000 18604 33028
rect 18279 32997 18291 33000
rect 18233 32991 18291 32997
rect 18598 32988 18604 33000
rect 18656 32988 18662 33040
rect 20809 33031 20867 33037
rect 20809 33028 20821 33031
rect 19720 33000 20821 33028
rect 17543 32932 17908 32960
rect 17972 32932 19196 32960
rect 17543 32929 17555 32932
rect 17497 32923 17555 32929
rect 15712 32864 15889 32892
rect 15712 32852 15718 32864
rect 15930 32852 15936 32904
rect 15988 32892 15994 32904
rect 16393 32895 16451 32901
rect 16393 32892 16405 32895
rect 15988 32864 16405 32892
rect 15988 32852 15994 32864
rect 16393 32861 16405 32864
rect 16439 32861 16451 32895
rect 16393 32855 16451 32861
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 17770 32892 17776 32904
rect 16540 32864 17776 32892
rect 16540 32852 16546 32864
rect 17770 32852 17776 32864
rect 17828 32852 17834 32904
rect 17972 32901 18000 32932
rect 19168 32904 19196 32932
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 18414 32852 18420 32904
rect 18472 32852 18478 32904
rect 19058 32852 19064 32904
rect 19116 32852 19122 32904
rect 19150 32852 19156 32904
rect 19208 32852 19214 32904
rect 19720 32901 19748 33000
rect 20809 32997 20821 33000
rect 20855 32997 20867 33031
rect 25685 33031 25743 33037
rect 25685 33028 25697 33031
rect 20809 32991 20867 32997
rect 22066 33000 25697 33028
rect 19978 32960 19984 32972
rect 19812 32932 19984 32960
rect 19812 32901 19840 32932
rect 19978 32920 19984 32932
rect 20036 32920 20042 32972
rect 20162 32960 20168 32972
rect 20088 32932 20168 32960
rect 20088 32901 20116 32932
rect 20162 32920 20168 32932
rect 20220 32920 20226 32972
rect 20530 32920 20536 32972
rect 20588 32920 20594 32972
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 19797 32895 19855 32901
rect 19797 32861 19809 32895
rect 19843 32861 19855 32895
rect 19797 32855 19855 32861
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 20073 32895 20131 32901
rect 20073 32861 20085 32895
rect 20119 32861 20131 32895
rect 20073 32855 20131 32861
rect 20257 32895 20315 32901
rect 20257 32861 20269 32895
rect 20303 32892 20315 32895
rect 20548 32892 20576 32920
rect 20303 32864 20576 32892
rect 20303 32861 20315 32864
rect 20257 32855 20315 32861
rect 12637 32787 12695 32793
rect 12729 32796 14044 32824
rect 15096 32827 15154 32833
rect 10475 32728 10548 32756
rect 10597 32759 10655 32765
rect 10475 32725 10487 32728
rect 10429 32719 10487 32725
rect 10597 32725 10609 32759
rect 10643 32756 10655 32759
rect 10686 32756 10692 32768
rect 10643 32728 10692 32756
rect 10643 32725 10655 32728
rect 10597 32719 10655 32725
rect 10686 32716 10692 32728
rect 10744 32716 10750 32768
rect 12066 32716 12072 32768
rect 12124 32756 12130 32768
rect 12729 32756 12757 32796
rect 15096 32793 15108 32827
rect 15142 32824 15154 32827
rect 18049 32827 18107 32833
rect 15142 32796 16988 32824
rect 15142 32793 15154 32796
rect 15096 32787 15154 32793
rect 16960 32768 16988 32796
rect 18049 32793 18061 32827
rect 18095 32824 18107 32827
rect 18506 32824 18512 32836
rect 18095 32796 18512 32824
rect 18095 32793 18107 32796
rect 18049 32787 18107 32793
rect 18506 32784 18512 32796
rect 18564 32824 18570 32836
rect 19076 32824 19104 32852
rect 18564 32796 19104 32824
rect 19904 32824 19932 32855
rect 20898 32852 20904 32904
rect 20956 32852 20962 32904
rect 22066 32892 22094 33000
rect 25685 32997 25697 33000
rect 25731 32997 25743 33031
rect 25685 32991 25743 32997
rect 26237 33031 26295 33037
rect 26237 32997 26249 33031
rect 26283 33028 26295 33031
rect 26283 33000 27844 33028
rect 26283 32997 26295 33000
rect 26237 32991 26295 32997
rect 22370 32920 22376 32972
rect 22428 32920 22434 32972
rect 27338 32960 27344 32972
rect 25148 32932 27344 32960
rect 21100 32864 22094 32892
rect 21100 32824 21128 32864
rect 23198 32852 23204 32904
rect 23256 32892 23262 32904
rect 23293 32895 23351 32901
rect 23293 32892 23305 32895
rect 23256 32864 23305 32892
rect 23256 32852 23262 32864
rect 23293 32861 23305 32864
rect 23339 32861 23351 32895
rect 23293 32855 23351 32861
rect 23569 32895 23627 32901
rect 23569 32861 23581 32895
rect 23615 32892 23627 32895
rect 23934 32892 23940 32904
rect 23615 32864 23940 32892
rect 23615 32861 23627 32864
rect 23569 32855 23627 32861
rect 23934 32852 23940 32864
rect 23992 32852 23998 32904
rect 24486 32852 24492 32904
rect 24544 32852 24550 32904
rect 25148 32901 25176 32932
rect 27338 32920 27344 32932
rect 27396 32920 27402 32972
rect 27614 32960 27620 32972
rect 27448 32932 27620 32960
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 25409 32855 25467 32861
rect 19904 32796 21128 32824
rect 21168 32827 21226 32833
rect 18564 32784 18570 32796
rect 21168 32793 21180 32827
rect 21214 32824 21226 32827
rect 23017 32827 23075 32833
rect 23017 32824 23029 32827
rect 21214 32796 23029 32824
rect 21214 32793 21226 32796
rect 21168 32787 21226 32793
rect 23017 32793 23029 32796
rect 23063 32793 23075 32827
rect 23017 32787 23075 32793
rect 24121 32827 24179 32833
rect 24121 32793 24133 32827
rect 24167 32793 24179 32827
rect 24121 32787 24179 32793
rect 12124 32728 12757 32756
rect 12124 32716 12130 32728
rect 12802 32716 12808 32768
rect 12860 32716 12866 32768
rect 14737 32759 14795 32765
rect 14737 32725 14749 32759
rect 14783 32756 14795 32759
rect 15654 32756 15660 32768
rect 14783 32728 15660 32756
rect 14783 32725 14795 32728
rect 14737 32719 14795 32725
rect 15654 32716 15660 32728
rect 15712 32716 15718 32768
rect 16942 32716 16948 32768
rect 17000 32716 17006 32768
rect 17034 32716 17040 32768
rect 17092 32716 17098 32768
rect 17126 32716 17132 32768
rect 17184 32756 17190 32768
rect 17862 32756 17868 32768
rect 17184 32728 17868 32756
rect 17184 32716 17190 32728
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 19058 32716 19064 32768
rect 19116 32716 19122 32768
rect 19429 32759 19487 32765
rect 19429 32725 19441 32759
rect 19475 32756 19487 32759
rect 19978 32756 19984 32768
rect 19475 32728 19984 32756
rect 19475 32725 19487 32728
rect 19429 32719 19487 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20070 32716 20076 32768
rect 20128 32756 20134 32768
rect 24136 32756 24164 32787
rect 24854 32784 24860 32836
rect 24912 32824 24918 32836
rect 25424 32824 25452 32855
rect 25498 32852 25504 32904
rect 25556 32852 25562 32904
rect 25774 32852 25780 32904
rect 25832 32892 25838 32904
rect 26053 32895 26111 32901
rect 26053 32892 26065 32895
rect 25832 32864 26065 32892
rect 25832 32852 25838 32864
rect 26053 32861 26065 32864
rect 26099 32861 26111 32895
rect 26053 32855 26111 32861
rect 26234 32852 26240 32904
rect 26292 32852 26298 32904
rect 26329 32895 26387 32901
rect 26329 32861 26341 32895
rect 26375 32892 26387 32895
rect 26418 32892 26424 32904
rect 26375 32864 26424 32892
rect 26375 32861 26387 32864
rect 26329 32855 26387 32861
rect 26418 32852 26424 32864
rect 26476 32852 26482 32904
rect 26881 32895 26939 32901
rect 26881 32892 26893 32895
rect 26528 32864 26893 32892
rect 24912 32796 25452 32824
rect 25516 32824 25544 32852
rect 25869 32827 25927 32833
rect 25869 32824 25881 32827
rect 25516 32796 25881 32824
rect 24912 32784 24918 32796
rect 25869 32793 25881 32796
rect 25915 32793 25927 32827
rect 26252 32824 26280 32852
rect 26528 32824 26556 32864
rect 26881 32861 26893 32864
rect 26927 32861 26939 32895
rect 26881 32855 26939 32861
rect 26970 32852 26976 32904
rect 27028 32892 27034 32904
rect 27448 32901 27476 32932
rect 27614 32920 27620 32932
rect 27672 32920 27678 32972
rect 27816 32960 27844 33000
rect 28902 32960 28908 32972
rect 27816 32932 28908 32960
rect 27816 32904 27844 32932
rect 28902 32920 28908 32932
rect 28960 32920 28966 32972
rect 29270 32920 29276 32972
rect 29328 32920 29334 32972
rect 29362 32920 29368 32972
rect 29420 32960 29426 32972
rect 29825 32963 29883 32969
rect 29825 32960 29837 32963
rect 29420 32932 29837 32960
rect 29420 32920 29426 32932
rect 29825 32929 29837 32932
rect 29871 32929 29883 32963
rect 29825 32923 29883 32929
rect 27065 32895 27123 32901
rect 27065 32892 27077 32895
rect 27028 32864 27077 32892
rect 27028 32852 27034 32864
rect 27065 32861 27077 32864
rect 27111 32861 27123 32895
rect 27065 32855 27123 32861
rect 27433 32895 27491 32901
rect 27433 32861 27445 32895
rect 27479 32861 27491 32895
rect 27433 32855 27491 32861
rect 27522 32852 27528 32904
rect 27580 32852 27586 32904
rect 27706 32852 27712 32904
rect 27764 32852 27770 32904
rect 27798 32852 27804 32904
rect 27856 32852 27862 32904
rect 28169 32895 28227 32901
rect 28169 32861 28181 32895
rect 28215 32892 28227 32895
rect 28442 32892 28448 32904
rect 28215 32864 28448 32892
rect 28215 32861 28227 32864
rect 28169 32855 28227 32861
rect 28442 32852 28448 32864
rect 28500 32852 28506 32904
rect 29086 32852 29092 32904
rect 29144 32852 29150 32904
rect 29181 32895 29239 32901
rect 29181 32861 29193 32895
rect 29227 32892 29239 32895
rect 29288 32892 29316 32920
rect 29730 32892 29736 32904
rect 29227 32864 29736 32892
rect 29227 32861 29239 32864
rect 29181 32855 29239 32861
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 29840 32892 29868 32923
rect 30374 32892 30380 32904
rect 29840 32864 30380 32892
rect 30374 32852 30380 32864
rect 30432 32852 30438 32904
rect 26252 32796 26556 32824
rect 26605 32827 26663 32833
rect 25869 32787 25927 32793
rect 26605 32793 26617 32827
rect 26651 32824 26663 32827
rect 27893 32827 27951 32833
rect 27893 32824 27905 32827
rect 26651 32796 27905 32824
rect 26651 32793 26663 32796
rect 26605 32787 26663 32793
rect 27893 32793 27905 32796
rect 27939 32824 27951 32827
rect 28994 32824 29000 32836
rect 27939 32796 29000 32824
rect 27939 32793 27951 32796
rect 27893 32787 27951 32793
rect 24578 32756 24584 32768
rect 20128 32728 24584 32756
rect 20128 32716 20134 32728
rect 24578 32716 24584 32728
rect 24636 32716 24642 32768
rect 25038 32716 25044 32768
rect 25096 32716 25102 32768
rect 26418 32716 26424 32768
rect 26476 32756 26482 32768
rect 26620 32756 26648 32787
rect 28994 32784 29000 32796
rect 29052 32824 29058 32836
rect 29270 32824 29276 32836
rect 29052 32796 29276 32824
rect 29052 32784 29058 32796
rect 29270 32784 29276 32796
rect 29328 32784 29334 32836
rect 29362 32784 29368 32836
rect 29420 32784 29426 32836
rect 29638 32784 29644 32836
rect 29696 32824 29702 32836
rect 30070 32827 30128 32833
rect 30070 32824 30082 32827
rect 29696 32796 30082 32824
rect 29696 32784 29702 32796
rect 30070 32793 30082 32796
rect 30116 32793 30128 32827
rect 30070 32787 30128 32793
rect 26476 32728 26648 32756
rect 26476 32716 26482 32728
rect 26694 32716 26700 32768
rect 26752 32756 26758 32768
rect 26878 32756 26884 32768
rect 26752 32728 26884 32756
rect 26752 32716 26758 32728
rect 26878 32716 26884 32728
rect 26936 32756 26942 32768
rect 26973 32759 27031 32765
rect 26973 32756 26985 32759
rect 26936 32728 26985 32756
rect 26936 32716 26942 32728
rect 26973 32725 26985 32728
rect 27019 32725 27031 32759
rect 26973 32719 27031 32725
rect 27246 32716 27252 32768
rect 27304 32716 27310 32768
rect 28077 32759 28135 32765
rect 28077 32725 28089 32759
rect 28123 32756 28135 32759
rect 28166 32756 28172 32768
rect 28123 32728 28172 32756
rect 28123 32725 28135 32728
rect 28077 32719 28135 32725
rect 28166 32716 28172 32728
rect 28224 32756 28230 32768
rect 28718 32756 28724 32768
rect 28224 32728 28724 32756
rect 28224 32716 28230 32728
rect 28718 32716 28724 32728
rect 28776 32716 28782 32768
rect 28810 32716 28816 32768
rect 28868 32716 28874 32768
rect 29914 32716 29920 32768
rect 29972 32756 29978 32768
rect 31205 32759 31263 32765
rect 31205 32756 31217 32759
rect 29972 32728 31217 32756
rect 29972 32716 29978 32728
rect 31205 32725 31217 32728
rect 31251 32725 31263 32759
rect 31205 32719 31263 32725
rect 1104 32666 43884 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 43884 32666
rect 1104 32592 43884 32614
rect 7374 32512 7380 32564
rect 7432 32552 7438 32564
rect 7929 32555 7987 32561
rect 7929 32552 7941 32555
rect 7432 32524 7941 32552
rect 7432 32512 7438 32524
rect 7929 32521 7941 32524
rect 7975 32521 7987 32555
rect 7929 32515 7987 32521
rect 8294 32512 8300 32564
rect 8352 32512 8358 32564
rect 9306 32552 9312 32564
rect 8588 32524 9312 32552
rect 4632 32456 6408 32484
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 1670 32416 1676 32428
rect 1627 32388 1676 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 4632 32425 4660 32456
rect 3697 32419 3755 32425
rect 3697 32385 3709 32419
rect 3743 32416 3755 32419
rect 4617 32419 4675 32425
rect 3743 32388 4568 32416
rect 3743 32385 3755 32388
rect 3697 32379 3755 32385
rect 1486 32308 1492 32360
rect 1544 32348 1550 32360
rect 1857 32351 1915 32357
rect 1857 32348 1869 32351
rect 1544 32320 1869 32348
rect 1544 32308 1550 32320
rect 1857 32317 1869 32320
rect 1903 32317 1915 32351
rect 1857 32311 1915 32317
rect 2958 32308 2964 32360
rect 3016 32308 3022 32360
rect 3973 32351 4031 32357
rect 3973 32317 3985 32351
rect 4019 32348 4031 32351
rect 4540 32348 4568 32388
rect 4617 32385 4629 32419
rect 4663 32385 4675 32419
rect 4617 32379 4675 32385
rect 4884 32419 4942 32425
rect 4884 32385 4896 32419
rect 4930 32416 4942 32419
rect 5626 32416 5632 32428
rect 4930 32388 5632 32416
rect 4930 32385 4942 32388
rect 4884 32379 4942 32385
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 6380 32357 6408 32456
rect 6632 32419 6690 32425
rect 6632 32385 6644 32419
rect 6678 32416 6690 32419
rect 7374 32416 7380 32428
rect 6678 32388 7380 32416
rect 6678 32385 6690 32388
rect 6632 32379 6690 32385
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 8588 32416 8616 32524
rect 9306 32512 9312 32524
rect 9364 32552 9370 32564
rect 9364 32524 11100 32552
rect 9364 32512 9370 32524
rect 8662 32444 8668 32496
rect 8720 32484 8726 32496
rect 8757 32487 8815 32493
rect 8757 32484 8769 32487
rect 8720 32456 8769 32484
rect 8720 32444 8726 32456
rect 8757 32453 8769 32456
rect 8803 32453 8815 32487
rect 8757 32447 8815 32453
rect 8973 32487 9031 32493
rect 8973 32453 8985 32487
rect 9019 32484 9031 32487
rect 9214 32484 9220 32496
rect 9019 32456 9220 32484
rect 9019 32453 9031 32456
rect 8973 32447 9031 32453
rect 8496 32388 8616 32416
rect 8772 32416 8800 32447
rect 9214 32444 9220 32456
rect 9272 32484 9278 32496
rect 11072 32484 11100 32524
rect 11146 32512 11152 32564
rect 11204 32552 11210 32564
rect 11333 32555 11391 32561
rect 11333 32552 11345 32555
rect 11204 32524 11345 32552
rect 11204 32512 11210 32524
rect 11333 32521 11345 32524
rect 11379 32552 11391 32555
rect 11698 32552 11704 32564
rect 11379 32524 11704 32552
rect 11379 32521 11391 32524
rect 11333 32515 11391 32521
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 13630 32512 13636 32564
rect 13688 32512 13694 32564
rect 14093 32555 14151 32561
rect 14093 32521 14105 32555
rect 14139 32552 14151 32555
rect 14918 32552 14924 32564
rect 14139 32524 14924 32552
rect 14139 32521 14151 32524
rect 14093 32515 14151 32521
rect 14918 32512 14924 32524
rect 14976 32512 14982 32564
rect 15197 32555 15255 32561
rect 15197 32521 15209 32555
rect 15243 32521 15255 32555
rect 15197 32515 15255 32521
rect 13265 32487 13323 32493
rect 9272 32456 10548 32484
rect 11072 32456 11836 32484
rect 9272 32444 9278 32456
rect 10318 32416 10324 32428
rect 8772 32388 10324 32416
rect 6365 32351 6423 32357
rect 4019 32320 4108 32348
rect 4540 32320 4660 32348
rect 4019 32317 4031 32320
rect 3973 32311 4031 32317
rect 4080 32224 4108 32320
rect 3510 32172 3516 32224
rect 3568 32172 3574 32224
rect 4062 32172 4068 32224
rect 4120 32172 4126 32224
rect 4632 32212 4660 32320
rect 6365 32317 6377 32351
rect 6411 32317 6423 32351
rect 6365 32311 6423 32317
rect 5902 32240 5908 32292
rect 5960 32280 5966 32292
rect 5997 32283 6055 32289
rect 5997 32280 6009 32283
rect 5960 32252 6009 32280
rect 5960 32240 5966 32252
rect 5997 32249 6009 32252
rect 6043 32249 6055 32283
rect 5997 32243 6055 32249
rect 6270 32240 6276 32292
rect 6328 32240 6334 32292
rect 6288 32212 6316 32240
rect 4632 32184 6316 32212
rect 6380 32212 6408 32311
rect 7834 32308 7840 32360
rect 7892 32348 7898 32360
rect 8389 32351 8447 32357
rect 8389 32348 8401 32351
rect 7892 32320 8401 32348
rect 7892 32308 7898 32320
rect 8389 32317 8401 32320
rect 8435 32317 8447 32351
rect 8389 32311 8447 32317
rect 7745 32283 7803 32289
rect 7745 32249 7757 32283
rect 7791 32280 7803 32283
rect 8202 32280 8208 32292
rect 7791 32252 8208 32280
rect 7791 32249 7803 32252
rect 7745 32243 7803 32249
rect 8202 32240 8208 32252
rect 8260 32240 8266 32292
rect 7006 32212 7012 32224
rect 6380 32184 7012 32212
rect 7006 32172 7012 32184
rect 7064 32172 7070 32224
rect 8496 32212 8524 32388
rect 10318 32376 10324 32388
rect 10376 32376 10382 32428
rect 10520 32360 10548 32456
rect 11808 32425 11836 32456
rect 13265 32453 13277 32487
rect 13311 32484 13323 32487
rect 13538 32484 13544 32496
rect 13311 32456 13544 32484
rect 13311 32453 13323 32456
rect 13265 32447 13323 32453
rect 13538 32444 13544 32456
rect 13596 32484 13602 32496
rect 15212 32484 15240 32515
rect 15562 32512 15568 32564
rect 15620 32512 15626 32564
rect 15654 32512 15660 32564
rect 15712 32512 15718 32564
rect 15930 32512 15936 32564
rect 15988 32512 15994 32564
rect 16298 32552 16304 32564
rect 16132 32524 16304 32552
rect 15948 32484 15976 32512
rect 13596 32456 14872 32484
rect 15212 32456 15976 32484
rect 13596 32444 13602 32456
rect 11793 32419 11851 32425
rect 11793 32385 11805 32419
rect 11839 32416 11851 32419
rect 13906 32416 13912 32428
rect 11839 32388 13912 32416
rect 11839 32385 11851 32388
rect 11793 32379 11851 32385
rect 13906 32376 13912 32388
rect 13964 32376 13970 32428
rect 13998 32376 14004 32428
rect 14056 32376 14062 32428
rect 14274 32376 14280 32428
rect 14332 32376 14338 32428
rect 14366 32376 14372 32428
rect 14424 32376 14430 32428
rect 14458 32376 14464 32428
rect 14516 32376 14522 32428
rect 14550 32376 14556 32428
rect 14608 32425 14614 32428
rect 14608 32419 14637 32425
rect 14625 32385 14637 32419
rect 14608 32379 14637 32385
rect 14608 32376 14614 32379
rect 8570 32308 8576 32360
rect 8628 32348 8634 32360
rect 9217 32351 9275 32357
rect 8628 32320 9016 32348
rect 8628 32308 8634 32320
rect 8901 32215 8959 32221
rect 8901 32212 8913 32215
rect 8496 32184 8913 32212
rect 8901 32181 8913 32184
rect 8947 32181 8959 32215
rect 8988 32212 9016 32320
rect 9217 32317 9229 32351
rect 9263 32348 9275 32351
rect 9306 32348 9312 32360
rect 9263 32320 9312 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 9490 32308 9496 32360
rect 9548 32308 9554 32360
rect 10226 32308 10232 32360
rect 10284 32308 10290 32360
rect 10502 32308 10508 32360
rect 10560 32348 10566 32360
rect 12529 32351 12587 32357
rect 10560 32320 11100 32348
rect 10560 32308 10566 32320
rect 9122 32240 9128 32292
rect 9180 32240 9186 32292
rect 10244 32280 10272 32308
rect 10244 32252 10916 32280
rect 10318 32212 10324 32224
rect 8988 32184 10324 32212
rect 8901 32175 8959 32181
rect 10318 32172 10324 32184
rect 10376 32172 10382 32224
rect 10888 32212 10916 32252
rect 10962 32240 10968 32292
rect 11020 32240 11026 32292
rect 11072 32280 11100 32320
rect 12529 32317 12541 32351
rect 12575 32348 12587 32351
rect 14734 32348 14740 32360
rect 12575 32320 14740 32348
rect 12575 32317 12587 32320
rect 12529 32311 12587 32317
rect 14734 32308 14740 32320
rect 14792 32308 14798 32360
rect 14844 32348 14872 32456
rect 16022 32444 16028 32496
rect 16080 32484 16086 32496
rect 16132 32493 16160 32524
rect 16298 32512 16304 32524
rect 16356 32512 16362 32564
rect 16482 32512 16488 32564
rect 16540 32512 16546 32564
rect 17034 32512 17040 32564
rect 17092 32512 17098 32564
rect 17862 32512 17868 32564
rect 17920 32552 17926 32564
rect 20070 32552 20076 32564
rect 17920 32524 20076 32552
rect 17920 32512 17926 32524
rect 20070 32512 20076 32524
rect 20128 32512 20134 32564
rect 20438 32512 20444 32564
rect 20496 32552 20502 32564
rect 20533 32555 20591 32561
rect 20533 32552 20545 32555
rect 20496 32524 20545 32552
rect 20496 32512 20502 32524
rect 20533 32521 20545 32524
rect 20579 32521 20591 32555
rect 20533 32515 20591 32521
rect 20714 32512 20720 32564
rect 20772 32552 20778 32564
rect 20993 32555 21051 32561
rect 20993 32552 21005 32555
rect 20772 32524 21005 32552
rect 20772 32512 20778 32524
rect 20993 32521 21005 32524
rect 21039 32521 21051 32555
rect 20993 32515 21051 32521
rect 22462 32512 22468 32564
rect 22520 32512 22526 32564
rect 24486 32512 24492 32564
rect 24544 32552 24550 32564
rect 24765 32555 24823 32561
rect 24765 32552 24777 32555
rect 24544 32524 24777 32552
rect 24544 32512 24550 32524
rect 24765 32521 24777 32524
rect 24811 32521 24823 32555
rect 24765 32515 24823 32521
rect 24854 32512 24860 32564
rect 24912 32512 24918 32564
rect 25038 32512 25044 32564
rect 25096 32512 25102 32564
rect 25685 32555 25743 32561
rect 25685 32552 25697 32555
rect 25424 32524 25697 32552
rect 16117 32487 16175 32493
rect 16117 32484 16129 32487
rect 16080 32456 16129 32484
rect 16080 32444 16086 32456
rect 16117 32453 16129 32456
rect 16163 32453 16175 32487
rect 16758 32484 16764 32496
rect 16117 32447 16175 32453
rect 16684 32456 16764 32484
rect 14921 32419 14979 32425
rect 14921 32385 14933 32419
rect 14967 32416 14979 32419
rect 15654 32416 15660 32428
rect 14967 32388 15660 32416
rect 14967 32385 14979 32388
rect 14921 32379 14979 32385
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15930 32416 15936 32428
rect 15764 32388 15936 32416
rect 15764 32348 15792 32388
rect 15930 32376 15936 32388
rect 15988 32416 15994 32428
rect 16684 32425 16712 32456
rect 16758 32444 16764 32456
rect 16816 32444 16822 32496
rect 16301 32419 16359 32425
rect 16301 32416 16313 32419
rect 15988 32388 16313 32416
rect 15988 32376 15994 32388
rect 16301 32385 16313 32388
rect 16347 32385 16359 32419
rect 16301 32379 16359 32385
rect 16669 32419 16727 32425
rect 16669 32385 16681 32419
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 16853 32419 16911 32425
rect 16853 32385 16865 32419
rect 16899 32416 16911 32419
rect 17052 32416 17080 32512
rect 19426 32484 19432 32496
rect 17972 32456 19432 32484
rect 17972 32425 18000 32456
rect 19426 32444 19432 32456
rect 19484 32484 19490 32496
rect 20898 32484 20904 32496
rect 19484 32456 20904 32484
rect 19484 32444 19490 32456
rect 20898 32444 20904 32456
rect 20956 32444 20962 32496
rect 16899 32388 17080 32416
rect 17957 32419 18015 32425
rect 16899 32385 16911 32388
rect 16853 32379 16911 32385
rect 17957 32385 17969 32419
rect 18003 32385 18015 32419
rect 17957 32379 18015 32385
rect 18224 32419 18282 32425
rect 18224 32385 18236 32419
rect 18270 32416 18282 32419
rect 18506 32416 18512 32428
rect 18270 32388 18512 32416
rect 18270 32385 18282 32388
rect 18224 32379 18282 32385
rect 18506 32376 18512 32388
rect 18564 32376 18570 32428
rect 19242 32376 19248 32428
rect 19300 32416 19306 32428
rect 19613 32419 19671 32425
rect 19613 32416 19625 32419
rect 19300 32388 19625 32416
rect 19300 32376 19306 32388
rect 19613 32385 19625 32388
rect 19659 32385 19671 32419
rect 19613 32379 19671 32385
rect 14844 32320 15792 32348
rect 15841 32351 15899 32357
rect 15841 32317 15853 32351
rect 15887 32348 15899 32351
rect 16574 32348 16580 32360
rect 15887 32320 16580 32348
rect 15887 32317 15899 32320
rect 15841 32311 15899 32317
rect 16574 32308 16580 32320
rect 16632 32308 16638 32360
rect 16942 32308 16948 32360
rect 17000 32348 17006 32360
rect 17037 32351 17095 32357
rect 17037 32348 17049 32351
rect 17000 32320 17049 32348
rect 17000 32308 17006 32320
rect 17037 32317 17049 32320
rect 17083 32317 17095 32351
rect 17037 32311 17095 32317
rect 17218 32308 17224 32360
rect 17276 32308 17282 32360
rect 19334 32308 19340 32360
rect 19392 32348 19398 32360
rect 19429 32351 19487 32357
rect 19429 32348 19441 32351
rect 19392 32320 19441 32348
rect 19392 32308 19398 32320
rect 19429 32317 19441 32320
rect 19475 32317 19487 32351
rect 19631 32348 19659 32379
rect 19978 32376 19984 32428
rect 20036 32376 20042 32428
rect 20438 32416 20444 32428
rect 20079 32388 20444 32416
rect 20079 32348 20107 32388
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 20548 32388 20760 32416
rect 20548 32348 20576 32388
rect 19631 32320 20107 32348
rect 20272 32320 20576 32348
rect 19429 32311 19487 32317
rect 15013 32283 15071 32289
rect 11072 32252 13860 32280
rect 12066 32212 12072 32224
rect 10888 32184 12072 32212
rect 12066 32172 12072 32184
rect 12124 32172 12130 32224
rect 12897 32215 12955 32221
rect 12897 32181 12909 32215
rect 12943 32212 12955 32215
rect 13722 32212 13728 32224
rect 12943 32184 13728 32212
rect 12943 32181 12955 32184
rect 12897 32175 12955 32181
rect 13722 32172 13728 32184
rect 13780 32172 13786 32224
rect 13832 32212 13860 32252
rect 15013 32249 15025 32283
rect 15059 32280 15071 32283
rect 17954 32280 17960 32292
rect 15059 32252 17960 32280
rect 15059 32249 15071 32252
rect 15013 32243 15071 32249
rect 17954 32240 17960 32252
rect 18012 32240 18018 32292
rect 20272 32280 20300 32320
rect 20622 32308 20628 32360
rect 20680 32308 20686 32360
rect 20732 32348 20760 32388
rect 20806 32376 20812 32428
rect 20864 32416 20870 32428
rect 22480 32416 22508 32512
rect 22824 32487 22882 32493
rect 22824 32453 22836 32487
rect 22870 32484 22882 32487
rect 25056 32484 25084 32512
rect 22870 32456 25084 32484
rect 22870 32453 22882 32456
rect 22824 32447 22882 32453
rect 25424 32428 25452 32524
rect 25685 32521 25697 32524
rect 25731 32521 25743 32555
rect 25685 32515 25743 32521
rect 26349 32524 26832 32552
rect 26349 32484 26377 32524
rect 25516 32456 26377 32484
rect 25516 32428 25544 32456
rect 26418 32444 26424 32496
rect 26476 32444 26482 32496
rect 20864 32388 22508 32416
rect 20864 32376 20870 32388
rect 23750 32376 23756 32428
rect 23808 32376 23814 32428
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32416 24087 32419
rect 24118 32416 24124 32428
rect 24075 32388 24124 32416
rect 24075 32385 24087 32388
rect 24029 32379 24087 32385
rect 20990 32348 20996 32360
rect 20732 32320 20996 32348
rect 20990 32308 20996 32320
rect 21048 32308 21054 32360
rect 22094 32308 22100 32360
rect 22152 32348 22158 32360
rect 22557 32351 22615 32357
rect 22557 32348 22569 32351
rect 22152 32320 22569 32348
rect 22152 32308 22158 32320
rect 22557 32317 22569 32320
rect 22603 32317 22615 32351
rect 22557 32311 22615 32317
rect 18892 32252 20300 32280
rect 23768 32280 23796 32376
rect 23842 32308 23848 32360
rect 23900 32348 23906 32360
rect 24044 32348 24072 32379
rect 24118 32376 24124 32388
rect 24176 32376 24182 32428
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32416 24271 32419
rect 24259 32388 24532 32416
rect 24259 32385 24271 32388
rect 24213 32379 24271 32385
rect 23900 32320 24072 32348
rect 23900 32308 23906 32320
rect 24302 32308 24308 32360
rect 24360 32308 24366 32360
rect 24397 32351 24455 32357
rect 24397 32317 24409 32351
rect 24443 32317 24455 32351
rect 24504 32348 24532 32388
rect 24578 32376 24584 32428
rect 24636 32376 24642 32428
rect 24854 32376 24860 32428
rect 24912 32376 24918 32428
rect 24946 32376 24952 32428
rect 25004 32416 25010 32428
rect 25225 32419 25283 32425
rect 25225 32416 25237 32419
rect 25004 32388 25237 32416
rect 25004 32376 25010 32388
rect 25225 32385 25237 32388
rect 25271 32385 25283 32419
rect 25225 32379 25283 32385
rect 25406 32376 25412 32428
rect 25464 32376 25470 32428
rect 25498 32376 25504 32428
rect 25556 32376 25562 32428
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32416 25835 32419
rect 25866 32416 25872 32428
rect 25823 32388 25872 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 25866 32376 25872 32388
rect 25924 32376 25930 32428
rect 26050 32376 26056 32428
rect 26108 32376 26114 32428
rect 26234 32376 26240 32428
rect 26292 32376 26298 32428
rect 26329 32419 26387 32425
rect 26329 32385 26341 32419
rect 26375 32416 26387 32419
rect 26436 32416 26464 32444
rect 26804 32425 26832 32524
rect 26878 32512 26884 32564
rect 26936 32552 26942 32564
rect 27157 32555 27215 32561
rect 27157 32552 27169 32555
rect 26936 32524 27169 32552
rect 26936 32512 26942 32524
rect 27157 32521 27169 32524
rect 27203 32521 27215 32555
rect 27157 32515 27215 32521
rect 27338 32512 27344 32564
rect 27396 32552 27402 32564
rect 27709 32555 27767 32561
rect 27709 32552 27721 32555
rect 27396 32524 27721 32552
rect 27396 32512 27402 32524
rect 27709 32521 27721 32524
rect 27755 32521 27767 32555
rect 28258 32552 28264 32564
rect 27709 32515 27767 32521
rect 27816 32524 28264 32552
rect 27816 32484 27844 32524
rect 28258 32512 28264 32524
rect 28316 32512 28322 32564
rect 28718 32512 28724 32564
rect 28776 32552 28782 32564
rect 28813 32555 28871 32561
rect 28813 32552 28825 32555
rect 28776 32524 28825 32552
rect 28776 32512 28782 32524
rect 28813 32521 28825 32524
rect 28859 32521 28871 32555
rect 28813 32515 28871 32521
rect 29454 32512 29460 32564
rect 29512 32512 29518 32564
rect 29638 32512 29644 32564
rect 29696 32512 29702 32564
rect 30006 32512 30012 32564
rect 30064 32552 30070 32564
rect 30742 32552 30748 32564
rect 30064 32524 30748 32552
rect 30064 32512 30070 32524
rect 29273 32487 29331 32493
rect 29273 32484 29285 32487
rect 27169 32456 27844 32484
rect 28460 32456 29285 32484
rect 26375 32388 26464 32416
rect 26605 32419 26663 32425
rect 26375 32385 26387 32388
rect 26329 32379 26387 32385
rect 26605 32385 26617 32419
rect 26651 32385 26663 32419
rect 26605 32379 26663 32385
rect 26789 32419 26847 32425
rect 26789 32385 26801 32419
rect 26835 32385 26847 32419
rect 26789 32379 26847 32385
rect 24872 32348 24900 32376
rect 24504 32320 24900 32348
rect 25041 32351 25099 32357
rect 24397 32311 24455 32317
rect 25041 32317 25053 32351
rect 25087 32317 25099 32351
rect 25041 32311 25099 32317
rect 24118 32280 24124 32292
rect 23768 32252 24124 32280
rect 16390 32212 16396 32224
rect 13832 32184 16396 32212
rect 16390 32172 16396 32184
rect 16448 32172 16454 32224
rect 16666 32172 16672 32224
rect 16724 32212 16730 32224
rect 17865 32215 17923 32221
rect 17865 32212 17877 32215
rect 16724 32184 17877 32212
rect 16724 32172 16730 32184
rect 17865 32181 17877 32184
rect 17911 32181 17923 32215
rect 17865 32175 17923 32181
rect 18598 32172 18604 32224
rect 18656 32212 18662 32224
rect 18892 32212 18920 32252
rect 24118 32240 24124 32252
rect 24176 32280 24182 32292
rect 24412 32280 24440 32311
rect 24176 32252 24440 32280
rect 24176 32240 24182 32252
rect 24670 32240 24676 32292
rect 24728 32280 24734 32292
rect 25056 32280 25084 32311
rect 25130 32308 25136 32360
rect 25188 32308 25194 32360
rect 25317 32351 25375 32357
rect 25317 32317 25329 32351
rect 25363 32317 25375 32351
rect 25424 32348 25452 32376
rect 26620 32348 26648 32379
rect 25424 32320 26648 32348
rect 25317 32311 25375 32317
rect 24728 32252 25084 32280
rect 25332 32280 25360 32311
rect 25332 32252 26464 32280
rect 24728 32240 24734 32252
rect 18656 32184 18920 32212
rect 18656 32172 18662 32184
rect 18966 32172 18972 32224
rect 19024 32212 19030 32224
rect 19337 32215 19395 32221
rect 19337 32212 19349 32215
rect 19024 32184 19349 32212
rect 19024 32172 19030 32184
rect 19337 32181 19349 32184
rect 19383 32181 19395 32215
rect 19337 32175 19395 32181
rect 19797 32215 19855 32221
rect 19797 32181 19809 32215
rect 19843 32212 19855 32215
rect 20070 32212 20076 32224
rect 19843 32184 20076 32212
rect 19843 32181 19855 32184
rect 19797 32175 19855 32181
rect 20070 32172 20076 32184
rect 20128 32172 20134 32224
rect 20346 32172 20352 32224
rect 20404 32212 20410 32224
rect 21266 32212 21272 32224
rect 20404 32184 21272 32212
rect 20404 32172 20410 32184
rect 21266 32172 21272 32184
rect 21324 32172 21330 32224
rect 22002 32172 22008 32224
rect 22060 32172 22066 32224
rect 23934 32172 23940 32224
rect 23992 32172 23998 32224
rect 25222 32172 25228 32224
rect 25280 32212 25286 32224
rect 25501 32215 25559 32221
rect 25501 32212 25513 32215
rect 25280 32184 25513 32212
rect 25280 32172 25286 32184
rect 25501 32181 25513 32184
rect 25547 32181 25559 32215
rect 25501 32175 25559 32181
rect 25590 32172 25596 32224
rect 25648 32212 25654 32224
rect 26326 32212 26332 32224
rect 25648 32184 26332 32212
rect 25648 32172 25654 32184
rect 26326 32172 26332 32184
rect 26384 32172 26390 32224
rect 26436 32212 26464 32252
rect 26510 32240 26516 32292
rect 26568 32240 26574 32292
rect 26605 32283 26663 32289
rect 26605 32249 26617 32283
rect 26651 32249 26663 32283
rect 26804 32280 26832 32379
rect 26878 32376 26884 32428
rect 26936 32416 26942 32428
rect 27169 32425 27197 32456
rect 27154 32419 27212 32425
rect 27154 32416 27166 32419
rect 26936 32388 27166 32416
rect 26936 32376 26942 32388
rect 27154 32385 27166 32388
rect 27200 32385 27212 32419
rect 27154 32379 27212 32385
rect 27246 32376 27252 32428
rect 27304 32416 27310 32428
rect 27617 32419 27675 32425
rect 27617 32416 27629 32419
rect 27304 32388 27629 32416
rect 27304 32376 27310 32388
rect 27617 32385 27629 32388
rect 27663 32385 27675 32419
rect 27617 32379 27675 32385
rect 27798 32376 27804 32428
rect 27856 32416 27862 32428
rect 27893 32419 27951 32425
rect 27893 32416 27905 32419
rect 27856 32388 27905 32416
rect 27856 32376 27862 32388
rect 27893 32385 27905 32388
rect 27939 32385 27951 32419
rect 27893 32379 27951 32385
rect 28166 32376 28172 32428
rect 28224 32376 28230 32428
rect 28350 32376 28356 32428
rect 28408 32376 28414 32428
rect 26970 32308 26976 32360
rect 27028 32348 27034 32360
rect 27338 32348 27344 32360
rect 27028 32320 27344 32348
rect 27028 32308 27034 32320
rect 27338 32308 27344 32320
rect 27396 32308 27402 32360
rect 27522 32308 27528 32360
rect 27580 32348 27586 32360
rect 28460 32348 28488 32456
rect 29273 32453 29285 32456
rect 29319 32453 29331 32487
rect 29472 32484 29500 32512
rect 29472 32456 30144 32484
rect 29273 32447 29331 32453
rect 28629 32419 28687 32425
rect 28629 32385 28641 32419
rect 28675 32416 28687 32419
rect 28718 32416 28724 32428
rect 28675 32388 28724 32416
rect 28675 32385 28687 32388
rect 28629 32379 28687 32385
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32416 28963 32419
rect 28994 32416 29000 32428
rect 28951 32388 29000 32416
rect 28951 32385 28963 32388
rect 28905 32379 28963 32385
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 29089 32419 29147 32425
rect 29089 32385 29101 32419
rect 29135 32385 29147 32419
rect 29089 32379 29147 32385
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32385 29975 32419
rect 29917 32379 29975 32385
rect 27580 32320 28488 32348
rect 28537 32351 28595 32357
rect 27580 32308 27586 32320
rect 28537 32317 28549 32351
rect 28583 32348 28595 32351
rect 28810 32348 28816 32360
rect 28583 32320 28816 32348
rect 28583 32317 28595 32320
rect 28537 32311 28595 32317
rect 28810 32308 28816 32320
rect 28868 32348 28874 32360
rect 29104 32348 29132 32379
rect 28868 32320 29132 32348
rect 28868 32308 28874 32320
rect 26804 32252 27936 32280
rect 26605 32243 26663 32249
rect 26618 32212 26646 32243
rect 26436 32184 26646 32212
rect 26970 32172 26976 32224
rect 27028 32172 27034 32224
rect 27908 32212 27936 32252
rect 27982 32240 27988 32292
rect 28040 32240 28046 32292
rect 28077 32283 28135 32289
rect 28077 32249 28089 32283
rect 28123 32280 28135 32283
rect 29932 32280 29960 32379
rect 30006 32376 30012 32428
rect 30064 32376 30070 32428
rect 30116 32425 30144 32456
rect 30300 32425 30328 32524
rect 30742 32512 30748 32524
rect 30800 32552 30806 32564
rect 32214 32552 32220 32564
rect 30800 32524 32220 32552
rect 30800 32512 30806 32524
rect 32214 32512 32220 32524
rect 32272 32512 32278 32564
rect 30828 32487 30886 32493
rect 30828 32453 30840 32487
rect 30874 32484 30886 32487
rect 33042 32484 33048 32496
rect 30874 32456 33048 32484
rect 30874 32453 30886 32456
rect 30828 32447 30886 32453
rect 33042 32444 33048 32456
rect 33100 32444 33106 32496
rect 30101 32419 30159 32425
rect 30101 32385 30113 32419
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 30285 32419 30343 32425
rect 30285 32385 30297 32419
rect 30331 32385 30343 32419
rect 30285 32379 30343 32385
rect 30374 32376 30380 32428
rect 30432 32416 30438 32428
rect 30561 32419 30619 32425
rect 30561 32416 30573 32419
rect 30432 32388 30573 32416
rect 30432 32376 30438 32388
rect 30561 32385 30573 32388
rect 30607 32385 30619 32419
rect 30561 32379 30619 32385
rect 31386 32376 31392 32428
rect 31444 32416 31450 32428
rect 32125 32419 32183 32425
rect 32125 32416 32137 32419
rect 31444 32388 32137 32416
rect 31444 32376 31450 32388
rect 32125 32385 32137 32388
rect 32171 32385 32183 32419
rect 32125 32379 32183 32385
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 32355 32388 32720 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 30466 32280 30472 32292
rect 28123 32252 28994 32280
rect 29932 32252 30472 32280
rect 28123 32249 28135 32252
rect 28077 32243 28135 32249
rect 28092 32212 28120 32243
rect 27908 32184 28120 32212
rect 28626 32172 28632 32224
rect 28684 32172 28690 32224
rect 28966 32212 28994 32252
rect 30466 32240 30472 32252
rect 30524 32240 30530 32292
rect 29362 32212 29368 32224
rect 28966 32184 29368 32212
rect 29362 32172 29368 32184
rect 29420 32172 29426 32224
rect 30834 32172 30840 32224
rect 30892 32212 30898 32224
rect 31941 32215 31999 32221
rect 31941 32212 31953 32215
rect 30892 32184 31953 32212
rect 30892 32172 30898 32184
rect 31941 32181 31953 32184
rect 31987 32181 31999 32215
rect 31941 32175 31999 32181
rect 32122 32172 32128 32224
rect 32180 32172 32186 32224
rect 32692 32221 32720 32388
rect 32677 32215 32735 32221
rect 32677 32181 32689 32215
rect 32723 32212 32735 32215
rect 32766 32212 32772 32224
rect 32723 32184 32772 32212
rect 32723 32181 32735 32184
rect 32677 32175 32735 32181
rect 32766 32172 32772 32184
rect 32824 32172 32830 32224
rect 1104 32122 43884 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 43884 32122
rect 1104 32048 43884 32070
rect 1854 32008 1860 32020
rect 1688 31980 1860 32008
rect 1688 31881 1716 31980
rect 1854 31968 1860 31980
rect 1912 31968 1918 32020
rect 3510 32008 3516 32020
rect 2746 31980 3516 32008
rect 1673 31875 1731 31881
rect 1673 31841 1685 31875
rect 1719 31841 1731 31875
rect 1673 31835 1731 31841
rect 1940 31807 1998 31813
rect 1940 31773 1952 31807
rect 1986 31804 1998 31807
rect 2746 31804 2774 31980
rect 3510 31968 3516 31980
rect 3568 31968 3574 32020
rect 3789 32011 3847 32017
rect 3789 31977 3801 32011
rect 3835 32008 3847 32011
rect 4706 32008 4712 32020
rect 3835 31980 4712 32008
rect 3835 31977 3847 31980
rect 3789 31971 3847 31977
rect 4706 31968 4712 31980
rect 4764 31968 4770 32020
rect 4801 32011 4859 32017
rect 4801 31977 4813 32011
rect 4847 32008 4859 32011
rect 4890 32008 4896 32020
rect 4847 31980 4896 32008
rect 4847 31977 4859 31980
rect 4801 31971 4859 31977
rect 4890 31968 4896 31980
rect 4948 31968 4954 32020
rect 5350 32008 5356 32020
rect 4992 31980 5356 32008
rect 4992 31940 5020 31980
rect 5350 31968 5356 31980
rect 5408 32008 5414 32020
rect 5905 32011 5963 32017
rect 5905 32008 5917 32011
rect 5408 31980 5917 32008
rect 5408 31968 5414 31980
rect 5905 31977 5917 31980
rect 5951 32008 5963 32011
rect 5951 31980 6500 32008
rect 5951 31977 5963 31980
rect 5905 31971 5963 31977
rect 6365 31943 6423 31949
rect 6365 31940 6377 31943
rect 4356 31912 5020 31940
rect 5276 31912 6377 31940
rect 4356 31884 4384 31912
rect 4338 31832 4344 31884
rect 4396 31832 4402 31884
rect 4890 31832 4896 31884
rect 4948 31872 4954 31884
rect 5276 31881 5304 31912
rect 6365 31909 6377 31912
rect 6411 31909 6423 31943
rect 6472 31940 6500 31980
rect 7374 31968 7380 32020
rect 7432 31968 7438 32020
rect 8570 31968 8576 32020
rect 8628 31968 8634 32020
rect 9306 31968 9312 32020
rect 9364 32008 9370 32020
rect 10321 32011 10379 32017
rect 10321 32008 10333 32011
rect 9364 31980 10333 32008
rect 9364 31968 9370 31980
rect 10321 31977 10333 31980
rect 10367 32008 10379 32011
rect 11790 32008 11796 32020
rect 10367 31980 11796 32008
rect 10367 31977 10379 31980
rect 10321 31971 10379 31977
rect 11790 31968 11796 31980
rect 11848 31968 11854 32020
rect 12250 31968 12256 32020
rect 12308 32008 12314 32020
rect 12308 31980 12756 32008
rect 12308 31968 12314 31980
rect 8588 31940 8616 31968
rect 6472 31912 8616 31940
rect 6365 31903 6423 31909
rect 11606 31900 11612 31952
rect 11664 31940 11670 31952
rect 12728 31940 12756 31980
rect 14182 31968 14188 32020
rect 14240 31968 14246 32020
rect 14274 31968 14280 32020
rect 14332 32008 14338 32020
rect 15381 32011 15439 32017
rect 15381 32008 15393 32011
rect 14332 31980 15393 32008
rect 14332 31968 14338 31980
rect 15381 31977 15393 31980
rect 15427 31977 15439 32011
rect 15381 31971 15439 31977
rect 16574 31968 16580 32020
rect 16632 32008 16638 32020
rect 17865 32011 17923 32017
rect 17865 32008 17877 32011
rect 16632 31980 17877 32008
rect 16632 31968 16638 31980
rect 17865 31977 17877 31980
rect 17911 31977 17923 32011
rect 17865 31971 17923 31977
rect 17954 31968 17960 32020
rect 18012 32008 18018 32020
rect 18012 31980 18276 32008
rect 18012 31968 18018 31980
rect 11664 31912 12296 31940
rect 12728 31912 12848 31940
rect 11664 31900 11670 31912
rect 5261 31875 5319 31881
rect 5261 31872 5273 31875
rect 4948 31844 5273 31872
rect 4948 31832 4954 31844
rect 5261 31841 5273 31844
rect 5307 31841 5319 31875
rect 5261 31835 5319 31841
rect 5350 31832 5356 31884
rect 5408 31832 5414 31884
rect 5442 31832 5448 31884
rect 5500 31872 5506 31884
rect 5500 31844 6592 31872
rect 5500 31832 5506 31844
rect 6089 31807 6147 31813
rect 6089 31804 6101 31807
rect 1986 31776 2774 31804
rect 5920 31776 6101 31804
rect 1986 31773 1998 31776
rect 1940 31767 1998 31773
rect 5920 31748 5948 31776
rect 6089 31773 6101 31776
rect 6135 31773 6147 31807
rect 6089 31767 6147 31773
rect 6362 31764 6368 31816
rect 6420 31764 6426 31816
rect 6564 31813 6592 31844
rect 7006 31832 7012 31884
rect 7064 31872 7070 31884
rect 7064 31844 8984 31872
rect 7064 31832 7070 31844
rect 6549 31807 6607 31813
rect 6549 31773 6561 31807
rect 6595 31773 6607 31807
rect 6549 31767 6607 31773
rect 6822 31764 6828 31816
rect 6880 31764 6886 31816
rect 7558 31764 7564 31816
rect 7616 31804 7622 31816
rect 8018 31804 8024 31816
rect 7616 31776 8024 31804
rect 7616 31764 7622 31776
rect 8018 31764 8024 31776
rect 8076 31764 8082 31816
rect 8113 31807 8171 31813
rect 8113 31773 8125 31807
rect 8159 31804 8171 31807
rect 8202 31804 8208 31816
rect 8159 31776 8208 31804
rect 8159 31773 8171 31776
rect 8113 31767 8171 31773
rect 8202 31764 8208 31776
rect 8260 31764 8266 31816
rect 8956 31813 8984 31844
rect 8941 31807 8999 31813
rect 8941 31773 8953 31807
rect 8987 31804 8999 31807
rect 9582 31804 9588 31816
rect 8987 31776 9588 31804
rect 8987 31773 8999 31776
rect 8941 31767 8999 31773
rect 9582 31764 9588 31776
rect 9640 31764 9646 31816
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31804 10747 31807
rect 10962 31804 10968 31816
rect 10735 31776 10968 31804
rect 10735 31773 10747 31776
rect 10689 31767 10747 31773
rect 10962 31764 10968 31776
rect 11020 31804 11026 31816
rect 11517 31807 11575 31813
rect 11517 31804 11529 31807
rect 11020 31776 11529 31804
rect 11020 31764 11026 31776
rect 11517 31773 11529 31776
rect 11563 31804 11575 31807
rect 11885 31807 11943 31813
rect 11885 31804 11897 31807
rect 11563 31776 11897 31804
rect 11563 31773 11575 31776
rect 11517 31767 11575 31773
rect 11885 31773 11897 31776
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12268 31804 12296 31912
rect 12820 31881 12848 31912
rect 12986 31900 12992 31952
rect 13044 31940 13050 31952
rect 13081 31943 13139 31949
rect 13081 31940 13093 31943
rect 13044 31912 13093 31940
rect 13044 31900 13050 31912
rect 13081 31909 13093 31912
rect 13127 31909 13139 31943
rect 13081 31903 13139 31909
rect 13538 31900 13544 31952
rect 13596 31900 13602 31952
rect 14200 31940 14228 31968
rect 18046 31940 18052 31952
rect 14200 31912 15238 31940
rect 12805 31875 12863 31881
rect 12805 31841 12817 31875
rect 12851 31872 12863 31875
rect 13556 31872 13584 31900
rect 12851 31844 13584 31872
rect 14093 31875 14151 31881
rect 12851 31841 12863 31844
rect 12805 31835 12863 31841
rect 14093 31841 14105 31875
rect 14139 31872 14151 31875
rect 14550 31872 14556 31884
rect 14139 31844 14556 31872
rect 14139 31841 14151 31844
rect 14093 31835 14151 31841
rect 14550 31832 14556 31844
rect 14608 31832 14614 31884
rect 12342 31804 12348 31816
rect 12115 31776 12348 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 15210 31813 15238 31912
rect 17972 31912 18052 31940
rect 15470 31832 15476 31884
rect 15528 31872 15534 31884
rect 15657 31875 15715 31881
rect 15657 31872 15669 31875
rect 15528 31844 15669 31872
rect 15528 31832 15534 31844
rect 15657 31841 15669 31844
rect 15703 31872 15715 31875
rect 16022 31872 16028 31884
rect 15703 31844 16028 31872
rect 15703 31841 15715 31844
rect 15657 31835 15715 31841
rect 16022 31832 16028 31844
rect 16080 31832 16086 31884
rect 14369 31807 14427 31813
rect 14369 31773 14381 31807
rect 14415 31804 14427 31807
rect 15195 31807 15253 31813
rect 14415 31776 14504 31804
rect 14415 31773 14427 31776
rect 14369 31767 14427 31773
rect 3418 31736 3424 31748
rect 3068 31708 3424 31736
rect 3068 31677 3096 31708
rect 3418 31696 3424 31708
rect 3476 31696 3482 31748
rect 4154 31696 4160 31748
rect 4212 31696 4218 31748
rect 5902 31696 5908 31748
rect 5960 31696 5966 31748
rect 8478 31696 8484 31748
rect 8536 31736 8542 31748
rect 9186 31739 9244 31745
rect 9186 31736 9198 31739
rect 8536 31708 9198 31736
rect 8536 31696 8542 31708
rect 9186 31705 9198 31708
rect 9232 31705 9244 31739
rect 9186 31699 9244 31705
rect 14476 31680 14504 31776
rect 15195 31773 15207 31807
rect 15241 31773 15253 31807
rect 15195 31767 15253 31773
rect 15746 31764 15752 31816
rect 15804 31764 15810 31816
rect 16393 31807 16451 31813
rect 16393 31773 16405 31807
rect 16439 31804 16451 31807
rect 17972 31806 18000 31912
rect 18046 31900 18052 31912
rect 18104 31900 18110 31952
rect 18138 31832 18144 31884
rect 18196 31832 18202 31884
rect 18248 31881 18276 31980
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 18877 32011 18935 32017
rect 18877 32008 18889 32011
rect 18564 31980 18889 32008
rect 18564 31968 18570 31980
rect 18877 31977 18889 31980
rect 18923 31977 18935 32011
rect 18877 31971 18935 31977
rect 19058 31968 19064 32020
rect 19116 31968 19122 32020
rect 19610 31968 19616 32020
rect 19668 32008 19674 32020
rect 20254 32008 20260 32020
rect 19668 31980 20260 32008
rect 19668 31968 19674 31980
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 21545 32011 21603 32017
rect 21545 32008 21557 32011
rect 20824 31980 21557 32008
rect 18233 31875 18291 31881
rect 18233 31841 18245 31875
rect 18279 31841 18291 31875
rect 19076 31872 19104 31968
rect 19150 31900 19156 31952
rect 19208 31940 19214 31952
rect 19521 31943 19579 31949
rect 19521 31940 19533 31943
rect 19208 31912 19533 31940
rect 19208 31900 19214 31912
rect 19521 31909 19533 31912
rect 19567 31909 19579 31943
rect 19521 31903 19579 31909
rect 18233 31835 18291 31841
rect 18708 31844 19104 31872
rect 18708 31813 18736 31844
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 19484 31844 19625 31872
rect 19484 31832 19490 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 19613 31835 19671 31841
rect 19886 31813 19892 31816
rect 18049 31807 18107 31813
rect 18049 31806 18061 31807
rect 16439 31776 16804 31804
rect 17972 31778 18061 31806
rect 16439 31773 16451 31776
rect 16393 31767 16451 31773
rect 15013 31739 15071 31745
rect 15013 31705 15025 31739
rect 15059 31736 15071 31739
rect 15059 31708 15139 31736
rect 15059 31705 15071 31708
rect 15013 31699 15071 31705
rect 3053 31671 3111 31677
rect 3053 31637 3065 31671
rect 3099 31637 3111 31671
rect 3053 31631 3111 31637
rect 3513 31671 3571 31677
rect 3513 31637 3525 31671
rect 3559 31668 3571 31671
rect 3878 31668 3884 31680
rect 3559 31640 3884 31668
rect 3559 31637 3571 31640
rect 3513 31631 3571 31637
rect 3878 31628 3884 31640
rect 3936 31628 3942 31680
rect 4249 31671 4307 31677
rect 4249 31637 4261 31671
rect 4295 31668 4307 31671
rect 4982 31668 4988 31680
rect 4295 31640 4988 31668
rect 4295 31637 4307 31640
rect 4249 31631 4307 31637
rect 4982 31628 4988 31640
rect 5040 31628 5046 31680
rect 5166 31628 5172 31680
rect 5224 31668 5230 31680
rect 6273 31671 6331 31677
rect 6273 31668 6285 31671
rect 5224 31640 6285 31668
rect 5224 31628 5230 31640
rect 6273 31637 6285 31640
rect 6319 31637 6331 31671
rect 6273 31631 6331 31637
rect 7466 31628 7472 31680
rect 7524 31668 7530 31680
rect 8297 31671 8355 31677
rect 8297 31668 8309 31671
rect 7524 31640 8309 31668
rect 7524 31628 7530 31640
rect 8297 31637 8309 31640
rect 8343 31637 8355 31671
rect 8297 31631 8355 31637
rect 8754 31628 8760 31680
rect 8812 31668 8818 31680
rect 9490 31668 9496 31680
rect 8812 31640 9496 31668
rect 8812 31628 8818 31640
rect 9490 31628 9496 31640
rect 9548 31628 9554 31680
rect 10042 31628 10048 31680
rect 10100 31668 10106 31680
rect 11241 31671 11299 31677
rect 11241 31668 11253 31671
rect 10100 31640 11253 31668
rect 10100 31628 10106 31640
rect 11241 31637 11253 31640
rect 11287 31637 11299 31671
rect 11241 31631 11299 31637
rect 12066 31628 12072 31680
rect 12124 31668 12130 31680
rect 12253 31671 12311 31677
rect 12253 31668 12265 31671
rect 12124 31640 12265 31668
rect 12124 31628 12130 31640
rect 12253 31637 12265 31640
rect 12299 31637 12311 31671
rect 12253 31631 12311 31637
rect 13538 31628 13544 31680
rect 13596 31628 13602 31680
rect 13722 31628 13728 31680
rect 13780 31668 13786 31680
rect 13909 31671 13967 31677
rect 13909 31668 13921 31671
rect 13780 31640 13921 31668
rect 13780 31628 13786 31640
rect 13909 31637 13921 31640
rect 13955 31668 13967 31671
rect 14182 31668 14188 31680
rect 13955 31640 14188 31668
rect 13955 31637 13967 31640
rect 13909 31631 13967 31637
rect 14182 31628 14188 31640
rect 14240 31628 14246 31680
rect 14458 31628 14464 31680
rect 14516 31628 14522 31680
rect 15111 31668 15139 31708
rect 15470 31696 15476 31748
rect 15528 31736 15534 31748
rect 15764 31736 15792 31764
rect 16408 31736 16436 31767
rect 16776 31748 16804 31776
rect 18049 31773 18061 31778
rect 18095 31773 18107 31807
rect 18049 31767 18107 31773
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31773 18383 31807
rect 18325 31767 18383 31773
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18693 31807 18751 31813
rect 18555 31776 18644 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 16666 31745 16672 31748
rect 15528 31708 16436 31736
rect 15528 31696 15534 31708
rect 16660 31699 16672 31745
rect 16666 31696 16672 31699
rect 16724 31696 16730 31748
rect 16758 31696 16764 31748
rect 16816 31696 16822 31748
rect 17586 31696 17592 31748
rect 17644 31736 17650 31748
rect 18340 31736 18368 31767
rect 17644 31708 18368 31736
rect 18616 31736 18644 31776
rect 18693 31773 18705 31807
rect 18739 31773 18751 31807
rect 18693 31767 18751 31773
rect 19337 31807 19395 31813
rect 19337 31773 19349 31807
rect 19383 31804 19395 31807
rect 19383 31776 19847 31804
rect 19383 31773 19395 31776
rect 19337 31767 19395 31773
rect 19819 31736 19847 31776
rect 19880 31767 19892 31813
rect 19886 31764 19892 31767
rect 19944 31764 19950 31816
rect 20824 31804 20852 31980
rect 21545 31977 21557 31980
rect 21591 32008 21603 32011
rect 24670 32008 24676 32020
rect 21591 31980 24676 32008
rect 21591 31977 21603 31980
rect 21545 31971 21603 31977
rect 24670 31968 24676 31980
rect 24728 31968 24734 32020
rect 25501 32011 25559 32017
rect 25501 31977 25513 32011
rect 25547 31977 25559 32011
rect 25501 31971 25559 31977
rect 25685 32011 25743 32017
rect 25685 31977 25697 32011
rect 25731 32008 25743 32011
rect 26234 32008 26240 32020
rect 25731 31980 26240 32008
rect 25731 31977 25743 31980
rect 25685 31971 25743 31977
rect 20990 31900 20996 31952
rect 21048 31900 21054 31952
rect 23477 31943 23535 31949
rect 23477 31909 23489 31943
rect 23523 31909 23535 31943
rect 23477 31903 23535 31909
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 22094 31872 22100 31884
rect 20956 31844 22100 31872
rect 20956 31832 20962 31844
rect 22094 31832 22100 31844
rect 22152 31832 22158 31884
rect 21085 31807 21143 31813
rect 21085 31804 21097 31807
rect 20824 31776 21097 31804
rect 21085 31773 21097 31776
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 21453 31807 21511 31813
rect 21453 31773 21465 31807
rect 21499 31773 21511 31807
rect 21637 31807 21695 31813
rect 21637 31804 21649 31807
rect 21453 31767 21511 31773
rect 21560 31776 21649 31804
rect 20254 31736 20260 31748
rect 18616 31708 19334 31736
rect 19819 31708 20260 31736
rect 17644 31696 17650 31708
rect 15562 31668 15568 31680
rect 15111 31640 15568 31668
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 15746 31628 15752 31680
rect 15804 31668 15810 31680
rect 16301 31671 16359 31677
rect 16301 31668 16313 31671
rect 15804 31640 16313 31668
rect 15804 31628 15810 31640
rect 16301 31637 16313 31640
rect 16347 31637 16359 31671
rect 16301 31631 16359 31637
rect 16390 31628 16396 31680
rect 16448 31668 16454 31680
rect 17773 31671 17831 31677
rect 17773 31668 17785 31671
rect 16448 31640 17785 31668
rect 16448 31628 16454 31640
rect 17773 31637 17785 31640
rect 17819 31637 17831 31671
rect 19306 31668 19334 31708
rect 20254 31696 20260 31708
rect 20312 31696 20318 31748
rect 20530 31696 20536 31748
rect 20588 31736 20594 31748
rect 21192 31736 21220 31767
rect 20588 31708 21220 31736
rect 20588 31696 20594 31708
rect 21266 31696 21272 31748
rect 21324 31736 21330 31748
rect 21361 31739 21419 31745
rect 21361 31736 21373 31739
rect 21324 31708 21373 31736
rect 21324 31696 21330 31708
rect 21361 31705 21373 31708
rect 21407 31705 21419 31739
rect 21361 31699 21419 31705
rect 21468 31680 21496 31767
rect 21560 31680 21588 31776
rect 21637 31773 21649 31776
rect 21683 31773 21695 31807
rect 21637 31767 21695 31773
rect 22364 31807 22422 31813
rect 22364 31773 22376 31807
rect 22410 31804 22422 31807
rect 22410 31776 23244 31804
rect 22410 31773 22422 31776
rect 22364 31767 22422 31773
rect 23216 31736 23244 31776
rect 23290 31764 23296 31816
rect 23348 31804 23354 31816
rect 23492 31804 23520 31903
rect 25130 31900 25136 31952
rect 25188 31900 25194 31952
rect 25516 31940 25544 31971
rect 26234 31968 26240 31980
rect 26292 31968 26298 32020
rect 26786 31968 26792 32020
rect 26844 32008 26850 32020
rect 26844 31980 30512 32008
rect 26844 31968 26850 31980
rect 26326 31940 26332 31952
rect 25516 31912 26332 31940
rect 26326 31900 26332 31912
rect 26384 31940 26390 31952
rect 27798 31940 27804 31952
rect 26384 31912 26740 31940
rect 26384 31900 26390 31912
rect 23842 31832 23848 31884
rect 23900 31872 23906 31884
rect 24581 31875 24639 31881
rect 24581 31872 24593 31875
rect 23900 31844 24593 31872
rect 23900 31832 23906 31844
rect 24581 31841 24593 31844
rect 24627 31841 24639 31875
rect 24581 31835 24639 31841
rect 25148 31844 25820 31872
rect 23569 31807 23627 31813
rect 23569 31804 23581 31807
rect 23348 31776 23581 31804
rect 23348 31764 23354 31776
rect 23569 31773 23581 31776
rect 23615 31773 23627 31807
rect 23569 31767 23627 31773
rect 24394 31764 24400 31816
rect 24452 31764 24458 31816
rect 24762 31764 24768 31816
rect 24820 31764 24826 31816
rect 25148 31813 25176 31844
rect 25792 31816 25820 31844
rect 26234 31832 26240 31884
rect 26292 31872 26298 31884
rect 26513 31875 26571 31881
rect 26513 31872 26525 31875
rect 26292 31844 26525 31872
rect 26292 31832 26298 31844
rect 26513 31841 26525 31844
rect 26559 31841 26571 31875
rect 26513 31835 26571 31841
rect 25133 31807 25191 31813
rect 25133 31773 25145 31807
rect 25179 31773 25191 31807
rect 25133 31767 25191 31773
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 25317 31807 25375 31813
rect 25317 31804 25329 31807
rect 25280 31776 25329 31804
rect 25280 31764 25286 31776
rect 25317 31773 25329 31776
rect 25363 31804 25375 31807
rect 25409 31807 25467 31813
rect 25409 31804 25421 31807
rect 25363 31776 25421 31804
rect 25363 31773 25375 31776
rect 25317 31767 25375 31773
rect 25409 31773 25421 31776
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 25774 31764 25780 31816
rect 25832 31764 25838 31816
rect 25866 31764 25872 31816
rect 25924 31804 25930 31816
rect 26053 31807 26111 31813
rect 26053 31804 26065 31807
rect 25924 31776 26065 31804
rect 25924 31764 25930 31776
rect 26053 31773 26065 31776
rect 26099 31773 26111 31807
rect 26053 31767 26111 31773
rect 26142 31764 26148 31816
rect 26200 31764 26206 31816
rect 26712 31813 26740 31912
rect 26804 31912 27804 31940
rect 26804 31816 26832 31912
rect 27798 31900 27804 31912
rect 27856 31900 27862 31952
rect 27982 31900 27988 31952
rect 28040 31940 28046 31952
rect 28353 31943 28411 31949
rect 28353 31940 28365 31943
rect 28040 31912 28365 31940
rect 28040 31900 28046 31912
rect 28353 31909 28365 31912
rect 28399 31909 28411 31943
rect 30098 31940 30104 31952
rect 28353 31903 28411 31909
rect 28644 31912 30104 31940
rect 28644 31884 28672 31912
rect 30098 31900 30104 31912
rect 30156 31900 30162 31952
rect 26878 31832 26884 31884
rect 26936 31832 26942 31884
rect 26973 31875 27031 31881
rect 26973 31841 26985 31875
rect 27019 31872 27031 31875
rect 27338 31872 27344 31884
rect 27019 31844 27344 31872
rect 27019 31841 27031 31844
rect 26973 31835 27031 31841
rect 27338 31832 27344 31844
rect 27396 31872 27402 31884
rect 28626 31872 28632 31884
rect 27396 31844 28632 31872
rect 27396 31832 27402 31844
rect 28626 31832 28632 31844
rect 28684 31832 28690 31884
rect 29086 31832 29092 31884
rect 29144 31872 29150 31884
rect 29144 31844 30328 31872
rect 29144 31832 29150 31844
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31773 26387 31807
rect 26329 31767 26387 31773
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31773 26479 31807
rect 26421 31767 26479 31773
rect 26697 31807 26755 31813
rect 26697 31773 26709 31807
rect 26743 31773 26755 31807
rect 26697 31767 26755 31773
rect 23658 31736 23664 31748
rect 23216 31708 23664 31736
rect 23658 31696 23664 31708
rect 23716 31696 23722 31748
rect 19518 31668 19524 31680
rect 19306 31640 19524 31668
rect 17773 31631 17831 31637
rect 19518 31628 19524 31640
rect 19576 31628 19582 31680
rect 21082 31628 21088 31680
rect 21140 31628 21146 31680
rect 21450 31628 21456 31680
rect 21508 31628 21514 31680
rect 21542 31628 21548 31680
rect 21600 31628 21606 31680
rect 21910 31628 21916 31680
rect 21968 31628 21974 31680
rect 23474 31628 23480 31680
rect 23532 31668 23538 31680
rect 24213 31671 24271 31677
rect 24213 31668 24225 31671
rect 23532 31640 24225 31668
rect 23532 31628 23538 31640
rect 24213 31637 24225 31640
rect 24259 31637 24271 31671
rect 24412 31668 24440 31764
rect 24780 31736 24808 31764
rect 25967 31739 26025 31745
rect 24780 31708 25912 31736
rect 25590 31668 25596 31680
rect 24412 31640 25596 31668
rect 24213 31631 24271 31637
rect 25590 31628 25596 31640
rect 25648 31628 25654 31680
rect 25884 31668 25912 31708
rect 25967 31705 25979 31739
rect 26013 31736 26025 31739
rect 26160 31736 26188 31764
rect 26013 31708 26188 31736
rect 26013 31705 26025 31708
rect 25967 31699 26025 31705
rect 26145 31671 26203 31677
rect 26145 31668 26157 31671
rect 25884 31640 26157 31668
rect 26145 31637 26157 31640
rect 26191 31637 26203 31671
rect 26344 31668 26372 31767
rect 26436 31736 26464 31767
rect 26786 31764 26792 31816
rect 26844 31764 26850 31816
rect 27062 31764 27068 31816
rect 27120 31764 27126 31816
rect 27157 31807 27215 31813
rect 27157 31773 27169 31807
rect 27203 31804 27215 31807
rect 27203 31776 27292 31804
rect 27203 31773 27215 31776
rect 27157 31767 27215 31773
rect 27080 31736 27108 31764
rect 27264 31748 27292 31776
rect 26436 31708 27108 31736
rect 27246 31696 27252 31748
rect 27304 31696 27310 31748
rect 26970 31668 26976 31680
rect 26344 31640 26976 31668
rect 26145 31631 26203 31637
rect 26970 31628 26976 31640
rect 27028 31628 27034 31680
rect 27062 31628 27068 31680
rect 27120 31668 27126 31680
rect 27356 31668 27384 31832
rect 27614 31764 27620 31816
rect 27672 31804 27678 31816
rect 28074 31804 28080 31816
rect 27672 31776 28080 31804
rect 27672 31764 27678 31776
rect 28074 31764 28080 31776
rect 28132 31804 28138 31816
rect 28169 31807 28227 31813
rect 28169 31804 28181 31807
rect 28132 31776 28181 31804
rect 28132 31764 28138 31776
rect 28169 31773 28181 31776
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 28810 31764 28816 31816
rect 28868 31764 28874 31816
rect 28902 31764 28908 31816
rect 28960 31764 28966 31816
rect 29546 31764 29552 31816
rect 29604 31804 29610 31816
rect 30300 31813 30328 31844
rect 30484 31813 30512 31980
rect 31386 31968 31392 32020
rect 31444 31968 31450 32020
rect 33042 31968 33048 32020
rect 33100 31968 33106 32020
rect 31404 31940 31432 31968
rect 30944 31912 31432 31940
rect 30834 31832 30840 31884
rect 30892 31832 30898 31884
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29604 31776 29745 31804
rect 29604 31764 29610 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 30101 31807 30159 31813
rect 30101 31773 30113 31807
rect 30147 31773 30159 31807
rect 30101 31767 30159 31773
rect 30285 31807 30343 31813
rect 30285 31773 30297 31807
rect 30331 31773 30343 31807
rect 30285 31767 30343 31773
rect 30373 31807 30431 31813
rect 30373 31773 30385 31807
rect 30419 31773 30431 31807
rect 30373 31767 30431 31773
rect 30469 31807 30527 31813
rect 30469 31773 30481 31807
rect 30515 31773 30527 31807
rect 30944 31804 30972 31912
rect 31018 31832 31024 31884
rect 31076 31872 31082 31884
rect 31076 31844 31524 31872
rect 31076 31832 31082 31844
rect 31496 31813 31524 31844
rect 32214 31832 32220 31884
rect 32272 31872 32278 31884
rect 32677 31875 32735 31881
rect 32677 31872 32689 31875
rect 32272 31844 32689 31872
rect 32272 31832 32278 31844
rect 32677 31841 32689 31844
rect 32723 31841 32735 31875
rect 32677 31835 32735 31841
rect 30469 31767 30527 31773
rect 30576 31776 30972 31804
rect 31481 31807 31539 31813
rect 27706 31696 27712 31748
rect 27764 31736 27770 31748
rect 27985 31739 28043 31745
rect 27985 31736 27997 31739
rect 27764 31708 27997 31736
rect 27764 31696 27770 31708
rect 27985 31705 27997 31708
rect 28031 31736 28043 31739
rect 28031 31708 29408 31736
rect 28031 31705 28043 31708
rect 27985 31699 28043 31705
rect 29380 31680 29408 31708
rect 27120 31640 27384 31668
rect 27120 31628 27126 31640
rect 28166 31628 28172 31680
rect 28224 31668 28230 31680
rect 28813 31671 28871 31677
rect 28813 31668 28825 31671
rect 28224 31640 28825 31668
rect 28224 31628 28230 31640
rect 28813 31637 28825 31640
rect 28859 31668 28871 31671
rect 29086 31668 29092 31680
rect 28859 31640 29092 31668
rect 28859 31637 28871 31640
rect 28813 31631 28871 31637
rect 29086 31628 29092 31640
rect 29144 31628 29150 31680
rect 29362 31628 29368 31680
rect 29420 31628 29426 31680
rect 30116 31668 30144 31767
rect 30392 31736 30420 31767
rect 30576 31736 30604 31776
rect 31481 31773 31493 31807
rect 31527 31773 31539 31807
rect 31481 31767 31539 31773
rect 32398 31764 32404 31816
rect 32456 31764 32462 31816
rect 32861 31807 32919 31813
rect 32861 31773 32873 31807
rect 32907 31773 32919 31807
rect 32861 31767 32919 31773
rect 32876 31736 32904 31767
rect 30392 31708 30604 31736
rect 30668 31708 32904 31736
rect 30374 31668 30380 31680
rect 30116 31640 30380 31668
rect 30374 31628 30380 31640
rect 30432 31628 30438 31680
rect 30668 31677 30696 31708
rect 30653 31671 30711 31677
rect 30653 31637 30665 31671
rect 30699 31637 30711 31671
rect 30653 31631 30711 31637
rect 32122 31628 32128 31680
rect 32180 31628 32186 31680
rect 32214 31628 32220 31680
rect 32272 31668 32278 31680
rect 32585 31671 32643 31677
rect 32585 31668 32597 31671
rect 32272 31640 32597 31668
rect 32272 31628 32278 31640
rect 32585 31637 32597 31640
rect 32631 31637 32643 31671
rect 32585 31631 32643 31637
rect 1104 31578 43884 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 43884 31578
rect 1104 31504 43884 31526
rect 2958 31424 2964 31476
rect 3016 31464 3022 31476
rect 3697 31467 3755 31473
rect 3697 31464 3709 31467
rect 3016 31436 3709 31464
rect 3016 31424 3022 31436
rect 3697 31433 3709 31436
rect 3743 31433 3755 31467
rect 3697 31427 3755 31433
rect 6822 31424 6828 31476
rect 6880 31424 6886 31476
rect 7576 31436 7880 31464
rect 7576 31408 7604 31436
rect 3142 31356 3148 31408
rect 3200 31396 3206 31408
rect 5442 31396 5448 31408
rect 3200 31368 5448 31396
rect 3200 31356 3206 31368
rect 5442 31356 5448 31368
rect 5500 31356 5506 31408
rect 6181 31399 6239 31405
rect 6181 31365 6193 31399
rect 6227 31396 6239 31399
rect 6549 31399 6607 31405
rect 6549 31396 6561 31399
rect 6227 31368 6561 31396
rect 6227 31365 6239 31368
rect 6181 31359 6239 31365
rect 6549 31365 6561 31368
rect 6595 31396 6607 31399
rect 6914 31396 6920 31408
rect 6595 31368 6920 31396
rect 6595 31365 6607 31368
rect 6549 31359 6607 31365
rect 6914 31356 6920 31368
rect 6972 31396 6978 31408
rect 7377 31399 7435 31405
rect 7377 31396 7389 31399
rect 6972 31368 7389 31396
rect 6972 31356 6978 31368
rect 7377 31365 7389 31368
rect 7423 31396 7435 31399
rect 7558 31396 7564 31408
rect 7423 31368 7564 31396
rect 7423 31365 7435 31368
rect 7377 31359 7435 31365
rect 7558 31356 7564 31368
rect 7616 31356 7622 31408
rect 7742 31356 7748 31408
rect 7800 31356 7806 31408
rect 1946 31288 1952 31340
rect 2004 31288 2010 31340
rect 2216 31331 2274 31337
rect 2216 31297 2228 31331
rect 2262 31328 2274 31331
rect 2498 31328 2504 31340
rect 2262 31300 2504 31328
rect 2262 31297 2274 31300
rect 2216 31291 2274 31297
rect 2498 31288 2504 31300
rect 2556 31288 2562 31340
rect 3878 31288 3884 31340
rect 3936 31328 3942 31340
rect 4065 31331 4123 31337
rect 4065 31328 4077 31331
rect 3936 31300 4077 31328
rect 3936 31288 3942 31300
rect 4065 31297 4077 31300
rect 4111 31297 4123 31331
rect 4065 31291 4123 31297
rect 4890 31288 4896 31340
rect 4948 31288 4954 31340
rect 4982 31288 4988 31340
rect 5040 31288 5046 31340
rect 5077 31331 5135 31337
rect 5077 31297 5089 31331
rect 5123 31297 5135 31331
rect 5077 31291 5135 31297
rect 5273 31331 5331 31337
rect 5273 31297 5285 31331
rect 5319 31297 5331 31331
rect 5273 31291 5331 31297
rect 6365 31331 6423 31337
rect 6365 31297 6377 31331
rect 6411 31328 6423 31331
rect 6454 31328 6460 31340
rect 6411 31300 6460 31328
rect 6411 31297 6423 31300
rect 6365 31291 6423 31297
rect 4157 31263 4215 31269
rect 4157 31229 4169 31263
rect 4203 31229 4215 31263
rect 4157 31223 4215 31229
rect 4062 31152 4068 31204
rect 4120 31192 4126 31204
rect 4172 31192 4200 31223
rect 4338 31220 4344 31272
rect 4396 31260 4402 31272
rect 4798 31260 4804 31272
rect 4396 31232 4804 31260
rect 4396 31220 4402 31232
rect 4798 31220 4804 31232
rect 4856 31220 4862 31272
rect 4120 31164 4200 31192
rect 5092 31192 5120 31291
rect 5276 31260 5304 31291
rect 6454 31288 6460 31300
rect 6512 31288 6518 31340
rect 7098 31288 7104 31340
rect 7156 31288 7162 31340
rect 7653 31331 7711 31337
rect 7653 31297 7665 31331
rect 7699 31328 7711 31331
rect 7760 31328 7788 31356
rect 7852 31337 7880 31436
rect 8478 31424 8484 31476
rect 8536 31424 8542 31476
rect 10134 31424 10140 31476
rect 10192 31464 10198 31476
rect 11514 31464 11520 31476
rect 10192 31436 11520 31464
rect 10192 31424 10198 31436
rect 11514 31424 11520 31436
rect 11572 31424 11578 31476
rect 13538 31424 13544 31476
rect 13596 31464 13602 31476
rect 17037 31467 17095 31473
rect 13596 31436 15608 31464
rect 13596 31424 13602 31436
rect 8110 31356 8116 31408
rect 8168 31396 8174 31408
rect 9033 31399 9091 31405
rect 9033 31396 9045 31399
rect 8168 31368 9045 31396
rect 8168 31356 8174 31368
rect 9033 31365 9045 31368
rect 9079 31365 9091 31399
rect 15470 31396 15476 31408
rect 9033 31359 9091 31365
rect 11532 31368 15476 31396
rect 7699 31300 7788 31328
rect 7837 31331 7895 31337
rect 7699 31297 7711 31300
rect 7653 31291 7711 31297
rect 7837 31297 7849 31331
rect 7883 31297 7895 31331
rect 7837 31291 7895 31297
rect 7929 31331 7987 31337
rect 7929 31297 7941 31331
rect 7975 31297 7987 31331
rect 7929 31291 7987 31297
rect 5534 31260 5540 31272
rect 5276 31232 5540 31260
rect 5534 31220 5540 31232
rect 5592 31220 5598 31272
rect 6733 31263 6791 31269
rect 6733 31229 6745 31263
rect 6779 31260 6791 31263
rect 7009 31263 7067 31269
rect 7009 31260 7021 31263
rect 6779 31232 7021 31260
rect 6779 31229 6791 31232
rect 6733 31223 6791 31229
rect 7009 31229 7021 31232
rect 7055 31229 7067 31263
rect 7009 31223 7067 31229
rect 7466 31220 7472 31272
rect 7524 31220 7530 31272
rect 7745 31263 7803 31269
rect 7745 31229 7757 31263
rect 7791 31260 7803 31263
rect 7944 31260 7972 31291
rect 8202 31288 8208 31340
rect 8260 31288 8266 31340
rect 8297 31331 8355 31337
rect 8297 31297 8309 31331
rect 8343 31328 8355 31331
rect 8754 31328 8760 31340
rect 8343 31300 8760 31328
rect 8343 31297 8355 31300
rect 8297 31291 8355 31297
rect 8754 31288 8760 31300
rect 8812 31288 8818 31340
rect 8849 31331 8907 31337
rect 8849 31297 8861 31331
rect 8895 31297 8907 31331
rect 8849 31291 8907 31297
rect 7791 31232 7972 31260
rect 7791 31229 7803 31232
rect 7745 31223 7803 31229
rect 8662 31192 8668 31204
rect 5092 31164 8668 31192
rect 4120 31152 4126 31164
rect 8662 31152 8668 31164
rect 8720 31192 8726 31204
rect 8864 31192 8892 31291
rect 8938 31288 8944 31340
rect 8996 31288 9002 31340
rect 9582 31288 9588 31340
rect 9640 31288 9646 31340
rect 11532 31337 11560 31368
rect 11517 31331 11575 31337
rect 11517 31297 11529 31331
rect 11563 31297 11575 31331
rect 11517 31291 11575 31297
rect 11606 31288 11612 31340
rect 11664 31328 11670 31340
rect 13188 31337 13216 31368
rect 11773 31331 11831 31337
rect 11773 31328 11785 31331
rect 11664 31300 11785 31328
rect 11664 31288 11670 31300
rect 11773 31297 11785 31300
rect 11819 31297 11831 31331
rect 11773 31291 11831 31297
rect 13173 31331 13231 31337
rect 13173 31297 13185 31331
rect 13219 31297 13231 31331
rect 13173 31291 13231 31297
rect 13440 31331 13498 31337
rect 13440 31297 13452 31331
rect 13486 31328 13498 31331
rect 13722 31328 13728 31340
rect 13486 31300 13728 31328
rect 13486 31297 13498 31300
rect 13440 31291 13498 31297
rect 13722 31288 13728 31300
rect 13780 31288 13786 31340
rect 15028 31337 15056 31368
rect 15470 31356 15476 31368
rect 15528 31356 15534 31408
rect 15013 31331 15071 31337
rect 15013 31297 15025 31331
rect 15059 31297 15071 31331
rect 15269 31331 15327 31337
rect 15269 31328 15281 31331
rect 15013 31291 15071 31297
rect 15120 31300 15281 31328
rect 9306 31220 9312 31272
rect 9364 31220 9370 31272
rect 9858 31220 9864 31272
rect 9916 31220 9922 31272
rect 14274 31220 14280 31272
rect 14332 31260 14338 31272
rect 15120 31260 15148 31300
rect 15269 31297 15281 31300
rect 15315 31297 15327 31331
rect 15580 31328 15608 31436
rect 17037 31433 17049 31467
rect 17083 31464 17095 31467
rect 17218 31464 17224 31476
rect 17083 31436 17224 31464
rect 17083 31433 17095 31436
rect 17037 31427 17095 31433
rect 17218 31424 17224 31436
rect 17276 31424 17282 31476
rect 17862 31424 17868 31476
rect 17920 31424 17926 31476
rect 18414 31424 18420 31476
rect 18472 31424 18478 31476
rect 18598 31424 18604 31476
rect 18656 31464 18662 31476
rect 19242 31464 19248 31476
rect 18656 31436 18736 31464
rect 18656 31424 18662 31436
rect 15654 31356 15660 31408
rect 15712 31396 15718 31408
rect 18322 31396 18328 31408
rect 15712 31368 17908 31396
rect 15712 31356 15718 31368
rect 16776 31337 16804 31368
rect 17880 31340 17908 31368
rect 17972 31368 18328 31396
rect 16761 31331 16819 31337
rect 15580 31300 16712 31328
rect 15269 31291 15327 31297
rect 14332 31232 15148 31260
rect 14332 31220 14338 31232
rect 16022 31220 16028 31272
rect 16080 31260 16086 31272
rect 16390 31260 16396 31272
rect 16080 31232 16396 31260
rect 16080 31220 16086 31232
rect 16390 31220 16396 31232
rect 16448 31220 16454 31272
rect 16684 31260 16712 31300
rect 16761 31297 16773 31331
rect 16807 31297 16819 31331
rect 16761 31291 16819 31297
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 16868 31260 16896 31291
rect 17678 31288 17684 31340
rect 17736 31288 17742 31340
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 17972 31337 18000 31368
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 18708 31405 18736 31436
rect 18938 31436 19248 31464
rect 18693 31399 18751 31405
rect 18693 31365 18705 31399
rect 18739 31365 18751 31399
rect 18693 31359 18751 31365
rect 18782 31356 18788 31408
rect 18840 31356 18846 31408
rect 18938 31405 18966 31436
rect 19242 31424 19248 31436
rect 19300 31464 19306 31476
rect 19417 31464 19423 31476
rect 19300 31436 19423 31464
rect 19300 31424 19306 31436
rect 19417 31424 19423 31436
rect 19475 31424 19481 31476
rect 19705 31467 19763 31473
rect 19705 31433 19717 31467
rect 19751 31464 19763 31467
rect 19978 31464 19984 31476
rect 19751 31436 19984 31464
rect 19751 31433 19763 31436
rect 19705 31427 19763 31433
rect 19978 31424 19984 31436
rect 20036 31424 20042 31476
rect 20530 31424 20536 31476
rect 20588 31464 20594 31476
rect 23474 31464 23480 31476
rect 20588 31436 23480 31464
rect 20588 31424 20594 31436
rect 18923 31399 18981 31405
rect 18923 31365 18935 31399
rect 18969 31365 18981 31399
rect 21082 31396 21088 31408
rect 18923 31359 18981 31365
rect 19076 31368 21088 31396
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31297 18015 31331
rect 17957 31291 18015 31297
rect 18141 31331 18199 31337
rect 18141 31297 18153 31331
rect 18187 31328 18199 31331
rect 18506 31328 18512 31340
rect 18187 31300 18512 31328
rect 18187 31297 18199 31300
rect 18141 31291 18199 31297
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18601 31331 18659 31337
rect 18601 31297 18613 31331
rect 18647 31328 18659 31331
rect 19076 31328 19104 31368
rect 18647 31300 19104 31328
rect 18647 31297 18659 31300
rect 18601 31291 18659 31297
rect 19150 31288 19156 31340
rect 19208 31288 19214 31340
rect 19337 31331 19395 31337
rect 19337 31297 19349 31331
rect 19383 31297 19395 31331
rect 19337 31291 19395 31297
rect 17218 31260 17224 31272
rect 16684 31232 17224 31260
rect 17218 31220 17224 31232
rect 17276 31220 17282 31272
rect 17589 31263 17647 31269
rect 17589 31260 17601 31263
rect 17328 31232 17601 31260
rect 17328 31192 17356 31232
rect 17589 31229 17601 31232
rect 17635 31260 17647 31263
rect 18046 31260 18052 31272
rect 17635 31232 18052 31260
rect 17635 31229 17647 31232
rect 17589 31223 17647 31229
rect 18046 31220 18052 31232
rect 18104 31220 18110 31272
rect 19058 31220 19064 31272
rect 19116 31220 19122 31272
rect 19352 31260 19380 31291
rect 19702 31288 19708 31340
rect 19760 31328 19766 31340
rect 19889 31331 19947 31337
rect 19889 31328 19901 31331
rect 19760 31300 19901 31328
rect 19760 31288 19766 31300
rect 19889 31297 19901 31300
rect 19935 31328 19947 31331
rect 19978 31328 19984 31340
rect 19935 31300 19984 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 19978 31288 19984 31300
rect 20036 31288 20042 31340
rect 20070 31288 20076 31340
rect 20128 31288 20134 31340
rect 20180 31337 20208 31368
rect 21082 31356 21088 31368
rect 21140 31356 21146 31408
rect 21174 31356 21180 31408
rect 21232 31396 21238 31408
rect 22020 31405 22048 31436
rect 23474 31424 23480 31436
rect 23532 31424 23538 31476
rect 23658 31424 23664 31476
rect 23716 31424 23722 31476
rect 24394 31424 24400 31476
rect 24452 31424 24458 31476
rect 24486 31424 24492 31476
rect 24544 31424 24550 31476
rect 24578 31424 24584 31476
rect 24636 31424 24642 31476
rect 25866 31464 25872 31476
rect 25424 31436 25872 31464
rect 22005 31399 22063 31405
rect 21232 31368 21956 31396
rect 21232 31356 21238 31368
rect 20165 31331 20223 31337
rect 20165 31297 20177 31331
rect 20211 31297 20223 31331
rect 20165 31291 20223 31297
rect 20349 31331 20407 31337
rect 20349 31297 20361 31331
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20533 31331 20591 31337
rect 20622 31331 20628 31340
rect 20533 31297 20545 31331
rect 20579 31303 20628 31331
rect 20579 31297 20591 31303
rect 20533 31291 20591 31297
rect 19168 31232 19380 31260
rect 20364 31260 20392 31291
rect 20622 31288 20628 31303
rect 20680 31288 20686 31340
rect 21818 31288 21824 31340
rect 21876 31288 21882 31340
rect 21928 31328 21956 31368
rect 22005 31365 22017 31399
rect 22051 31396 22063 31399
rect 22281 31399 22339 31405
rect 22051 31368 22085 31396
rect 22051 31365 22063 31368
rect 22005 31359 22063 31365
rect 22281 31365 22293 31399
rect 22327 31396 22339 31399
rect 22327 31368 22867 31396
rect 22327 31365 22339 31368
rect 22281 31359 22339 31365
rect 22186 31328 22192 31340
rect 21928 31300 22192 31328
rect 22186 31288 22192 31300
rect 22244 31328 22250 31340
rect 22511 31331 22569 31337
rect 22511 31328 22523 31331
rect 22244 31300 22523 31328
rect 22244 31288 22250 31300
rect 22511 31297 22523 31300
rect 22557 31297 22569 31331
rect 22511 31291 22569 31297
rect 22630 31331 22688 31337
rect 22630 31297 22642 31331
rect 22676 31328 22688 31331
rect 22676 31297 22692 31328
rect 22630 31291 22692 31297
rect 20438 31260 20444 31272
rect 20364 31232 20444 31260
rect 19168 31204 19196 31232
rect 20438 31220 20444 31232
rect 20496 31260 20502 31272
rect 20496 31232 20944 31260
rect 20496 31220 20502 31232
rect 8720 31164 8892 31192
rect 15948 31164 17356 31192
rect 17497 31195 17555 31201
rect 8720 31152 8726 31164
rect 1857 31127 1915 31133
rect 1857 31093 1869 31127
rect 1903 31124 1915 31127
rect 3329 31127 3387 31133
rect 3329 31124 3341 31127
rect 1903 31096 3341 31124
rect 1903 31093 1915 31096
rect 1857 31087 1915 31093
rect 3329 31093 3341 31096
rect 3375 31124 3387 31127
rect 3694 31124 3700 31136
rect 3375 31096 3700 31124
rect 3375 31093 3387 31096
rect 3329 31087 3387 31093
rect 3694 31084 3700 31096
rect 3752 31084 3758 31136
rect 4614 31084 4620 31136
rect 4672 31084 4678 31136
rect 7650 31084 7656 31136
rect 7708 31124 7714 31136
rect 8573 31127 8631 31133
rect 8573 31124 8585 31127
rect 7708 31096 8585 31124
rect 7708 31084 7714 31096
rect 8573 31093 8585 31096
rect 8619 31093 8631 31127
rect 8573 31087 8631 31093
rect 9217 31127 9275 31133
rect 9217 31093 9229 31127
rect 9263 31124 9275 31127
rect 10778 31124 10784 31136
rect 9263 31096 10784 31124
rect 9263 31093 9275 31096
rect 9217 31087 9275 31093
rect 10778 31084 10784 31096
rect 10836 31084 10842 31136
rect 10962 31084 10968 31136
rect 11020 31084 11026 31136
rect 11698 31084 11704 31136
rect 11756 31124 11762 31136
rect 12434 31124 12440 31136
rect 11756 31096 12440 31124
rect 11756 31084 11762 31096
rect 12434 31084 12440 31096
rect 12492 31124 12498 31136
rect 12897 31127 12955 31133
rect 12897 31124 12909 31127
rect 12492 31096 12909 31124
rect 12492 31084 12498 31096
rect 12897 31093 12909 31096
rect 12943 31093 12955 31127
rect 12897 31087 12955 31093
rect 14550 31084 14556 31136
rect 14608 31084 14614 31136
rect 14826 31084 14832 31136
rect 14884 31124 14890 31136
rect 15948 31124 15976 31164
rect 17497 31161 17509 31195
rect 17543 31192 17555 31195
rect 17543 31164 18644 31192
rect 17543 31161 17555 31164
rect 17497 31155 17555 31161
rect 14884 31096 15976 31124
rect 14884 31084 14890 31096
rect 16390 31084 16396 31136
rect 16448 31084 16454 31136
rect 17126 31084 17132 31136
rect 17184 31124 17190 31136
rect 17221 31127 17279 31133
rect 17221 31124 17233 31127
rect 17184 31096 17233 31124
rect 17184 31084 17190 31096
rect 17221 31093 17233 31096
rect 17267 31093 17279 31127
rect 17221 31087 17279 31093
rect 17862 31084 17868 31136
rect 17920 31124 17926 31136
rect 18325 31127 18383 31133
rect 18325 31124 18337 31127
rect 17920 31096 18337 31124
rect 17920 31084 17926 31096
rect 18325 31093 18337 31096
rect 18371 31124 18383 31127
rect 18414 31124 18420 31136
rect 18371 31096 18420 31124
rect 18371 31093 18383 31096
rect 18325 31087 18383 31093
rect 18414 31084 18420 31096
rect 18472 31084 18478 31136
rect 18616 31124 18644 31164
rect 19150 31152 19156 31204
rect 19208 31152 19214 31204
rect 19242 31152 19248 31204
rect 19300 31192 19306 31204
rect 19429 31195 19487 31201
rect 19429 31192 19441 31195
rect 19300 31164 19441 31192
rect 19300 31152 19306 31164
rect 19429 31161 19441 31164
rect 19475 31192 19487 31195
rect 20806 31192 20812 31204
rect 19475 31164 20812 31192
rect 19475 31161 19487 31164
rect 19429 31155 19487 31161
rect 20806 31152 20812 31164
rect 20864 31152 20870 31204
rect 20916 31192 20944 31232
rect 20990 31220 20996 31272
rect 21048 31220 21054 31272
rect 21836 31192 21864 31288
rect 20916 31164 21864 31192
rect 22189 31195 22247 31201
rect 21376 31136 21404 31164
rect 22189 31161 22201 31195
rect 22235 31192 22247 31195
rect 22554 31192 22560 31204
rect 22235 31164 22560 31192
rect 22235 31161 22247 31164
rect 22189 31155 22247 31161
rect 22554 31152 22560 31164
rect 22612 31152 22618 31204
rect 22664 31192 22692 31291
rect 22738 31288 22744 31340
rect 22796 31288 22802 31340
rect 22839 31260 22867 31368
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 23842 31328 23848 31340
rect 22980 31300 23848 31328
rect 22980 31288 22986 31300
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24596 31328 24624 31424
rect 24762 31356 24768 31408
rect 24820 31356 24826 31408
rect 24854 31356 24860 31408
rect 24912 31356 24918 31408
rect 25314 31396 25320 31408
rect 25240 31368 25320 31396
rect 24673 31331 24731 31337
rect 24673 31328 24685 31331
rect 24596 31300 24685 31328
rect 24673 31297 24685 31300
rect 24719 31297 24731 31331
rect 24673 31291 24731 31297
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 25240 31337 25268 31368
rect 25314 31356 25320 31368
rect 25372 31356 25378 31408
rect 25424 31405 25452 31436
rect 25866 31424 25872 31436
rect 25924 31424 25930 31476
rect 25958 31424 25964 31476
rect 26016 31464 26022 31476
rect 26697 31467 26755 31473
rect 26697 31464 26709 31467
rect 26016 31436 26709 31464
rect 26016 31424 26022 31436
rect 26697 31433 26709 31436
rect 26743 31433 26755 31467
rect 26697 31427 26755 31433
rect 27617 31467 27675 31473
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 28350 31464 28356 31476
rect 27663 31436 28356 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 28350 31424 28356 31436
rect 28408 31424 28414 31476
rect 29457 31467 29515 31473
rect 29457 31433 29469 31467
rect 29503 31464 29515 31467
rect 29503 31436 29776 31464
rect 29503 31433 29515 31436
rect 29457 31427 29515 31433
rect 25409 31399 25467 31405
rect 25409 31365 25421 31399
rect 25455 31365 25467 31399
rect 25409 31359 25467 31365
rect 25608 31368 25820 31396
rect 25608 31340 25636 31368
rect 25041 31331 25099 31337
rect 25041 31328 25053 31331
rect 25004 31300 25053 31328
rect 25004 31288 25010 31300
rect 25041 31297 25053 31300
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31297 25283 31331
rect 25225 31291 25283 31297
rect 23017 31263 23075 31269
rect 23017 31260 23029 31263
rect 22839 31232 23029 31260
rect 23017 31229 23029 31232
rect 23063 31229 23075 31263
rect 23017 31223 23075 31229
rect 24394 31220 24400 31272
rect 24452 31260 24458 31272
rect 25148 31260 25176 31291
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31297 25743 31331
rect 25792 31328 25820 31368
rect 26234 31356 26240 31408
rect 26292 31356 26298 31408
rect 27724 31368 28672 31396
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 25792 31300 25881 31328
rect 25685 31291 25743 31297
rect 25869 31297 25881 31300
rect 25915 31297 25927 31331
rect 26252 31328 26280 31356
rect 27724 31340 27752 31368
rect 25869 31291 25927 31297
rect 25976 31300 26280 31328
rect 24452 31232 25176 31260
rect 25700 31260 25728 31291
rect 25976 31260 26004 31300
rect 26326 31288 26332 31340
rect 26384 31288 26390 31340
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31328 26479 31331
rect 26510 31328 26516 31340
rect 26467 31300 26516 31328
rect 26467 31297 26479 31300
rect 26421 31291 26479 31297
rect 26510 31288 26516 31300
rect 26568 31288 26574 31340
rect 26605 31331 26663 31337
rect 26605 31297 26617 31331
rect 26651 31328 26663 31331
rect 26694 31328 26700 31340
rect 26651 31300 26700 31328
rect 26651 31297 26663 31300
rect 26605 31291 26663 31297
rect 26694 31288 26700 31300
rect 26752 31288 26758 31340
rect 26789 31331 26847 31337
rect 26789 31297 26801 31331
rect 26835 31328 26847 31331
rect 27338 31328 27344 31340
rect 26835 31300 27344 31328
rect 26835 31297 26847 31300
rect 26789 31291 26847 31297
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27614 31328 27620 31340
rect 27586 31288 27620 31328
rect 27672 31288 27678 31340
rect 27706 31288 27712 31340
rect 27764 31288 27770 31340
rect 27798 31288 27804 31340
rect 27856 31328 27862 31340
rect 27985 31331 28043 31337
rect 27985 31328 27997 31331
rect 27856 31300 27997 31328
rect 27856 31288 27862 31300
rect 27985 31297 27997 31300
rect 28031 31297 28043 31331
rect 27985 31291 28043 31297
rect 28074 31288 28080 31340
rect 28132 31328 28138 31340
rect 28350 31328 28356 31340
rect 28132 31300 28356 31328
rect 28132 31288 28138 31300
rect 28350 31288 28356 31300
rect 28408 31328 28414 31340
rect 28644 31337 28672 31368
rect 28445 31331 28503 31337
rect 28445 31328 28457 31331
rect 28408 31300 28457 31328
rect 28408 31288 28414 31300
rect 28445 31297 28457 31300
rect 28491 31297 28503 31331
rect 28445 31291 28503 31297
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31328 28687 31331
rect 29089 31331 29147 31337
rect 29089 31328 29101 31331
rect 28675 31300 29101 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 29089 31297 29101 31300
rect 29135 31297 29147 31331
rect 29089 31291 29147 31297
rect 29365 31331 29423 31337
rect 29365 31297 29377 31331
rect 29411 31297 29423 31331
rect 29365 31291 29423 31297
rect 25700 31232 26004 31260
rect 24452 31220 24458 31232
rect 26142 31220 26148 31272
rect 26200 31220 26206 31272
rect 26237 31263 26295 31269
rect 26237 31229 26249 31263
rect 26283 31260 26295 31263
rect 27586 31260 27614 31288
rect 28169 31263 28227 31269
rect 28169 31260 28181 31263
rect 26283 31232 27614 31260
rect 27693 31232 28181 31260
rect 26283 31229 26295 31232
rect 26237 31223 26295 31229
rect 25685 31195 25743 31201
rect 25685 31192 25697 31195
rect 22664 31164 25697 31192
rect 25332 31136 25360 31164
rect 25685 31161 25697 31164
rect 25731 31161 25743 31195
rect 25685 31155 25743 31161
rect 25958 31152 25964 31204
rect 26016 31152 26022 31204
rect 27693 31192 27721 31232
rect 28169 31229 28181 31232
rect 28215 31260 28227 31263
rect 28902 31260 28908 31272
rect 28215 31232 28908 31260
rect 28215 31229 28227 31232
rect 28169 31223 28227 31229
rect 28902 31220 28908 31232
rect 28960 31220 28966 31272
rect 29380 31260 29408 31291
rect 29546 31288 29552 31340
rect 29604 31288 29610 31340
rect 29748 31328 29776 31436
rect 29897 31331 29955 31337
rect 29897 31328 29909 31331
rect 29748 31300 29909 31328
rect 29897 31297 29909 31300
rect 29943 31297 29955 31331
rect 29897 31291 29955 31297
rect 31573 31331 31631 31337
rect 31573 31297 31585 31331
rect 31619 31328 31631 31331
rect 32122 31328 32128 31340
rect 31619 31300 32128 31328
rect 31619 31297 31631 31300
rect 31573 31291 31631 31297
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 29641 31263 29699 31269
rect 29380 31232 29592 31260
rect 28537 31195 28595 31201
rect 28537 31192 28549 31195
rect 27264 31164 27721 31192
rect 27816 31164 28549 31192
rect 27264 31136 27292 31164
rect 20530 31124 20536 31136
rect 18616 31096 20536 31124
rect 20530 31084 20536 31096
rect 20588 31084 20594 31136
rect 20717 31127 20775 31133
rect 20717 31093 20729 31127
rect 20763 31124 20775 31127
rect 21174 31124 21180 31136
rect 20763 31096 21180 31124
rect 20763 31093 20775 31096
rect 20717 31087 20775 31093
rect 21174 31084 21180 31096
rect 21232 31084 21238 31136
rect 21358 31084 21364 31136
rect 21416 31084 21422 31136
rect 21634 31084 21640 31136
rect 21692 31084 21698 31136
rect 22278 31084 22284 31136
rect 22336 31124 22342 31136
rect 23750 31124 23756 31136
rect 22336 31096 23756 31124
rect 22336 31084 22342 31096
rect 23750 31084 23756 31096
rect 23808 31084 23814 31136
rect 25314 31084 25320 31136
rect 25372 31084 25378 31136
rect 25501 31127 25559 31133
rect 25501 31093 25513 31127
rect 25547 31124 25559 31127
rect 25866 31124 25872 31136
rect 25547 31096 25872 31124
rect 25547 31093 25559 31096
rect 25501 31087 25559 31093
rect 25866 31084 25872 31096
rect 25924 31084 25930 31136
rect 26050 31084 26056 31136
rect 26108 31124 26114 31136
rect 26418 31124 26424 31136
rect 26108 31096 26424 31124
rect 26108 31084 26114 31096
rect 26418 31084 26424 31096
rect 26476 31084 26482 31136
rect 27246 31084 27252 31136
rect 27304 31084 27310 31136
rect 27614 31084 27620 31136
rect 27672 31124 27678 31136
rect 27816 31124 27844 31164
rect 28537 31161 28549 31164
rect 28583 31161 28595 31195
rect 28537 31155 28595 31161
rect 29564 31136 29592 31232
rect 29641 31229 29653 31263
rect 29687 31229 29699 31263
rect 29641 31223 29699 31229
rect 27672 31096 27844 31124
rect 27672 31084 27678 31096
rect 27890 31084 27896 31136
rect 27948 31124 27954 31136
rect 28902 31124 28908 31136
rect 27948 31096 28908 31124
rect 27948 31084 27954 31096
rect 28902 31084 28908 31096
rect 28960 31084 28966 31136
rect 29546 31084 29552 31136
rect 29604 31084 29610 31136
rect 29656 31124 29684 31223
rect 30926 31192 30932 31204
rect 30668 31164 30932 31192
rect 30282 31124 30288 31136
rect 29656 31096 30288 31124
rect 30282 31084 30288 31096
rect 30340 31124 30346 31136
rect 30668 31124 30696 31164
rect 30926 31152 30932 31164
rect 30984 31152 30990 31204
rect 30340 31096 30696 31124
rect 30340 31084 30346 31096
rect 30742 31084 30748 31136
rect 30800 31124 30806 31136
rect 31018 31124 31024 31136
rect 30800 31096 31024 31124
rect 30800 31084 30806 31096
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 31389 31127 31447 31133
rect 31389 31093 31401 31127
rect 31435 31124 31447 31127
rect 31662 31124 31668 31136
rect 31435 31096 31668 31124
rect 31435 31093 31447 31096
rect 31389 31087 31447 31093
rect 31662 31084 31668 31096
rect 31720 31084 31726 31136
rect 31754 31084 31760 31136
rect 31812 31084 31818 31136
rect 1104 31034 43884 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 43884 31034
rect 1104 30960 43884 30982
rect 2498 30880 2504 30932
rect 2556 30920 2562 30932
rect 2869 30923 2927 30929
rect 2869 30920 2881 30923
rect 2556 30892 2881 30920
rect 2556 30880 2562 30892
rect 2869 30889 2881 30892
rect 2915 30889 2927 30923
rect 2869 30883 2927 30889
rect 3970 30880 3976 30932
rect 4028 30880 4034 30932
rect 4062 30880 4068 30932
rect 4120 30920 4126 30932
rect 4525 30923 4583 30929
rect 4525 30920 4537 30923
rect 4120 30892 4537 30920
rect 4120 30880 4126 30892
rect 4525 30889 4537 30892
rect 4571 30889 4583 30923
rect 4525 30883 4583 30889
rect 4798 30880 4804 30932
rect 4856 30880 4862 30932
rect 4982 30880 4988 30932
rect 5040 30920 5046 30932
rect 5721 30923 5779 30929
rect 5721 30920 5733 30923
rect 5040 30892 5733 30920
rect 5040 30880 5046 30892
rect 5721 30889 5733 30892
rect 5767 30889 5779 30923
rect 5721 30883 5779 30889
rect 6641 30923 6699 30929
rect 6641 30889 6653 30923
rect 6687 30920 6699 30923
rect 6914 30920 6920 30932
rect 6687 30892 6920 30920
rect 6687 30889 6699 30892
rect 6641 30883 6699 30889
rect 6914 30880 6920 30892
rect 6972 30880 6978 30932
rect 7098 30880 7104 30932
rect 7156 30880 7162 30932
rect 8757 30923 8815 30929
rect 8757 30889 8769 30923
rect 8803 30920 8815 30923
rect 8938 30920 8944 30932
rect 8803 30892 8944 30920
rect 8803 30889 8815 30892
rect 8757 30883 8815 30889
rect 8938 30880 8944 30892
rect 8996 30880 9002 30932
rect 9677 30923 9735 30929
rect 9677 30889 9689 30923
rect 9723 30920 9735 30923
rect 9858 30920 9864 30932
rect 9723 30892 9864 30920
rect 9723 30889 9735 30892
rect 9677 30883 9735 30889
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 10594 30880 10600 30932
rect 10652 30920 10658 30932
rect 10965 30923 11023 30929
rect 10965 30920 10977 30923
rect 10652 30892 10977 30920
rect 10652 30880 10658 30892
rect 10965 30889 10977 30892
rect 11011 30889 11023 30923
rect 10965 30883 11023 30889
rect 11149 30923 11207 30929
rect 11149 30889 11161 30923
rect 11195 30920 11207 30923
rect 11606 30920 11612 30932
rect 11195 30892 11612 30920
rect 11195 30889 11207 30892
rect 11149 30883 11207 30889
rect 11606 30880 11612 30892
rect 11664 30880 11670 30932
rect 13722 30880 13728 30932
rect 13780 30920 13786 30932
rect 14093 30923 14151 30929
rect 14093 30920 14105 30923
rect 13780 30892 14105 30920
rect 13780 30880 13786 30892
rect 14093 30889 14105 30892
rect 14139 30889 14151 30923
rect 14093 30883 14151 30889
rect 14550 30880 14556 30932
rect 14608 30920 14614 30932
rect 15010 30920 15016 30932
rect 14608 30892 15016 30920
rect 14608 30880 14614 30892
rect 15010 30880 15016 30892
rect 15068 30880 15074 30932
rect 15197 30923 15255 30929
rect 15197 30889 15209 30923
rect 15243 30920 15255 30923
rect 15470 30920 15476 30932
rect 15243 30892 15476 30920
rect 15243 30889 15255 30892
rect 15197 30883 15255 30889
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 16945 30923 17003 30929
rect 16945 30920 16957 30923
rect 16408 30892 16957 30920
rect 4433 30855 4491 30861
rect 4433 30852 4445 30855
rect 3528 30824 4445 30852
rect 1210 30744 1216 30796
rect 1268 30784 1274 30796
rect 1857 30787 1915 30793
rect 1857 30784 1869 30787
rect 1268 30756 1869 30784
rect 1268 30744 1274 30756
rect 1857 30753 1869 30756
rect 1903 30753 1915 30787
rect 1857 30747 1915 30753
rect 2038 30744 2044 30796
rect 2096 30784 2102 30796
rect 3528 30793 3556 30824
rect 4433 30821 4445 30824
rect 4479 30852 4491 30855
rect 4816 30852 4844 30880
rect 4479 30824 4844 30852
rect 5169 30855 5227 30861
rect 4479 30821 4491 30824
rect 4433 30815 4491 30821
rect 5169 30821 5181 30855
rect 5215 30852 5227 30855
rect 5442 30852 5448 30864
rect 5215 30824 5448 30852
rect 5215 30821 5227 30824
rect 5169 30815 5227 30821
rect 5442 30812 5448 30824
rect 5500 30812 5506 30864
rect 5534 30812 5540 30864
rect 5592 30852 5598 30864
rect 6454 30852 6460 30864
rect 5592 30824 6460 30852
rect 5592 30812 5598 30824
rect 6454 30812 6460 30824
rect 6512 30852 6518 30864
rect 7377 30855 7435 30861
rect 7377 30852 7389 30855
rect 6512 30824 7389 30852
rect 6512 30812 6518 30824
rect 7377 30821 7389 30824
rect 7423 30821 7435 30855
rect 7377 30815 7435 30821
rect 7650 30812 7656 30864
rect 7708 30812 7714 30864
rect 8202 30812 8208 30864
rect 8260 30852 8266 30864
rect 8389 30855 8447 30861
rect 8389 30852 8401 30855
rect 8260 30824 8401 30852
rect 8260 30812 8266 30824
rect 8389 30821 8401 30824
rect 8435 30852 8447 30855
rect 13630 30852 13636 30864
rect 8435 30824 13636 30852
rect 8435 30821 8447 30824
rect 8389 30815 8447 30821
rect 13630 30812 13636 30824
rect 13688 30812 13694 30864
rect 13909 30855 13967 30861
rect 13909 30821 13921 30855
rect 13955 30852 13967 30855
rect 14826 30852 14832 30864
rect 13955 30824 14832 30852
rect 13955 30821 13967 30824
rect 13909 30815 13967 30821
rect 14826 30812 14832 30824
rect 14884 30812 14890 30864
rect 15102 30812 15108 30864
rect 15160 30852 15166 30864
rect 15289 30855 15347 30861
rect 15289 30852 15301 30855
rect 15160 30824 15301 30852
rect 15160 30812 15166 30824
rect 15289 30821 15301 30824
rect 15335 30821 15347 30855
rect 15289 30815 15347 30821
rect 3513 30787 3571 30793
rect 3513 30784 3525 30787
rect 2096 30756 3525 30784
rect 2096 30744 2102 30756
rect 3513 30753 3525 30756
rect 3559 30753 3571 30787
rect 6825 30787 6883 30793
rect 3513 30747 3571 30753
rect 3620 30756 5764 30784
rect 1578 30676 1584 30728
rect 1636 30676 1642 30728
rect 3418 30676 3424 30728
rect 3476 30716 3482 30728
rect 3620 30716 3648 30756
rect 3476 30688 3648 30716
rect 3476 30676 3482 30688
rect 3694 30676 3700 30728
rect 3752 30716 3758 30728
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3752 30688 3801 30716
rect 3752 30676 3758 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 3970 30676 3976 30728
rect 4028 30716 4034 30728
rect 4522 30716 4528 30728
rect 4028 30688 4528 30716
rect 4028 30676 4034 30688
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 4709 30719 4767 30725
rect 4709 30716 4721 30719
rect 4672 30688 4721 30716
rect 4672 30676 4678 30688
rect 4709 30685 4721 30688
rect 4755 30685 4767 30719
rect 4709 30679 4767 30685
rect 4801 30719 4859 30725
rect 4801 30685 4813 30719
rect 4847 30716 4859 30719
rect 4890 30716 4896 30728
rect 4847 30688 4896 30716
rect 4847 30685 4859 30688
rect 4801 30679 4859 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 4982 30676 4988 30728
rect 5040 30676 5046 30728
rect 5077 30719 5135 30725
rect 5077 30685 5089 30719
rect 5123 30685 5135 30719
rect 5077 30679 5135 30685
rect 3326 30608 3332 30660
rect 3384 30608 3390 30660
rect 3988 30648 4016 30676
rect 5092 30648 5120 30679
rect 5350 30676 5356 30728
rect 5408 30676 5414 30728
rect 5626 30676 5632 30728
rect 5684 30676 5690 30728
rect 5736 30725 5764 30756
rect 6825 30753 6837 30787
rect 6871 30784 6883 30787
rect 6871 30756 7880 30784
rect 6871 30753 6883 30756
rect 6825 30747 6883 30753
rect 7300 30725 7328 30756
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30685 5779 30719
rect 5721 30679 5779 30685
rect 5905 30719 5963 30725
rect 5905 30685 5917 30719
rect 5951 30685 5963 30719
rect 5905 30679 5963 30685
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30685 6791 30719
rect 6733 30679 6791 30685
rect 6917 30719 6975 30725
rect 6917 30685 6929 30719
rect 6963 30716 6975 30719
rect 7101 30719 7159 30725
rect 6963 30688 7052 30716
rect 6963 30685 6975 30688
rect 6917 30679 6975 30685
rect 3712 30620 4016 30648
rect 4080 30620 5120 30648
rect 3050 30540 3056 30592
rect 3108 30580 3114 30592
rect 3237 30583 3295 30589
rect 3237 30580 3249 30583
rect 3108 30552 3249 30580
rect 3108 30540 3114 30552
rect 3237 30549 3249 30552
rect 3283 30580 3295 30583
rect 3712 30580 3740 30620
rect 3283 30552 3740 30580
rect 3283 30549 3295 30552
rect 3237 30543 3295 30549
rect 3970 30540 3976 30592
rect 4028 30580 4034 30592
rect 4080 30580 4108 30620
rect 5258 30608 5264 30660
rect 5316 30648 5322 30660
rect 5920 30648 5948 30679
rect 5316 30620 5948 30648
rect 6748 30648 6776 30679
rect 7024 30648 7052 30688
rect 7101 30685 7113 30719
rect 7147 30716 7159 30719
rect 7285 30719 7343 30725
rect 7147 30688 7236 30716
rect 7147 30685 7159 30688
rect 7101 30679 7159 30685
rect 7208 30648 7236 30688
rect 7285 30685 7297 30719
rect 7331 30685 7343 30719
rect 7285 30679 7343 30685
rect 7558 30676 7564 30728
rect 7616 30676 7622 30728
rect 7742 30676 7748 30728
rect 7800 30676 7806 30728
rect 7852 30725 7880 30756
rect 8570 30744 8576 30796
rect 8628 30784 8634 30796
rect 9585 30787 9643 30793
rect 9585 30784 9597 30787
rect 8628 30756 9597 30784
rect 8628 30744 8634 30756
rect 9585 30753 9597 30756
rect 9631 30753 9643 30787
rect 9585 30747 9643 30753
rect 10321 30787 10379 30793
rect 10321 30753 10333 30787
rect 10367 30784 10379 30787
rect 10594 30784 10600 30796
rect 10367 30756 10600 30784
rect 10367 30753 10379 30756
rect 10321 30747 10379 30753
rect 10594 30744 10600 30756
rect 10652 30744 10658 30796
rect 10778 30744 10784 30796
rect 10836 30784 10842 30796
rect 11609 30787 11667 30793
rect 11609 30784 11621 30787
rect 10836 30756 11621 30784
rect 10836 30744 10842 30756
rect 11609 30753 11621 30756
rect 11655 30753 11667 30787
rect 11609 30747 11667 30753
rect 11793 30787 11851 30793
rect 11793 30753 11805 30787
rect 11839 30784 11851 30787
rect 11882 30784 11888 30796
rect 11839 30756 11888 30784
rect 11839 30753 11851 30756
rect 11793 30747 11851 30753
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 12805 30787 12863 30793
rect 12805 30753 12817 30787
rect 12851 30784 12863 30787
rect 12986 30784 12992 30796
rect 12851 30756 12992 30784
rect 12851 30753 12863 30756
rect 12805 30747 12863 30753
rect 12986 30744 12992 30756
rect 13044 30744 13050 30796
rect 14737 30787 14795 30793
rect 14737 30753 14749 30787
rect 14783 30784 14795 30787
rect 14918 30784 14924 30796
rect 14783 30756 14924 30784
rect 14783 30753 14795 30756
rect 14737 30747 14795 30753
rect 14918 30744 14924 30756
rect 14976 30744 14982 30796
rect 15746 30744 15752 30796
rect 15804 30744 15810 30796
rect 15933 30787 15991 30793
rect 15933 30753 15945 30787
rect 15979 30784 15991 30787
rect 16408 30784 16436 30892
rect 16945 30889 16957 30892
rect 16991 30889 17003 30923
rect 16945 30883 17003 30889
rect 17310 30880 17316 30932
rect 17368 30920 17374 30932
rect 17497 30923 17555 30929
rect 17497 30920 17509 30923
rect 17368 30892 17509 30920
rect 17368 30880 17374 30892
rect 17497 30889 17509 30892
rect 17543 30889 17555 30923
rect 17497 30883 17555 30889
rect 17586 30880 17592 30932
rect 17644 30880 17650 30932
rect 18138 30880 18144 30932
rect 18196 30920 18202 30932
rect 18598 30920 18604 30932
rect 18196 30892 18604 30920
rect 18196 30880 18202 30892
rect 18598 30880 18604 30892
rect 18656 30880 18662 30932
rect 18690 30880 18696 30932
rect 18748 30880 18754 30932
rect 19812 30892 22094 30920
rect 17037 30855 17095 30861
rect 17037 30821 17049 30855
rect 17083 30852 17095 30855
rect 17604 30852 17632 30880
rect 17083 30824 17632 30852
rect 17865 30855 17923 30861
rect 17083 30821 17095 30824
rect 17037 30815 17095 30821
rect 17865 30821 17877 30855
rect 17911 30852 17923 30855
rect 18877 30855 18935 30861
rect 18877 30852 18889 30855
rect 17911 30824 18889 30852
rect 17911 30821 17923 30824
rect 17865 30815 17923 30821
rect 18877 30821 18889 30824
rect 18923 30821 18935 30855
rect 18877 30815 18935 30821
rect 17052 30784 17080 30815
rect 15979 30756 16436 30784
rect 16776 30756 17080 30784
rect 18049 30787 18107 30793
rect 15979 30753 15991 30756
rect 15933 30747 15991 30753
rect 7837 30719 7895 30725
rect 7837 30685 7849 30719
rect 7883 30685 7895 30719
rect 7837 30679 7895 30685
rect 9214 30676 9220 30728
rect 9272 30676 9278 30728
rect 9401 30719 9459 30725
rect 9401 30685 9413 30719
rect 9447 30716 9459 30719
rect 9490 30716 9496 30728
rect 9447 30688 9496 30716
rect 9447 30685 9459 30688
rect 9401 30679 9459 30685
rect 9490 30676 9496 30688
rect 9548 30676 9554 30728
rect 10042 30676 10048 30728
rect 10100 30676 10106 30728
rect 11517 30719 11575 30725
rect 11517 30685 11529 30719
rect 11563 30716 11575 30719
rect 11563 30688 12112 30716
rect 11563 30685 11575 30688
rect 11517 30679 11575 30685
rect 12084 30660 12112 30688
rect 12158 30676 12164 30728
rect 12216 30676 12222 30728
rect 12437 30719 12495 30725
rect 12437 30716 12449 30719
rect 12268 30688 12449 30716
rect 12268 30660 12296 30688
rect 12437 30685 12449 30688
rect 12483 30685 12495 30719
rect 12437 30679 12495 30685
rect 12710 30676 12716 30728
rect 12768 30676 12774 30728
rect 13449 30719 13507 30725
rect 13449 30716 13461 30719
rect 13004 30688 13461 30716
rect 6748 30620 6960 30648
rect 7024 30620 7144 30648
rect 7208 30620 7880 30648
rect 5316 30608 5322 30620
rect 6932 30592 6960 30620
rect 7116 30592 7144 30620
rect 7852 30592 7880 30620
rect 9306 30608 9312 30660
rect 9364 30648 9370 30660
rect 10137 30651 10195 30657
rect 10137 30648 10149 30651
rect 9364 30620 10149 30648
rect 9364 30608 9370 30620
rect 10137 30617 10149 30620
rect 10183 30617 10195 30651
rect 10137 30611 10195 30617
rect 10870 30608 10876 30660
rect 10928 30648 10934 30660
rect 11977 30651 12035 30657
rect 11977 30648 11989 30651
rect 10928 30620 11989 30648
rect 10928 30608 10934 30620
rect 11977 30617 11989 30620
rect 12023 30617 12035 30651
rect 11977 30611 12035 30617
rect 12066 30608 12072 30660
rect 12124 30608 12130 30660
rect 12250 30608 12256 30660
rect 12308 30608 12314 30660
rect 12345 30651 12403 30657
rect 12345 30617 12357 30651
rect 12391 30648 12403 30651
rect 12728 30648 12756 30676
rect 12391 30620 12756 30648
rect 12391 30617 12403 30620
rect 12345 30611 12403 30617
rect 4028 30552 4108 30580
rect 4028 30540 4034 30552
rect 4522 30540 4528 30592
rect 4580 30580 4586 30592
rect 6273 30583 6331 30589
rect 6273 30580 6285 30583
rect 4580 30552 6285 30580
rect 4580 30540 4586 30552
rect 6273 30549 6285 30552
rect 6319 30580 6331 30583
rect 6454 30580 6460 30592
rect 6319 30552 6460 30580
rect 6319 30549 6331 30552
rect 6273 30543 6331 30549
rect 6454 30540 6460 30552
rect 6512 30540 6518 30592
rect 6914 30540 6920 30592
rect 6972 30540 6978 30592
rect 7098 30540 7104 30592
rect 7156 30540 7162 30592
rect 7834 30540 7840 30592
rect 7892 30540 7898 30592
rect 8938 30540 8944 30592
rect 8996 30580 9002 30592
rect 13004 30580 13032 30688
rect 13449 30685 13461 30688
rect 13495 30716 13507 30719
rect 13495 30688 16620 30716
rect 13495 30685 13507 30688
rect 13449 30679 13507 30685
rect 14553 30651 14611 30657
rect 14553 30648 14565 30651
rect 13096 30620 14565 30648
rect 13096 30589 13124 30620
rect 14553 30617 14565 30620
rect 14599 30617 14611 30651
rect 14553 30611 14611 30617
rect 16301 30651 16359 30657
rect 16301 30617 16313 30651
rect 16347 30617 16359 30651
rect 16592 30648 16620 30688
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 16776 30725 16804 30756
rect 18049 30753 18061 30787
rect 18095 30784 18107 30787
rect 18690 30784 18696 30796
rect 18095 30756 18696 30784
rect 18095 30753 18107 30756
rect 18049 30747 18107 30753
rect 18690 30744 18696 30756
rect 18748 30744 18754 30796
rect 19334 30784 19340 30796
rect 18800 30756 19340 30784
rect 16761 30719 16819 30725
rect 16761 30685 16773 30719
rect 16807 30685 16819 30719
rect 17310 30716 17316 30728
rect 16761 30679 16819 30685
rect 16868 30688 17316 30716
rect 16868 30648 16896 30688
rect 17310 30676 17316 30688
rect 17368 30676 17374 30728
rect 17770 30676 17776 30728
rect 17828 30676 17834 30728
rect 17954 30676 17960 30728
rect 18012 30676 18018 30728
rect 18233 30719 18291 30725
rect 18233 30685 18245 30719
rect 18279 30685 18291 30719
rect 18233 30679 18291 30685
rect 16592 30620 16896 30648
rect 17037 30651 17095 30657
rect 16301 30611 16359 30617
rect 17037 30617 17049 30651
rect 17083 30648 17095 30651
rect 17678 30648 17684 30660
rect 17083 30620 17684 30648
rect 17083 30617 17095 30620
rect 17037 30611 17095 30617
rect 8996 30552 13032 30580
rect 13081 30583 13139 30589
rect 8996 30540 9002 30552
rect 13081 30549 13093 30583
rect 13127 30549 13139 30583
rect 13081 30543 13139 30549
rect 13722 30540 13728 30592
rect 13780 30580 13786 30592
rect 13906 30580 13912 30592
rect 13780 30552 13912 30580
rect 13780 30540 13786 30552
rect 13906 30540 13912 30552
rect 13964 30540 13970 30592
rect 13998 30540 14004 30592
rect 14056 30580 14062 30592
rect 14366 30580 14372 30592
rect 14056 30552 14372 30580
rect 14056 30540 14062 30552
rect 14366 30540 14372 30552
rect 14424 30540 14430 30592
rect 14458 30540 14464 30592
rect 14516 30540 14522 30592
rect 15654 30540 15660 30592
rect 15712 30540 15718 30592
rect 16316 30580 16344 30611
rect 17678 30608 17684 30620
rect 17736 30608 17742 30660
rect 18248 30648 18276 30679
rect 18322 30676 18328 30728
rect 18380 30676 18386 30728
rect 18414 30676 18420 30728
rect 18472 30716 18478 30728
rect 18800 30716 18828 30756
rect 19334 30744 19340 30756
rect 19392 30744 19398 30796
rect 18472 30688 18828 30716
rect 18472 30676 18478 30688
rect 19242 30676 19248 30728
rect 19300 30676 19306 30728
rect 19812 30725 19840 30892
rect 20438 30852 20444 30864
rect 19996 30824 20444 30852
rect 19996 30725 20024 30824
rect 20438 30812 20444 30824
rect 20496 30812 20502 30864
rect 22066 30852 22094 30892
rect 22462 30880 22468 30932
rect 22520 30920 22526 30932
rect 22922 30920 22928 30932
rect 22520 30892 22928 30920
rect 22520 30880 22526 30892
rect 22922 30880 22928 30892
rect 22980 30880 22986 30932
rect 23293 30923 23351 30929
rect 23293 30889 23305 30923
rect 23339 30920 23351 30923
rect 24302 30920 24308 30932
rect 23339 30892 24308 30920
rect 23339 30889 23351 30892
rect 23293 30883 23351 30889
rect 24302 30880 24308 30892
rect 24360 30880 24366 30932
rect 24394 30880 24400 30932
rect 24452 30880 24458 30932
rect 24486 30880 24492 30932
rect 24544 30880 24550 30932
rect 24578 30880 24584 30932
rect 24636 30920 24642 30932
rect 24636 30892 26096 30920
rect 24636 30880 24642 30892
rect 23934 30852 23940 30864
rect 22066 30824 23940 30852
rect 23934 30812 23940 30824
rect 23992 30812 23998 30864
rect 24118 30812 24124 30864
rect 24176 30812 24182 30864
rect 20346 30744 20352 30796
rect 20404 30784 20410 30796
rect 20404 30756 20484 30784
rect 20404 30744 20410 30756
rect 20456 30725 20484 30756
rect 20714 30744 20720 30796
rect 20772 30744 20778 30796
rect 20898 30744 20904 30796
rect 20956 30744 20962 30796
rect 23201 30787 23259 30793
rect 21928 30756 23152 30784
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30685 19855 30719
rect 19797 30679 19855 30685
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20165 30719 20223 30725
rect 20165 30685 20177 30719
rect 20211 30716 20223 30719
rect 20441 30719 20499 30725
rect 20211 30692 20224 30716
rect 20211 30685 20392 30692
rect 20165 30679 20392 30685
rect 20441 30685 20453 30719
rect 20487 30685 20499 30719
rect 20732 30716 20760 30744
rect 21928 30716 21956 30756
rect 20732 30688 21956 30716
rect 20441 30679 20499 30685
rect 18506 30648 18512 30660
rect 18248 30620 18512 30648
rect 18506 30608 18512 30620
rect 18564 30608 18570 30660
rect 18598 30608 18604 30660
rect 18656 30648 18662 30660
rect 18693 30651 18751 30657
rect 18693 30648 18705 30651
rect 18656 30620 18705 30648
rect 18656 30608 18662 30620
rect 18693 30617 18705 30620
rect 18739 30617 18751 30651
rect 18693 30611 18751 30617
rect 18782 30608 18788 30660
rect 18840 30648 18846 30660
rect 19334 30648 19340 30660
rect 18840 30620 19340 30648
rect 18840 30608 18846 30620
rect 19334 30608 19340 30620
rect 19392 30608 19398 30660
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30648 19579 30651
rect 19996 30648 20024 30679
rect 20196 30664 20392 30679
rect 22002 30676 22008 30728
rect 22060 30716 22066 30728
rect 23124 30725 23152 30756
rect 23201 30753 23213 30787
rect 23247 30784 23259 30787
rect 23474 30784 23480 30796
rect 23247 30756 23480 30784
rect 23247 30753 23259 30756
rect 23201 30747 23259 30753
rect 23474 30744 23480 30756
rect 23532 30744 23538 30796
rect 23566 30744 23572 30796
rect 23624 30784 23630 30796
rect 24136 30784 24164 30812
rect 23624 30756 24164 30784
rect 24412 30784 24440 30880
rect 24504 30852 24532 30880
rect 24504 30824 25176 30852
rect 24489 30787 24547 30793
rect 24489 30784 24501 30787
rect 24412 30756 24501 30784
rect 23624 30744 23630 30756
rect 24489 30753 24501 30756
rect 24535 30753 24547 30787
rect 24489 30747 24547 30753
rect 24578 30744 24584 30796
rect 24636 30744 24642 30796
rect 24670 30744 24676 30796
rect 24728 30744 24734 30796
rect 24762 30744 24768 30796
rect 24820 30744 24826 30796
rect 24946 30744 24952 30796
rect 25004 30744 25010 30796
rect 22373 30719 22431 30725
rect 22373 30716 22385 30719
rect 22060 30688 22385 30716
rect 22060 30676 22066 30688
rect 22373 30685 22385 30688
rect 22419 30685 22431 30719
rect 22373 30679 22431 30685
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 23842 30676 23848 30728
rect 23900 30676 23906 30728
rect 24596 30716 24624 30744
rect 25148 30725 25176 30824
rect 25774 30812 25780 30864
rect 25832 30812 25838 30864
rect 24857 30719 24915 30725
rect 24857 30716 24869 30719
rect 24596 30688 24869 30716
rect 24857 30685 24869 30688
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30685 25191 30719
rect 25133 30679 25191 30685
rect 25314 30676 25320 30728
rect 25372 30676 25378 30728
rect 25406 30676 25412 30728
rect 25464 30676 25470 30728
rect 25593 30719 25651 30725
rect 25593 30685 25605 30719
rect 25639 30716 25651 30719
rect 25792 30716 25820 30812
rect 25639 30688 25820 30716
rect 26068 30716 26096 30892
rect 26142 30880 26148 30932
rect 26200 30920 26206 30932
rect 27341 30923 27399 30929
rect 27341 30920 27353 30923
rect 26200 30892 27353 30920
rect 26200 30880 26206 30892
rect 27341 30889 27353 30892
rect 27387 30889 27399 30923
rect 27341 30883 27399 30889
rect 28166 30880 28172 30932
rect 28224 30880 28230 30932
rect 28442 30880 28448 30932
rect 28500 30880 28506 30932
rect 29546 30880 29552 30932
rect 29604 30880 29610 30932
rect 30653 30923 30711 30929
rect 30653 30889 30665 30923
rect 30699 30920 30711 30923
rect 32398 30920 32404 30932
rect 30699 30892 32404 30920
rect 30699 30889 30711 30892
rect 30653 30883 30711 30889
rect 32398 30880 32404 30892
rect 32456 30880 32462 30932
rect 26326 30812 26332 30864
rect 26384 30812 26390 30864
rect 26510 30812 26516 30864
rect 26568 30852 26574 30864
rect 26970 30852 26976 30864
rect 26568 30824 26976 30852
rect 26568 30812 26574 30824
rect 26970 30812 26976 30824
rect 27028 30852 27034 30864
rect 27614 30852 27620 30864
rect 27028 30824 27620 30852
rect 27028 30812 27034 30824
rect 27356 30784 27384 30824
rect 27614 30812 27620 30824
rect 27672 30812 27678 30864
rect 28718 30812 28724 30864
rect 28776 30852 28782 30864
rect 28776 30824 30788 30852
rect 28776 30812 28782 30824
rect 27356 30756 27476 30784
rect 26068 30688 26832 30716
rect 25639 30685 25651 30688
rect 25593 30679 25651 30685
rect 19567 30620 20024 30648
rect 20364 30648 20392 30664
rect 20714 30648 20720 30660
rect 20364 30620 20720 30648
rect 19567 30617 19579 30620
rect 19521 30611 19579 30617
rect 20714 30608 20720 30620
rect 20772 30608 20778 30660
rect 21168 30651 21226 30657
rect 21168 30617 21180 30651
rect 21214 30648 21226 30651
rect 23017 30651 23075 30657
rect 23017 30648 23029 30651
rect 21214 30620 23029 30648
rect 21214 30617 21226 30620
rect 21168 30611 21226 30617
rect 23017 30617 23029 30620
rect 23063 30617 23075 30651
rect 24486 30648 24492 30660
rect 23017 30611 23075 30617
rect 23492 30620 24492 30648
rect 17126 30580 17132 30592
rect 16316 30552 17132 30580
rect 17126 30540 17132 30552
rect 17184 30540 17190 30592
rect 17221 30583 17279 30589
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 19150 30580 19156 30592
rect 17267 30552 19156 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 19150 30540 19156 30552
rect 19208 30540 19214 30592
rect 19242 30540 19248 30592
rect 19300 30580 19306 30592
rect 19889 30583 19947 30589
rect 19889 30580 19901 30583
rect 19300 30552 19901 30580
rect 19300 30540 19306 30552
rect 19889 30549 19901 30552
rect 19935 30549 19947 30583
rect 19889 30543 19947 30549
rect 20070 30540 20076 30592
rect 20128 30580 20134 30592
rect 20349 30583 20407 30589
rect 20349 30580 20361 30583
rect 20128 30552 20361 30580
rect 20128 30540 20134 30552
rect 20349 30549 20361 30552
rect 20395 30580 20407 30583
rect 20438 30580 20444 30592
rect 20395 30552 20444 30580
rect 20395 30549 20407 30552
rect 20349 30543 20407 30549
rect 20438 30540 20444 30552
rect 20496 30540 20502 30592
rect 20530 30540 20536 30592
rect 20588 30540 20594 30592
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 22281 30583 22339 30589
rect 22281 30580 22293 30583
rect 20956 30552 22293 30580
rect 20956 30540 20962 30552
rect 22281 30549 22293 30552
rect 22327 30549 22339 30583
rect 22281 30543 22339 30549
rect 22738 30540 22744 30592
rect 22796 30580 22802 30592
rect 23106 30580 23112 30592
rect 22796 30552 23112 30580
rect 22796 30540 22802 30552
rect 23106 30540 23112 30552
rect 23164 30540 23170 30592
rect 23492 30589 23520 30620
rect 24486 30608 24492 30620
rect 24544 30608 24550 30660
rect 25038 30608 25044 30660
rect 25096 30648 25102 30660
rect 25096 30620 25453 30648
rect 25096 30608 25102 30620
rect 23477 30583 23535 30589
rect 23477 30549 23489 30583
rect 23523 30549 23535 30583
rect 23477 30543 23535 30549
rect 23658 30540 23664 30592
rect 23716 30580 23722 30592
rect 24394 30580 24400 30592
rect 23716 30552 24400 30580
rect 23716 30540 23722 30552
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 24762 30540 24768 30592
rect 24820 30580 24826 30592
rect 25225 30583 25283 30589
rect 25225 30580 25237 30583
rect 24820 30552 25237 30580
rect 24820 30540 24826 30552
rect 25225 30549 25237 30552
rect 25271 30549 25283 30583
rect 25425 30580 25453 30620
rect 25498 30608 25504 30660
rect 25556 30648 25562 30660
rect 25961 30651 26019 30657
rect 25961 30648 25973 30651
rect 25556 30620 25973 30648
rect 25556 30608 25562 30620
rect 25961 30617 25973 30620
rect 26007 30617 26019 30651
rect 25961 30611 26019 30617
rect 26050 30608 26056 30660
rect 26108 30648 26114 30660
rect 26145 30651 26203 30657
rect 26145 30648 26157 30651
rect 26108 30620 26157 30648
rect 26108 30608 26114 30620
rect 26145 30617 26157 30620
rect 26191 30617 26203 30651
rect 26145 30611 26203 30617
rect 26694 30580 26700 30592
rect 25425 30552 26700 30580
rect 25225 30543 25283 30549
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 26804 30580 26832 30688
rect 27448 30648 27476 30756
rect 27522 30744 27528 30796
rect 27580 30784 27586 30796
rect 28169 30787 28227 30793
rect 28169 30784 28181 30787
rect 27580 30756 28181 30784
rect 27580 30744 27586 30756
rect 28169 30753 28181 30756
rect 28215 30753 28227 30787
rect 28626 30784 28632 30796
rect 28169 30747 28227 30753
rect 28276 30756 28632 30784
rect 27617 30719 27675 30725
rect 27617 30685 27629 30719
rect 27663 30716 27675 30719
rect 28077 30719 28135 30725
rect 28077 30716 28089 30719
rect 27663 30688 28089 30716
rect 27663 30685 27675 30688
rect 27617 30679 27675 30685
rect 28077 30685 28089 30688
rect 28123 30716 28135 30719
rect 28123 30715 28212 30716
rect 28276 30715 28304 30756
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 28810 30744 28816 30796
rect 28868 30744 28874 30796
rect 28123 30688 28304 30715
rect 28123 30685 28135 30688
rect 28184 30687 28304 30688
rect 28077 30679 28135 30685
rect 27893 30651 27951 30657
rect 27893 30648 27905 30651
rect 27448 30620 27905 30648
rect 27893 30617 27905 30620
rect 27939 30617 27951 30651
rect 27893 30611 27951 30617
rect 27985 30651 28043 30657
rect 27985 30617 27997 30651
rect 28031 30648 28043 30651
rect 28442 30648 28448 30660
rect 28031 30620 28448 30648
rect 28031 30617 28043 30620
rect 27985 30611 28043 30617
rect 28000 30580 28028 30611
rect 28442 30608 28448 30620
rect 28500 30648 28506 30660
rect 28629 30651 28687 30657
rect 28629 30648 28641 30651
rect 28500 30620 28641 30648
rect 28500 30608 28506 30620
rect 28629 30617 28641 30620
rect 28675 30648 28687 30651
rect 28828 30648 28856 30744
rect 28902 30676 28908 30728
rect 28960 30676 28966 30728
rect 29012 30716 29040 30824
rect 29270 30744 29276 30796
rect 29328 30784 29334 30796
rect 29328 30756 30512 30784
rect 29328 30744 29334 30756
rect 29840 30725 29868 30756
rect 30484 30728 30512 30756
rect 29733 30719 29791 30725
rect 29733 30716 29745 30719
rect 29012 30688 29745 30716
rect 29733 30685 29745 30688
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 29825 30719 29883 30725
rect 29825 30685 29837 30719
rect 29871 30685 29883 30719
rect 29825 30679 29883 30685
rect 30098 30676 30104 30728
rect 30156 30676 30162 30728
rect 30466 30676 30472 30728
rect 30524 30676 30530 30728
rect 28675 30620 28856 30648
rect 29181 30651 29239 30657
rect 28675 30617 28687 30620
rect 28629 30611 28687 30617
rect 29181 30617 29193 30651
rect 29227 30648 29239 30651
rect 29549 30651 29607 30657
rect 29549 30648 29561 30651
rect 29227 30620 29561 30648
rect 29227 30617 29239 30620
rect 29181 30611 29239 30617
rect 29549 30617 29561 30620
rect 29595 30648 29607 30651
rect 30285 30651 30343 30657
rect 30285 30648 30297 30651
rect 29595 30620 30297 30648
rect 29595 30617 29607 30620
rect 29549 30611 29607 30617
rect 30285 30617 30297 30620
rect 30331 30617 30343 30651
rect 30285 30611 30343 30617
rect 30377 30651 30435 30657
rect 30377 30617 30389 30651
rect 30423 30648 30435 30651
rect 30650 30648 30656 30660
rect 30423 30620 30656 30648
rect 30423 30617 30435 30620
rect 30377 30611 30435 30617
rect 30650 30608 30656 30620
rect 30708 30608 30714 30660
rect 30760 30648 30788 30824
rect 30837 30719 30895 30725
rect 30837 30685 30849 30719
rect 30883 30716 30895 30719
rect 30926 30716 30932 30728
rect 30883 30688 30932 30716
rect 30883 30685 30895 30688
rect 30837 30679 30895 30685
rect 30926 30676 30932 30688
rect 30984 30676 30990 30728
rect 31104 30719 31162 30725
rect 31104 30685 31116 30719
rect 31150 30716 31162 30719
rect 32214 30716 32220 30728
rect 31150 30688 32220 30716
rect 31150 30685 31162 30688
rect 31104 30679 31162 30685
rect 32214 30676 32220 30688
rect 32272 30676 32278 30728
rect 32401 30719 32459 30725
rect 32401 30685 32413 30719
rect 32447 30716 32459 30719
rect 33502 30716 33508 30728
rect 32447 30688 33508 30716
rect 32447 30685 32459 30688
rect 32401 30679 32459 30685
rect 31754 30648 31760 30660
rect 30760 30620 31760 30648
rect 31754 30608 31760 30620
rect 31812 30608 31818 30660
rect 32416 30648 32444 30679
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 31864 30620 32444 30648
rect 26804 30552 28028 30580
rect 28810 30540 28816 30592
rect 28868 30540 28874 30592
rect 28997 30583 29055 30589
rect 28997 30549 29009 30583
rect 29043 30580 29055 30583
rect 30006 30580 30012 30592
rect 29043 30552 30012 30580
rect 29043 30549 29055 30552
rect 28997 30543 29055 30549
rect 30006 30540 30012 30552
rect 30064 30540 30070 30592
rect 31386 30540 31392 30592
rect 31444 30580 31450 30592
rect 31864 30580 31892 30620
rect 31444 30552 31892 30580
rect 31444 30540 31450 30552
rect 31938 30540 31944 30592
rect 31996 30580 32002 30592
rect 32217 30583 32275 30589
rect 32217 30580 32229 30583
rect 31996 30552 32229 30580
rect 31996 30540 32002 30552
rect 32217 30549 32229 30552
rect 32263 30549 32275 30583
rect 32217 30543 32275 30549
rect 32306 30540 32312 30592
rect 32364 30580 32370 30592
rect 32953 30583 33011 30589
rect 32953 30580 32965 30583
rect 32364 30552 32965 30580
rect 32364 30540 32370 30552
rect 32953 30549 32965 30552
rect 32999 30549 33011 30583
rect 32953 30543 33011 30549
rect 1104 30490 43884 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 43884 30490
rect 1104 30416 43884 30438
rect 2038 30336 2044 30388
rect 2096 30336 2102 30388
rect 2777 30379 2835 30385
rect 2777 30345 2789 30379
rect 2823 30376 2835 30379
rect 3326 30376 3332 30388
rect 2823 30348 3332 30376
rect 2823 30345 2835 30348
rect 2777 30339 2835 30345
rect 3326 30336 3332 30348
rect 3384 30336 3390 30388
rect 3804 30348 4292 30376
rect 2225 30311 2283 30317
rect 2225 30277 2237 30311
rect 2271 30308 2283 30311
rect 2271 30280 3096 30308
rect 2271 30277 2283 30280
rect 2225 30271 2283 30277
rect 2130 30200 2136 30252
rect 2188 30200 2194 30252
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30240 2375 30243
rect 2406 30240 2412 30252
rect 2363 30212 2412 30240
rect 2363 30209 2375 30212
rect 2317 30203 2375 30209
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 2498 30200 2504 30252
rect 2556 30200 2562 30252
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30240 2651 30243
rect 2866 30240 2872 30252
rect 2639 30212 2872 30240
rect 2639 30209 2651 30212
rect 2593 30203 2651 30209
rect 2866 30200 2872 30212
rect 2924 30200 2930 30252
rect 3068 30249 3096 30280
rect 3234 30268 3240 30320
rect 3292 30308 3298 30320
rect 3804 30317 3832 30348
rect 3789 30311 3847 30317
rect 3789 30308 3801 30311
rect 3292 30280 3801 30308
rect 3292 30268 3298 30280
rect 3789 30277 3801 30280
rect 3835 30277 3847 30311
rect 3789 30271 3847 30277
rect 3970 30268 3976 30320
rect 4028 30268 4034 30320
rect 4065 30311 4123 30317
rect 4065 30277 4077 30311
rect 4111 30308 4123 30311
rect 4154 30308 4160 30320
rect 4111 30280 4160 30308
rect 4111 30277 4123 30280
rect 4065 30271 4123 30277
rect 4154 30268 4160 30280
rect 4212 30268 4218 30320
rect 4264 30317 4292 30348
rect 4798 30336 4804 30388
rect 4856 30376 4862 30388
rect 4856 30348 5120 30376
rect 4856 30336 4862 30348
rect 4249 30311 4307 30317
rect 4249 30277 4261 30311
rect 4295 30277 4307 30311
rect 4249 30271 4307 30277
rect 4338 30268 4344 30320
rect 4396 30268 4402 30320
rect 4617 30311 4675 30317
rect 4617 30277 4629 30311
rect 4663 30308 4675 30311
rect 4706 30308 4712 30320
rect 4663 30280 4712 30308
rect 4663 30277 4675 30280
rect 4617 30271 4675 30277
rect 4706 30268 4712 30280
rect 4764 30268 4770 30320
rect 5092 30308 5120 30348
rect 5442 30336 5448 30388
rect 5500 30336 5506 30388
rect 5626 30336 5632 30388
rect 5684 30336 5690 30388
rect 6914 30336 6920 30388
rect 6972 30336 6978 30388
rect 7834 30336 7840 30388
rect 7892 30336 7898 30388
rect 8110 30336 8116 30388
rect 8168 30376 8174 30388
rect 8205 30379 8263 30385
rect 8205 30376 8217 30379
rect 8168 30348 8217 30376
rect 8168 30336 8174 30348
rect 8205 30345 8217 30348
rect 8251 30345 8263 30379
rect 8205 30339 8263 30345
rect 9582 30336 9588 30388
rect 9640 30376 9646 30388
rect 9858 30376 9864 30388
rect 9640 30348 9864 30376
rect 9640 30336 9646 30348
rect 9858 30336 9864 30348
rect 9916 30336 9922 30388
rect 10229 30379 10287 30385
rect 10229 30345 10241 30379
rect 10275 30376 10287 30379
rect 10594 30376 10600 30388
rect 10275 30348 10600 30376
rect 10275 30345 10287 30348
rect 10229 30339 10287 30345
rect 10594 30336 10600 30348
rect 10652 30336 10658 30388
rect 10778 30336 10784 30388
rect 10836 30376 10842 30388
rect 10873 30379 10931 30385
rect 10873 30376 10885 30379
rect 10836 30348 10885 30376
rect 10836 30336 10842 30348
rect 10873 30345 10885 30348
rect 10919 30345 10931 30379
rect 11882 30376 11888 30388
rect 10873 30339 10931 30345
rect 10980 30348 11888 30376
rect 5258 30308 5264 30320
rect 5092 30280 5264 30308
rect 3053 30243 3111 30249
rect 3053 30209 3065 30243
rect 3099 30209 3111 30243
rect 3053 30203 3111 30209
rect 2682 30064 2688 30116
rect 2740 30104 2746 30116
rect 3068 30104 3096 30203
rect 3142 30200 3148 30252
rect 3200 30240 3206 30252
rect 3329 30243 3387 30249
rect 3200 30212 3280 30240
rect 3200 30200 3206 30212
rect 3252 30181 3280 30212
rect 3329 30209 3341 30243
rect 3375 30240 3387 30243
rect 3510 30240 3516 30252
rect 3375 30212 3516 30240
rect 3375 30209 3387 30212
rect 3329 30203 3387 30209
rect 3510 30200 3516 30212
rect 3568 30200 3574 30252
rect 3605 30243 3663 30249
rect 3605 30209 3617 30243
rect 3651 30209 3663 30243
rect 3605 30203 3663 30209
rect 3697 30243 3755 30249
rect 3697 30209 3709 30243
rect 3743 30240 3755 30243
rect 4438 30243 4496 30249
rect 4438 30240 4450 30243
rect 3743 30230 3832 30240
rect 3988 30230 4450 30240
rect 3743 30212 4450 30230
rect 3743 30209 3755 30212
rect 3697 30203 3755 30209
rect 3237 30175 3295 30181
rect 3237 30141 3249 30175
rect 3283 30141 3295 30175
rect 3620 30172 3648 30203
rect 3804 30202 4016 30212
rect 4438 30209 4450 30212
rect 4484 30240 4496 30243
rect 4801 30243 4859 30249
rect 4484 30212 4752 30240
rect 4484 30209 4496 30212
rect 4438 30203 4496 30209
rect 4154 30172 4160 30184
rect 3620 30144 4160 30172
rect 3237 30135 3295 30141
rect 4154 30132 4160 30144
rect 4212 30132 4218 30184
rect 4341 30175 4399 30181
rect 4341 30141 4353 30175
rect 4387 30172 4399 30175
rect 4522 30172 4528 30184
rect 4387 30144 4528 30172
rect 4387 30141 4399 30144
rect 4341 30135 4399 30141
rect 4522 30132 4528 30144
rect 4580 30132 4586 30184
rect 3326 30104 3332 30116
rect 2740 30076 2912 30104
rect 3068 30076 3332 30104
rect 2740 30064 2746 30076
rect 2884 30045 2912 30076
rect 3326 30064 3332 30076
rect 3384 30064 3390 30116
rect 3421 30107 3479 30113
rect 3421 30073 3433 30107
rect 3467 30104 3479 30107
rect 4246 30104 4252 30116
rect 3467 30076 4252 30104
rect 3467 30073 3479 30076
rect 3421 30067 3479 30073
rect 4246 30064 4252 30076
rect 4304 30104 4310 30116
rect 4614 30104 4620 30116
rect 4304 30076 4620 30104
rect 4304 30064 4310 30076
rect 4614 30064 4620 30076
rect 4672 30064 4678 30116
rect 4724 30104 4752 30212
rect 4801 30209 4813 30243
rect 4847 30240 4859 30243
rect 4890 30240 4896 30252
rect 4847 30212 4896 30240
rect 4847 30209 4859 30212
rect 4801 30203 4859 30209
rect 4890 30200 4896 30212
rect 4948 30200 4954 30252
rect 5092 30249 5120 30280
rect 5258 30268 5264 30280
rect 5316 30268 5322 30320
rect 5644 30308 5672 30336
rect 5813 30311 5871 30317
rect 5813 30308 5825 30311
rect 5644 30280 5825 30308
rect 5813 30277 5825 30280
rect 5859 30308 5871 30311
rect 7098 30308 7104 30320
rect 5859 30280 7104 30308
rect 5859 30277 5871 30280
rect 5813 30271 5871 30277
rect 7098 30268 7104 30280
rect 7156 30268 7162 30320
rect 10612 30308 10640 30336
rect 10980 30308 11008 30348
rect 11882 30336 11888 30348
rect 11940 30336 11946 30388
rect 12158 30336 12164 30388
rect 12216 30376 12222 30388
rect 12253 30379 12311 30385
rect 12253 30376 12265 30379
rect 12216 30348 12265 30376
rect 12216 30336 12222 30348
rect 12253 30345 12265 30348
rect 12299 30345 12311 30379
rect 12253 30339 12311 30345
rect 8772 30280 9996 30308
rect 10612 30280 11008 30308
rect 12268 30308 12296 30339
rect 12342 30336 12348 30388
rect 12400 30376 12406 30388
rect 12400 30348 12757 30376
rect 12400 30336 12406 30348
rect 12268 30280 12664 30308
rect 5077 30243 5135 30249
rect 5077 30209 5089 30243
rect 5123 30209 5135 30243
rect 5537 30243 5595 30249
rect 5537 30240 5549 30243
rect 5077 30203 5135 30209
rect 5368 30212 5549 30240
rect 5368 30184 5396 30212
rect 5537 30209 5549 30212
rect 5583 30209 5595 30243
rect 5537 30203 5595 30209
rect 6178 30200 6184 30252
rect 6236 30240 6242 30252
rect 6641 30243 6699 30249
rect 6641 30240 6653 30243
rect 6236 30212 6653 30240
rect 6236 30200 6242 30212
rect 6641 30209 6653 30212
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30240 6791 30243
rect 6822 30240 6828 30252
rect 6779 30212 6828 30240
rect 6779 30209 6791 30212
rect 6733 30203 6791 30209
rect 5166 30132 5172 30184
rect 5224 30132 5230 30184
rect 5350 30132 5356 30184
rect 5408 30132 5414 30184
rect 6656 30172 6684 30203
rect 6822 30200 6828 30212
rect 6880 30240 6886 30252
rect 7009 30243 7067 30249
rect 7009 30240 7021 30243
rect 6880 30212 7021 30240
rect 6880 30200 6886 30212
rect 7009 30209 7021 30212
rect 7055 30209 7067 30243
rect 7009 30203 7067 30209
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 7469 30243 7527 30249
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 7742 30240 7748 30252
rect 7515 30212 7748 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 7208 30172 7236 30203
rect 7742 30200 7748 30212
rect 7800 30240 7806 30252
rect 8389 30243 8447 30249
rect 7800 30212 8248 30240
rect 7800 30200 7806 30212
rect 8220 30184 8248 30212
rect 8389 30209 8401 30243
rect 8435 30209 8447 30243
rect 8389 30203 8447 30209
rect 8481 30243 8539 30249
rect 8481 30209 8493 30243
rect 8527 30209 8539 30243
rect 8481 30203 8539 30209
rect 5460 30144 5764 30172
rect 6656 30144 7236 30172
rect 5460 30104 5488 30144
rect 4724 30076 5488 30104
rect 5534 30064 5540 30116
rect 5592 30104 5598 30116
rect 5629 30107 5687 30113
rect 5629 30104 5641 30107
rect 5592 30076 5641 30104
rect 5592 30064 5598 30076
rect 5629 30073 5641 30076
rect 5675 30073 5687 30107
rect 5736 30104 5764 30144
rect 7558 30132 7564 30184
rect 7616 30172 7622 30184
rect 8110 30172 8116 30184
rect 7616 30144 8116 30172
rect 7616 30132 7622 30144
rect 8110 30132 8116 30144
rect 8168 30132 8174 30184
rect 8202 30132 8208 30184
rect 8260 30132 8266 30184
rect 8404 30104 8432 30203
rect 8496 30172 8524 30203
rect 8662 30200 8668 30252
rect 8720 30200 8726 30252
rect 8772 30249 8800 30280
rect 9968 30252 9996 30280
rect 8757 30243 8815 30249
rect 8757 30209 8769 30243
rect 8803 30209 8815 30243
rect 8757 30203 8815 30209
rect 9033 30243 9091 30249
rect 9033 30209 9045 30243
rect 9079 30240 9091 30243
rect 9214 30240 9220 30252
rect 9079 30212 9220 30240
rect 9079 30209 9091 30212
rect 9033 30203 9091 30209
rect 9048 30172 9076 30203
rect 9214 30200 9220 30212
rect 9272 30200 9278 30252
rect 9950 30200 9956 30252
rect 10008 30200 10014 30252
rect 10410 30200 10416 30252
rect 10468 30240 10474 30252
rect 10505 30243 10563 30249
rect 10505 30240 10517 30243
rect 10468 30212 10517 30240
rect 10468 30200 10474 30212
rect 10505 30209 10517 30212
rect 10551 30240 10563 30243
rect 10870 30240 10876 30252
rect 10551 30212 10876 30240
rect 10551 30209 10563 30212
rect 10505 30203 10563 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 11330 30200 11336 30252
rect 11388 30200 11394 30252
rect 11514 30200 11520 30252
rect 11572 30200 11578 30252
rect 11606 30200 11612 30252
rect 11664 30200 11670 30252
rect 11974 30200 11980 30252
rect 12032 30240 12038 30252
rect 12636 30249 12664 30280
rect 12729 30249 12757 30348
rect 12986 30336 12992 30388
rect 13044 30336 13050 30388
rect 13998 30376 14004 30388
rect 13464 30348 14004 30376
rect 12161 30243 12219 30249
rect 12161 30240 12173 30243
rect 12032 30212 12173 30240
rect 12032 30200 12038 30212
rect 12161 30209 12173 30212
rect 12207 30209 12219 30243
rect 12161 30203 12219 30209
rect 12345 30243 12403 30249
rect 12345 30209 12357 30243
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 12621 30243 12679 30249
rect 12621 30209 12633 30243
rect 12667 30209 12679 30243
rect 12621 30203 12679 30209
rect 12714 30243 12772 30249
rect 12714 30209 12726 30243
rect 12760 30209 12772 30243
rect 12714 30203 12772 30209
rect 8496 30144 9076 30172
rect 9125 30175 9183 30181
rect 9125 30141 9137 30175
rect 9171 30141 9183 30175
rect 9125 30135 9183 30141
rect 9140 30104 9168 30135
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9401 30175 9459 30181
rect 9401 30172 9413 30175
rect 9364 30144 9413 30172
rect 9364 30132 9370 30144
rect 9401 30141 9413 30144
rect 9447 30141 9459 30175
rect 9401 30135 9459 30141
rect 9490 30132 9496 30184
rect 9548 30132 9554 30184
rect 10597 30175 10655 30181
rect 10597 30141 10609 30175
rect 10643 30172 10655 30175
rect 11885 30175 11943 30181
rect 11885 30172 11897 30175
rect 10643 30144 11897 30172
rect 10643 30141 10655 30144
rect 10597 30135 10655 30141
rect 11885 30141 11897 30144
rect 11931 30141 11943 30175
rect 11885 30135 11943 30141
rect 9508 30104 9536 30132
rect 11330 30104 11336 30116
rect 5736 30076 8294 30104
rect 8404 30076 9536 30104
rect 11164 30076 11336 30104
rect 5629 30067 5687 30073
rect 2869 30039 2927 30045
rect 2869 30005 2881 30039
rect 2915 30036 2927 30039
rect 2958 30036 2964 30048
rect 2915 30008 2964 30036
rect 2915 30005 2927 30008
rect 2869 29999 2927 30005
rect 2958 29996 2964 30008
rect 3016 29996 3022 30048
rect 4154 29996 4160 30048
rect 4212 30036 4218 30048
rect 4985 30039 5043 30045
rect 4985 30036 4997 30039
rect 4212 30008 4997 30036
rect 4212 29996 4218 30008
rect 4985 30005 4997 30008
rect 5031 30005 5043 30039
rect 4985 29999 5043 30005
rect 5258 29996 5264 30048
rect 5316 29996 5322 30048
rect 5721 30039 5779 30045
rect 5721 30005 5733 30039
rect 5767 30036 5779 30039
rect 6362 30036 6368 30048
rect 5767 30008 6368 30036
rect 5767 30005 5779 30008
rect 5721 29999 5779 30005
rect 6362 29996 6368 30008
rect 6420 29996 6426 30048
rect 7650 29996 7656 30048
rect 7708 29996 7714 30048
rect 8266 30036 8294 30076
rect 11164 30036 11192 30076
rect 11330 30064 11336 30076
rect 11388 30064 11394 30116
rect 8266 30008 11192 30036
rect 12250 29996 12256 30048
rect 12308 30036 12314 30048
rect 12360 30036 12388 30203
rect 12434 30132 12440 30184
rect 12492 30172 12498 30184
rect 13464 30172 13492 30348
rect 13998 30336 14004 30348
rect 14056 30336 14062 30388
rect 14274 30336 14280 30388
rect 14332 30336 14338 30388
rect 15105 30379 15163 30385
rect 15105 30345 15117 30379
rect 15151 30376 15163 30379
rect 15654 30376 15660 30388
rect 15151 30348 15660 30376
rect 15151 30345 15163 30348
rect 15105 30339 15163 30345
rect 15654 30336 15660 30348
rect 15712 30336 15718 30388
rect 16485 30379 16543 30385
rect 16485 30345 16497 30379
rect 16531 30376 16543 30379
rect 17770 30376 17776 30388
rect 16531 30348 17776 30376
rect 16531 30345 16543 30348
rect 16485 30339 16543 30345
rect 17770 30336 17776 30348
rect 17828 30376 17834 30388
rect 17828 30348 19380 30376
rect 17828 30336 17834 30348
rect 14826 30308 14832 30320
rect 13556 30280 14832 30308
rect 13556 30249 13584 30280
rect 14826 30268 14832 30280
rect 14884 30268 14890 30320
rect 16206 30308 16212 30320
rect 16132 30280 16212 30308
rect 13541 30243 13599 30249
rect 13541 30209 13553 30243
rect 13587 30209 13599 30243
rect 13541 30203 13599 30209
rect 13725 30243 13783 30249
rect 13725 30209 13737 30243
rect 13771 30240 13783 30243
rect 14093 30243 14151 30249
rect 13771 30212 14044 30240
rect 13771 30209 13783 30212
rect 13725 30203 13783 30209
rect 13909 30175 13967 30181
rect 13909 30172 13921 30175
rect 12492 30144 13124 30172
rect 13464 30144 13921 30172
rect 12492 30132 12498 30144
rect 13096 30116 13124 30144
rect 13909 30141 13921 30144
rect 13955 30141 13967 30175
rect 13909 30135 13967 30141
rect 12526 30064 12532 30116
rect 12584 30104 12590 30116
rect 12584 30076 12756 30104
rect 12584 30064 12590 30076
rect 12618 30036 12624 30048
rect 12308 30008 12624 30036
rect 12308 29996 12314 30008
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 12728 30036 12756 30076
rect 13078 30064 13084 30116
rect 13136 30064 13142 30116
rect 13265 30107 13323 30113
rect 13265 30073 13277 30107
rect 13311 30104 13323 30107
rect 14016 30104 14044 30212
rect 14093 30209 14105 30243
rect 14139 30240 14151 30243
rect 15013 30243 15071 30249
rect 15013 30240 15025 30243
rect 14139 30212 15025 30240
rect 14139 30209 14151 30212
rect 14093 30203 14151 30209
rect 15013 30209 15025 30212
rect 15059 30209 15071 30243
rect 15013 30203 15071 30209
rect 15102 30200 15108 30252
rect 15160 30200 15166 30252
rect 15470 30200 15476 30252
rect 15528 30200 15534 30252
rect 15654 30200 15660 30252
rect 15712 30240 15718 30252
rect 15930 30240 15936 30252
rect 15712 30212 15936 30240
rect 15712 30200 15718 30212
rect 15930 30200 15936 30212
rect 15988 30200 15994 30252
rect 16132 30249 16160 30280
rect 16206 30268 16212 30280
rect 16264 30268 16270 30320
rect 16942 30268 16948 30320
rect 17000 30268 17006 30320
rect 17052 30280 17540 30308
rect 17052 30249 17080 30280
rect 17512 30252 17540 30280
rect 18598 30268 18604 30320
rect 18656 30308 18662 30320
rect 19352 30308 19380 30348
rect 20714 30336 20720 30388
rect 20772 30376 20778 30388
rect 21177 30379 21235 30385
rect 21177 30376 21189 30379
rect 20772 30348 21189 30376
rect 20772 30336 20778 30348
rect 21177 30345 21189 30348
rect 21223 30345 21235 30379
rect 21177 30339 21235 30345
rect 21821 30379 21879 30385
rect 21821 30345 21833 30379
rect 21867 30376 21879 30379
rect 22002 30376 22008 30388
rect 21867 30348 22008 30376
rect 21867 30345 21879 30348
rect 21821 30339 21879 30345
rect 22002 30336 22008 30348
rect 22060 30336 22066 30388
rect 22922 30376 22928 30388
rect 22848 30348 22928 30376
rect 20346 30308 20352 30320
rect 18656 30280 19288 30308
rect 19352 30280 20352 30308
rect 18656 30268 18662 30280
rect 16117 30243 16175 30249
rect 16117 30209 16129 30243
rect 16163 30209 16175 30243
rect 16669 30243 16727 30249
rect 16669 30240 16681 30243
rect 16117 30203 16175 30209
rect 16224 30212 16681 30240
rect 14182 30132 14188 30184
rect 14240 30172 14246 30184
rect 14461 30175 14519 30181
rect 14240 30144 14412 30172
rect 14240 30132 14246 30144
rect 14274 30104 14280 30116
rect 13311 30076 13952 30104
rect 14016 30076 14280 30104
rect 13311 30073 13323 30076
rect 13265 30067 13323 30073
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 12728 30008 13553 30036
rect 13541 30005 13553 30008
rect 13587 30005 13599 30039
rect 13924 30036 13952 30076
rect 14274 30064 14280 30076
rect 14332 30064 14338 30116
rect 14384 30104 14412 30144
rect 14461 30141 14473 30175
rect 14507 30172 14519 30175
rect 15120 30172 15148 30200
rect 14507 30144 15148 30172
rect 14507 30141 14519 30144
rect 14461 30135 14519 30141
rect 15194 30132 15200 30184
rect 15252 30172 15258 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 15252 30144 15577 30172
rect 15252 30132 15258 30144
rect 15565 30141 15577 30144
rect 15611 30141 15623 30175
rect 15565 30135 15623 30141
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30172 15807 30175
rect 16025 30175 16083 30181
rect 16025 30172 16037 30175
rect 15795 30144 16037 30172
rect 15795 30141 15807 30144
rect 15749 30135 15807 30141
rect 16025 30141 16037 30144
rect 16071 30141 16083 30175
rect 16025 30135 16083 30141
rect 16132 30104 16160 30203
rect 16224 30184 16252 30212
rect 16669 30209 16681 30212
rect 16715 30209 16727 30243
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16669 30203 16727 30209
rect 16776 30212 16865 30240
rect 16206 30132 16212 30184
rect 16264 30132 16270 30184
rect 16482 30132 16488 30184
rect 16540 30172 16546 30184
rect 16776 30172 16804 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 17037 30243 17095 30249
rect 17037 30209 17049 30243
rect 17083 30209 17095 30243
rect 17037 30203 17095 30209
rect 17126 30200 17132 30252
rect 17184 30200 17190 30252
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 16540 30144 16804 30172
rect 17144 30172 17172 30200
rect 17328 30172 17356 30203
rect 17494 30200 17500 30252
rect 17552 30200 17558 30252
rect 17586 30200 17592 30252
rect 17644 30200 17650 30252
rect 17865 30243 17923 30249
rect 17865 30209 17877 30243
rect 17911 30209 17923 30243
rect 17865 30203 17923 30209
rect 17144 30144 17356 30172
rect 17681 30175 17739 30181
rect 16540 30132 16546 30144
rect 17681 30141 17693 30175
rect 17727 30141 17739 30175
rect 17681 30135 17739 30141
rect 14384 30076 16160 30104
rect 17126 30064 17132 30116
rect 17184 30104 17190 30116
rect 17696 30104 17724 30135
rect 17184 30076 17724 30104
rect 17184 30064 17190 30076
rect 13998 30036 14004 30048
rect 13924 30008 14004 30036
rect 13541 29999 13599 30005
rect 13998 29996 14004 30008
rect 14056 29996 14062 30048
rect 17218 29996 17224 30048
rect 17276 29996 17282 30048
rect 17678 29996 17684 30048
rect 17736 30036 17742 30048
rect 17880 30036 17908 30203
rect 17954 30200 17960 30252
rect 18012 30240 18018 30252
rect 18049 30243 18107 30249
rect 18049 30240 18061 30243
rect 18012 30212 18061 30240
rect 18012 30200 18018 30212
rect 18049 30209 18061 30212
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30209 19119 30243
rect 19260 30243 19288 30280
rect 19536 30249 19564 30280
rect 20346 30268 20352 30280
rect 20404 30268 20410 30320
rect 20438 30268 20444 30320
rect 20496 30308 20502 30320
rect 21453 30311 21511 30317
rect 21453 30308 21465 30311
rect 20496 30280 21465 30308
rect 20496 30268 20502 30280
rect 21453 30277 21465 30280
rect 21499 30277 21511 30311
rect 21453 30271 21511 30277
rect 21637 30311 21695 30317
rect 21637 30277 21649 30311
rect 21683 30308 21695 30311
rect 22848 30308 22876 30348
rect 22922 30336 22928 30348
rect 22980 30336 22986 30388
rect 23474 30376 23480 30388
rect 23216 30348 23480 30376
rect 23216 30317 23244 30348
rect 23474 30336 23480 30348
rect 23532 30336 23538 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 23992 30348 24532 30376
rect 23992 30336 23998 30348
rect 24504 30317 24532 30348
rect 25130 30336 25136 30388
rect 25188 30376 25194 30388
rect 25188 30348 26372 30376
rect 25188 30336 25194 30348
rect 23201 30311 23259 30317
rect 21683 30280 22324 30308
rect 22848 30280 23051 30308
rect 21683 30277 21695 30280
rect 21637 30271 21695 30277
rect 19337 30243 19395 30249
rect 19260 30215 19349 30243
rect 19061 30203 19119 30209
rect 19337 30209 19349 30215
rect 19383 30209 19395 30243
rect 19337 30203 19395 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 20064 30243 20122 30249
rect 20064 30209 20076 30243
rect 20110 30240 20122 30243
rect 21082 30240 21088 30252
rect 20110 30212 21088 30240
rect 20110 30209 20122 30212
rect 20064 30203 20122 30209
rect 18325 30175 18383 30181
rect 18325 30141 18337 30175
rect 18371 30141 18383 30175
rect 18325 30135 18383 30141
rect 18340 30048 18368 30135
rect 19076 30116 19104 30203
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 21358 30240 21364 30252
rect 21315 30212 21364 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 19306 30144 19656 30172
rect 19058 30064 19064 30116
rect 19116 30064 19122 30116
rect 19150 30064 19156 30116
rect 19208 30104 19214 30116
rect 19306 30104 19334 30144
rect 19208 30076 19334 30104
rect 19429 30107 19487 30113
rect 19208 30064 19214 30076
rect 19429 30073 19441 30107
rect 19475 30104 19487 30107
rect 19518 30104 19524 30116
rect 19475 30076 19524 30104
rect 19475 30073 19487 30076
rect 19429 30067 19487 30073
rect 19518 30064 19524 30076
rect 19576 30064 19582 30116
rect 17736 30008 17908 30036
rect 17736 29996 17742 30008
rect 18322 29996 18328 30048
rect 18380 29996 18386 30048
rect 18874 29996 18880 30048
rect 18932 29996 18938 30048
rect 19245 30039 19303 30045
rect 19245 30005 19257 30039
rect 19291 30036 19303 30039
rect 19334 30036 19340 30048
rect 19291 30008 19340 30036
rect 19291 30005 19303 30008
rect 19245 29999 19303 30005
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 19628 30036 19656 30144
rect 19794 30132 19800 30184
rect 19852 30132 19858 30184
rect 20806 30132 20812 30184
rect 20864 30172 20870 30184
rect 21284 30172 21312 30203
rect 21358 30200 21364 30212
rect 21416 30200 21422 30252
rect 20864 30144 21312 30172
rect 21468 30172 21496 30271
rect 22296 30249 22324 30280
rect 22097 30243 22155 30249
rect 22097 30209 22109 30243
rect 22143 30209 22155 30243
rect 22097 30203 22155 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 22281 30243 22339 30249
rect 22281 30209 22293 30243
rect 22327 30209 22339 30243
rect 22281 30203 22339 30209
rect 21634 30172 21640 30184
rect 21468 30144 21640 30172
rect 20864 30132 20870 30144
rect 21634 30132 21640 30144
rect 21692 30132 21698 30184
rect 20990 30064 20996 30116
rect 21048 30104 21054 30116
rect 22112 30104 22140 30203
rect 22204 30172 22232 30203
rect 22462 30200 22468 30252
rect 22520 30200 22526 30252
rect 22925 30243 22983 30249
rect 22925 30209 22937 30243
rect 22971 30209 22983 30243
rect 23023 30243 23051 30280
rect 23201 30277 23213 30311
rect 23247 30277 23259 30311
rect 24213 30311 24271 30317
rect 24213 30308 24225 30311
rect 23201 30271 23259 30277
rect 23492 30280 24225 30308
rect 23109 30243 23167 30249
rect 23023 30215 23121 30243
rect 22925 30203 22983 30209
rect 23109 30209 23121 30215
rect 23155 30209 23167 30243
rect 23109 30203 23167 30209
rect 22370 30172 22376 30184
rect 22204 30144 22376 30172
rect 22370 30132 22376 30144
rect 22428 30132 22434 30184
rect 22940 30172 22968 30203
rect 23290 30200 23296 30252
rect 23348 30200 23354 30252
rect 23492 30240 23520 30280
rect 24213 30277 24225 30280
rect 24259 30277 24271 30311
rect 24213 30271 24271 30277
rect 24489 30311 24547 30317
rect 24489 30277 24501 30311
rect 24535 30308 24547 30311
rect 24578 30308 24584 30320
rect 24535 30280 24584 30308
rect 24535 30277 24547 30280
rect 24489 30271 24547 30277
rect 24578 30268 24584 30280
rect 24636 30268 24642 30320
rect 25424 30280 25912 30308
rect 25424 30252 25452 30280
rect 23400 30212 23520 30240
rect 23569 30243 23627 30249
rect 23400 30172 23428 30212
rect 23569 30209 23581 30243
rect 23615 30240 23627 30243
rect 23658 30240 23664 30252
rect 23615 30212 23664 30240
rect 23615 30209 23627 30212
rect 23569 30203 23627 30209
rect 23658 30200 23664 30212
rect 23716 30200 23722 30252
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 22940 30144 23428 30172
rect 23474 30132 23480 30184
rect 23532 30132 23538 30184
rect 23842 30132 23848 30184
rect 23900 30132 23906 30184
rect 23952 30172 23980 30203
rect 24026 30200 24032 30252
rect 24084 30200 24090 30252
rect 24673 30243 24731 30249
rect 24673 30209 24685 30243
rect 24719 30240 24731 30243
rect 24762 30240 24768 30252
rect 24719 30212 24768 30240
rect 24719 30209 24731 30212
rect 24673 30203 24731 30209
rect 24762 30200 24768 30212
rect 24820 30200 24826 30252
rect 25314 30200 25320 30252
rect 25372 30200 25378 30252
rect 25406 30200 25412 30252
rect 25464 30200 25470 30252
rect 25498 30200 25504 30252
rect 25556 30200 25562 30252
rect 25590 30200 25596 30252
rect 25648 30200 25654 30252
rect 25774 30200 25780 30252
rect 25832 30200 25838 30252
rect 25884 30240 25912 30280
rect 26344 30249 26372 30348
rect 26528 30348 26924 30376
rect 26528 30252 26556 30348
rect 26053 30243 26111 30249
rect 26053 30240 26065 30243
rect 25884 30212 26065 30240
rect 26053 30209 26065 30212
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 26329 30243 26387 30249
rect 26329 30209 26341 30243
rect 26375 30209 26387 30243
rect 26329 30203 26387 30209
rect 26510 30200 26516 30252
rect 26568 30200 26574 30252
rect 26697 30243 26755 30249
rect 26697 30209 26709 30243
rect 26743 30240 26755 30243
rect 26786 30240 26792 30252
rect 26743 30212 26792 30240
rect 26743 30209 26755 30212
rect 26697 30203 26755 30209
rect 26786 30200 26792 30212
rect 26844 30200 26850 30252
rect 26896 30240 26924 30348
rect 27706 30336 27712 30388
rect 27764 30376 27770 30388
rect 28166 30376 28172 30388
rect 27764 30348 28172 30376
rect 27764 30336 27770 30348
rect 28166 30336 28172 30348
rect 28224 30376 28230 30388
rect 28810 30376 28816 30388
rect 28224 30348 28816 30376
rect 28224 30336 28230 30348
rect 28810 30336 28816 30348
rect 28868 30336 28874 30388
rect 29270 30336 29276 30388
rect 29328 30376 29334 30388
rect 29549 30379 29607 30385
rect 29328 30348 29500 30376
rect 29328 30336 29334 30348
rect 26973 30311 27031 30317
rect 26973 30277 26985 30311
rect 27019 30308 27031 30311
rect 28074 30308 28080 30320
rect 27019 30280 28080 30308
rect 27019 30277 27031 30280
rect 26973 30271 27031 30277
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 26896 30212 27353 30240
rect 27341 30209 27353 30212
rect 27387 30240 27399 30243
rect 27430 30240 27436 30252
rect 27387 30212 27436 30240
rect 27387 30209 27399 30212
rect 27341 30203 27399 30209
rect 27430 30200 27436 30212
rect 27488 30200 27494 30252
rect 28000 30249 28028 30280
rect 28074 30268 28080 30280
rect 28132 30268 28138 30320
rect 28534 30268 28540 30320
rect 28592 30308 28598 30320
rect 29472 30308 29500 30348
rect 29549 30345 29561 30379
rect 29595 30376 29607 30379
rect 29595 30348 30236 30376
rect 29595 30345 29607 30348
rect 29549 30339 29607 30345
rect 30208 30320 30236 30348
rect 30282 30336 30288 30388
rect 30340 30376 30346 30388
rect 30742 30376 30748 30388
rect 30340 30348 30748 30376
rect 30340 30336 30346 30348
rect 30742 30336 30748 30348
rect 30800 30336 30806 30388
rect 33502 30336 33508 30388
rect 33560 30336 33566 30388
rect 28592 30280 29132 30308
rect 29472 30280 29684 30308
rect 28592 30268 28598 30280
rect 27985 30243 28043 30249
rect 27985 30209 27997 30243
rect 28031 30209 28043 30243
rect 27985 30203 28043 30209
rect 28445 30243 28503 30249
rect 28445 30209 28457 30243
rect 28491 30238 28503 30243
rect 28552 30238 28580 30268
rect 28491 30210 28580 30238
rect 28629 30243 28687 30249
rect 28491 30209 28503 30210
rect 28445 30203 28503 30209
rect 28629 30209 28641 30243
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 24118 30172 24124 30184
rect 23952 30144 24124 30172
rect 24118 30132 24124 30144
rect 24176 30132 24182 30184
rect 24213 30175 24271 30181
rect 24213 30141 24225 30175
rect 24259 30141 24271 30175
rect 24213 30135 24271 30141
rect 24949 30175 25007 30181
rect 24949 30141 24961 30175
rect 24995 30172 25007 30175
rect 25682 30172 25688 30184
rect 24995 30144 25688 30172
rect 24995 30141 25007 30144
rect 24949 30135 25007 30141
rect 22186 30104 22192 30116
rect 21048 30076 22192 30104
rect 21048 30064 21054 30076
rect 22186 30064 22192 30076
rect 22244 30104 22250 30116
rect 23290 30104 23296 30116
rect 22244 30076 23296 30104
rect 22244 30064 22250 30076
rect 23290 30064 23296 30076
rect 23348 30064 23354 30116
rect 23492 30104 23520 30132
rect 24228 30104 24256 30135
rect 25682 30132 25688 30144
rect 25740 30132 25746 30184
rect 26145 30175 26203 30181
rect 26145 30141 26157 30175
rect 26191 30172 26203 30175
rect 28261 30175 28319 30181
rect 28261 30172 28273 30175
rect 26191 30144 28273 30172
rect 26191 30141 26203 30144
rect 26145 30135 26203 30141
rect 28261 30141 28273 30144
rect 28307 30172 28319 30175
rect 28350 30172 28356 30184
rect 28307 30144 28356 30172
rect 28307 30141 28319 30144
rect 28261 30135 28319 30141
rect 28350 30132 28356 30144
rect 28408 30172 28414 30184
rect 28644 30172 28672 30203
rect 28810 30200 28816 30252
rect 28868 30200 28874 30252
rect 28902 30200 28908 30252
rect 28960 30240 28966 30252
rect 29104 30249 29132 30280
rect 28997 30243 29055 30249
rect 28997 30240 29009 30243
rect 28960 30212 29009 30240
rect 28960 30200 28966 30212
rect 28997 30209 29009 30212
rect 29043 30209 29055 30243
rect 28997 30203 29055 30209
rect 29089 30243 29147 30249
rect 29089 30209 29101 30243
rect 29135 30209 29147 30243
rect 29089 30203 29147 30209
rect 29178 30200 29184 30252
rect 29236 30200 29242 30252
rect 29454 30200 29460 30252
rect 29512 30200 29518 30252
rect 29656 30249 29684 30280
rect 29748 30280 30144 30308
rect 29748 30249 29776 30280
rect 29641 30243 29699 30249
rect 29641 30209 29653 30243
rect 29687 30209 29699 30243
rect 29641 30203 29699 30209
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30209 29791 30243
rect 29733 30203 29791 30209
rect 30009 30243 30067 30249
rect 30009 30209 30021 30243
rect 30055 30209 30067 30243
rect 30116 30240 30144 30280
rect 30190 30268 30196 30320
rect 30248 30268 30254 30320
rect 30466 30268 30472 30320
rect 30524 30308 30530 30320
rect 31018 30308 31024 30320
rect 30524 30280 31024 30308
rect 30524 30268 30530 30280
rect 31018 30268 31024 30280
rect 31076 30268 31082 30320
rect 31665 30311 31723 30317
rect 31665 30308 31677 30311
rect 31119 30280 31677 30308
rect 30285 30243 30343 30249
rect 30116 30212 30236 30240
rect 30009 30203 30067 30209
rect 28408 30144 28672 30172
rect 28828 30172 28856 30200
rect 29273 30175 29331 30181
rect 29273 30172 29285 30175
rect 28828 30144 29285 30172
rect 28408 30132 28414 30144
rect 29273 30141 29285 30144
rect 29319 30141 29331 30175
rect 29273 30135 29331 30141
rect 23492 30076 25259 30104
rect 20070 30036 20076 30048
rect 19628 30008 20076 30036
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 22646 29996 22652 30048
rect 22704 30036 22710 30048
rect 22741 30039 22799 30045
rect 22741 30036 22753 30039
rect 22704 30008 22753 30036
rect 22704 29996 22710 30008
rect 22741 30005 22753 30008
rect 22787 30005 22799 30039
rect 22741 29999 22799 30005
rect 23474 29996 23480 30048
rect 23532 29996 23538 30048
rect 23658 29996 23664 30048
rect 23716 29996 23722 30048
rect 23750 29996 23756 30048
rect 23808 29996 23814 30048
rect 23842 29996 23848 30048
rect 23900 30036 23906 30048
rect 24302 30036 24308 30048
rect 23900 30008 24308 30036
rect 23900 29996 23906 30008
rect 24302 29996 24308 30008
rect 24360 29996 24366 30048
rect 24857 30039 24915 30045
rect 24857 30005 24869 30039
rect 24903 30036 24915 30039
rect 25133 30039 25191 30045
rect 25133 30036 25145 30039
rect 24903 30008 25145 30036
rect 24903 30005 24915 30008
rect 24857 29999 24915 30005
rect 25133 30005 25145 30008
rect 25179 30005 25191 30039
rect 25231 30036 25259 30076
rect 25406 30064 25412 30116
rect 25464 30064 25470 30116
rect 25774 30064 25780 30116
rect 25832 30064 25838 30116
rect 26234 30064 26240 30116
rect 26292 30064 26298 30116
rect 26878 30064 26884 30116
rect 26936 30104 26942 30116
rect 27249 30107 27307 30113
rect 27249 30104 27261 30107
rect 26936 30076 27261 30104
rect 26936 30064 26942 30076
rect 27249 30073 27261 30076
rect 27295 30073 27307 30107
rect 27249 30067 27307 30073
rect 28813 30107 28871 30113
rect 28813 30073 28825 30107
rect 28859 30104 28871 30107
rect 30024 30104 30052 30203
rect 28859 30076 30052 30104
rect 28859 30073 28871 30076
rect 28813 30067 28871 30073
rect 25792 30036 25820 30064
rect 25231 30008 25820 30036
rect 25869 30039 25927 30045
rect 25133 29999 25191 30005
rect 25869 30005 25881 30039
rect 25915 30036 25927 30039
rect 25958 30036 25964 30048
rect 25915 30008 25964 30036
rect 25915 30005 25927 30008
rect 25869 29999 25927 30005
rect 25958 29996 25964 30008
rect 26016 29996 26022 30048
rect 26050 29996 26056 30048
rect 26108 30036 26114 30048
rect 26605 30039 26663 30045
rect 26605 30036 26617 30039
rect 26108 30008 26617 30036
rect 26108 29996 26114 30008
rect 26605 30005 26617 30008
rect 26651 30005 26663 30039
rect 26605 29999 26663 30005
rect 26694 29996 26700 30048
rect 26752 30036 26758 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 26752 30008 26985 30036
rect 26752 29996 26758 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 26973 29999 27031 30005
rect 27062 29996 27068 30048
rect 27120 30036 27126 30048
rect 27157 30039 27215 30045
rect 27157 30036 27169 30039
rect 27120 30008 27169 30036
rect 27120 29996 27126 30008
rect 27157 30005 27169 30008
rect 27203 30005 27215 30039
rect 27157 29999 27215 30005
rect 27614 29996 27620 30048
rect 27672 30036 27678 30048
rect 27801 30039 27859 30045
rect 27801 30036 27813 30039
rect 27672 30008 27813 30036
rect 27672 29996 27678 30008
rect 27801 30005 27813 30008
rect 27847 30005 27859 30039
rect 27801 29999 27859 30005
rect 28169 30039 28227 30045
rect 28169 30005 28181 30039
rect 28215 30036 28227 30039
rect 28442 30036 28448 30048
rect 28215 30008 28448 30036
rect 28215 30005 28227 30008
rect 28169 29999 28227 30005
rect 28442 29996 28448 30008
rect 28500 29996 28506 30048
rect 28537 30039 28595 30045
rect 28537 30005 28549 30039
rect 28583 30036 28595 30039
rect 28626 30036 28632 30048
rect 28583 30008 28632 30036
rect 28583 30005 28595 30008
rect 28537 29999 28595 30005
rect 28626 29996 28632 30008
rect 28684 29996 28690 30048
rect 28718 29996 28724 30048
rect 28776 30036 28782 30048
rect 29825 30039 29883 30045
rect 29825 30036 29837 30039
rect 28776 30008 29837 30036
rect 28776 29996 28782 30008
rect 29825 30005 29837 30008
rect 29871 30005 29883 30039
rect 30208 30036 30236 30212
rect 30285 30209 30297 30243
rect 30331 30209 30343 30243
rect 30285 30203 30343 30209
rect 30377 30243 30435 30249
rect 30377 30209 30389 30243
rect 30423 30240 30435 30243
rect 30484 30240 30512 30268
rect 30423 30212 30512 30240
rect 30745 30243 30803 30249
rect 30423 30209 30435 30212
rect 30377 30203 30435 30209
rect 30745 30209 30757 30243
rect 30791 30240 30803 30243
rect 31119 30240 31147 30280
rect 31665 30277 31677 30280
rect 31711 30308 31723 30311
rect 31938 30308 31944 30320
rect 31711 30280 31944 30308
rect 31711 30277 31723 30280
rect 31665 30271 31723 30277
rect 31938 30268 31944 30280
rect 31996 30268 32002 30320
rect 30791 30212 31147 30240
rect 30791 30209 30803 30212
rect 30745 30203 30803 30209
rect 30300 30104 30328 30203
rect 30466 30132 30472 30184
rect 30524 30172 30530 30184
rect 30760 30172 30788 30203
rect 31386 30200 31392 30252
rect 31444 30200 31450 30252
rect 31570 30200 31576 30252
rect 31628 30200 31634 30252
rect 31754 30200 31760 30252
rect 31812 30200 31818 30252
rect 32214 30200 32220 30252
rect 32272 30240 32278 30252
rect 32381 30243 32439 30249
rect 32381 30240 32393 30243
rect 32272 30212 32393 30240
rect 32272 30200 32278 30212
rect 32381 30209 32393 30212
rect 32427 30209 32439 30243
rect 32381 30203 32439 30209
rect 30524 30144 30788 30172
rect 30524 30132 30530 30144
rect 30926 30132 30932 30184
rect 30984 30172 30990 30184
rect 32030 30172 32036 30184
rect 30984 30144 32036 30172
rect 30984 30132 30990 30144
rect 32030 30132 32036 30144
rect 32088 30172 32094 30184
rect 32125 30175 32183 30181
rect 32125 30172 32137 30175
rect 32088 30144 32137 30172
rect 32088 30132 32094 30144
rect 32125 30141 32137 30144
rect 32171 30141 32183 30175
rect 32125 30135 32183 30141
rect 30300 30076 32076 30104
rect 30466 30036 30472 30048
rect 30208 30008 30472 30036
rect 29825 29999 29883 30005
rect 30466 29996 30472 30008
rect 30524 29996 30530 30048
rect 30558 29996 30564 30048
rect 30616 29996 30622 30048
rect 30650 29996 30656 30048
rect 30708 30036 30714 30048
rect 31297 30039 31355 30045
rect 31297 30036 31309 30039
rect 30708 30008 31309 30036
rect 30708 29996 30714 30008
rect 31297 30005 31309 30008
rect 31343 30005 31355 30039
rect 31297 29999 31355 30005
rect 31938 29996 31944 30048
rect 31996 29996 32002 30048
rect 32048 30036 32076 30076
rect 32306 30036 32312 30048
rect 32048 30008 32312 30036
rect 32306 29996 32312 30008
rect 32364 29996 32370 30048
rect 1104 29946 43884 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 43884 29946
rect 1104 29872 43884 29894
rect 2498 29792 2504 29844
rect 2556 29832 2562 29844
rect 3145 29835 3203 29841
rect 3145 29832 3157 29835
rect 2556 29804 3157 29832
rect 2556 29792 2562 29804
rect 3145 29801 3157 29804
rect 3191 29832 3203 29835
rect 3234 29832 3240 29844
rect 3191 29804 3240 29832
rect 3191 29801 3203 29804
rect 3145 29795 3203 29801
rect 3234 29792 3240 29804
rect 3292 29792 3298 29844
rect 3418 29792 3424 29844
rect 3476 29832 3482 29844
rect 3513 29835 3571 29841
rect 3513 29832 3525 29835
rect 3476 29804 3525 29832
rect 3476 29792 3482 29804
rect 3513 29801 3525 29804
rect 3559 29801 3571 29835
rect 4433 29835 4491 29841
rect 4433 29832 4445 29835
rect 3513 29795 3571 29801
rect 4172 29804 4445 29832
rect 1578 29724 1584 29776
rect 1636 29764 1642 29776
rect 2958 29764 2964 29776
rect 1636 29736 2964 29764
rect 1636 29724 1642 29736
rect 2958 29724 2964 29736
rect 3016 29724 3022 29776
rect 1210 29656 1216 29708
rect 1268 29696 1274 29708
rect 1857 29699 1915 29705
rect 1857 29696 1869 29699
rect 1268 29668 1869 29696
rect 1268 29656 1274 29668
rect 1857 29665 1869 29668
rect 1903 29665 1915 29699
rect 1857 29659 1915 29665
rect 2682 29656 2688 29708
rect 2740 29696 2746 29708
rect 3053 29699 3111 29705
rect 3053 29696 3065 29699
rect 2740 29668 3065 29696
rect 2740 29656 2746 29668
rect 3053 29665 3065 29668
rect 3099 29665 3111 29699
rect 3053 29659 3111 29665
rect 3237 29669 3295 29675
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 2038 29628 2044 29640
rect 1627 29600 2044 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 2406 29588 2412 29640
rect 2464 29628 2470 29640
rect 2961 29631 3019 29637
rect 2961 29628 2973 29631
rect 2464 29600 2973 29628
rect 2464 29588 2470 29600
rect 2961 29597 2973 29600
rect 3007 29597 3019 29631
rect 3237 29635 3249 29669
rect 3283 29635 3295 29669
rect 3510 29656 3516 29708
rect 3568 29696 3574 29708
rect 3605 29699 3663 29705
rect 3605 29696 3617 29699
rect 3568 29668 3617 29696
rect 3568 29656 3574 29668
rect 3605 29665 3617 29668
rect 3651 29665 3663 29699
rect 3605 29659 3663 29665
rect 3881 29699 3939 29705
rect 3881 29665 3893 29699
rect 3927 29696 3939 29699
rect 3970 29696 3976 29708
rect 3927 29668 3976 29696
rect 3927 29665 3939 29668
rect 3881 29659 3939 29665
rect 3970 29656 3976 29668
rect 4028 29656 4034 29708
rect 3237 29629 3295 29635
rect 2961 29591 3019 29597
rect 1854 29452 1860 29504
rect 1912 29492 1918 29504
rect 2774 29492 2780 29504
rect 1912 29464 2780 29492
rect 1912 29452 1918 29464
rect 2774 29452 2780 29464
rect 2832 29452 2838 29504
rect 2976 29492 3004 29591
rect 3252 29560 3280 29629
rect 3326 29588 3332 29640
rect 3384 29588 3390 29640
rect 3418 29588 3424 29640
rect 3476 29588 3482 29640
rect 4065 29631 4123 29637
rect 4065 29597 4077 29631
rect 4111 29628 4123 29631
rect 4172 29628 4200 29804
rect 4433 29801 4445 29804
rect 4479 29801 4491 29835
rect 4433 29795 4491 29801
rect 4706 29792 4712 29844
rect 4764 29792 4770 29844
rect 5166 29792 5172 29844
rect 5224 29792 5230 29844
rect 6178 29792 6184 29844
rect 6236 29832 6242 29844
rect 6641 29835 6699 29841
rect 6236 29804 6597 29832
rect 6236 29792 6242 29804
rect 4249 29767 4307 29773
rect 4249 29733 4261 29767
rect 4295 29764 4307 29767
rect 5184 29764 5212 29792
rect 6454 29764 6460 29776
rect 4295 29736 5212 29764
rect 5552 29736 6460 29764
rect 4295 29733 4307 29736
rect 4249 29727 4307 29733
rect 4111 29600 4200 29628
rect 4111 29597 4123 29600
rect 4065 29591 4123 29597
rect 4264 29560 4292 29727
rect 5353 29699 5411 29705
rect 5353 29696 5365 29699
rect 4540 29668 5120 29696
rect 4540 29637 4568 29668
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29597 4583 29631
rect 4525 29591 4583 29597
rect 3252 29532 4292 29560
rect 4356 29560 4384 29591
rect 4706 29588 4712 29640
rect 4764 29588 4770 29640
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29597 4951 29631
rect 4893 29591 4951 29597
rect 4985 29631 5043 29637
rect 4985 29597 4997 29631
rect 5031 29597 5043 29631
rect 4985 29591 5043 29597
rect 4724 29560 4752 29588
rect 4356 29532 4752 29560
rect 4908 29504 4936 29591
rect 3970 29492 3976 29504
rect 2976 29464 3976 29492
rect 3970 29452 3976 29464
rect 4028 29452 4034 29504
rect 4890 29452 4896 29504
rect 4948 29452 4954 29504
rect 5000 29492 5028 29591
rect 5092 29572 5120 29668
rect 5184 29668 5365 29696
rect 5184 29637 5212 29668
rect 5353 29665 5365 29668
rect 5399 29665 5411 29699
rect 5353 29659 5411 29665
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29597 5227 29631
rect 5169 29591 5227 29597
rect 5258 29588 5264 29640
rect 5316 29588 5322 29640
rect 5552 29637 5580 29736
rect 6454 29724 6460 29736
rect 6512 29724 6518 29776
rect 6569 29764 6597 29804
rect 6641 29801 6653 29835
rect 6687 29832 6699 29835
rect 6822 29832 6828 29844
rect 6687 29804 6828 29832
rect 6687 29801 6699 29804
rect 6641 29795 6699 29801
rect 6822 29792 6828 29804
rect 6880 29792 6886 29844
rect 7653 29835 7711 29841
rect 7653 29832 7665 29835
rect 6932 29804 7665 29832
rect 6932 29764 6960 29804
rect 7653 29801 7665 29804
rect 7699 29801 7711 29835
rect 7653 29795 7711 29801
rect 8202 29792 8208 29844
rect 8260 29792 8266 29844
rect 8570 29792 8576 29844
rect 8628 29792 8634 29844
rect 8662 29792 8668 29844
rect 8720 29792 8726 29844
rect 9214 29792 9220 29844
rect 9272 29832 9278 29844
rect 9309 29835 9367 29841
rect 9309 29832 9321 29835
rect 9272 29804 9321 29832
rect 9272 29792 9278 29804
rect 9309 29801 9321 29804
rect 9355 29801 9367 29835
rect 9309 29795 9367 29801
rect 9953 29835 10011 29841
rect 9953 29801 9965 29835
rect 9999 29832 10011 29835
rect 10502 29832 10508 29844
rect 9999 29804 10508 29832
rect 9999 29801 10011 29804
rect 9953 29795 10011 29801
rect 10502 29792 10508 29804
rect 10560 29832 10566 29844
rect 11606 29832 11612 29844
rect 10560 29804 11612 29832
rect 10560 29792 10566 29804
rect 11606 29792 11612 29804
rect 11664 29792 11670 29844
rect 11701 29835 11759 29841
rect 11701 29801 11713 29835
rect 11747 29832 11759 29835
rect 11882 29832 11888 29844
rect 11747 29804 11888 29832
rect 11747 29801 11759 29804
rect 11701 29795 11759 29801
rect 11882 29792 11888 29804
rect 11940 29792 11946 29844
rect 12434 29792 12440 29844
rect 12492 29792 12498 29844
rect 13998 29792 14004 29844
rect 14056 29832 14062 29844
rect 16206 29832 16212 29844
rect 14056 29804 16212 29832
rect 14056 29792 14062 29804
rect 16206 29792 16212 29804
rect 16264 29792 16270 29844
rect 17218 29792 17224 29844
rect 17276 29792 17282 29844
rect 19058 29792 19064 29844
rect 19116 29832 19122 29844
rect 20625 29835 20683 29841
rect 20625 29832 20637 29835
rect 19116 29804 20637 29832
rect 19116 29792 19122 29804
rect 20625 29801 20637 29804
rect 20671 29801 20683 29835
rect 20625 29795 20683 29801
rect 21082 29792 21088 29844
rect 21140 29832 21146 29844
rect 22097 29835 22155 29841
rect 22097 29832 22109 29835
rect 21140 29804 22109 29832
rect 21140 29792 21146 29804
rect 22097 29801 22109 29804
rect 22143 29801 22155 29835
rect 22097 29795 22155 29801
rect 22186 29792 22192 29844
rect 22244 29832 22250 29844
rect 22738 29832 22744 29844
rect 22244 29804 22744 29832
rect 22244 29792 22250 29804
rect 22738 29792 22744 29804
rect 22796 29792 22802 29844
rect 23658 29792 23664 29844
rect 23716 29832 23722 29844
rect 24397 29835 24455 29841
rect 24397 29832 24409 29835
rect 23716 29804 24409 29832
rect 23716 29792 23722 29804
rect 24397 29801 24409 29804
rect 24443 29801 24455 29835
rect 24397 29795 24455 29801
rect 24765 29835 24823 29841
rect 24765 29801 24777 29835
rect 24811 29832 24823 29835
rect 25130 29832 25136 29844
rect 24811 29804 25136 29832
rect 24811 29801 24823 29804
rect 24765 29795 24823 29801
rect 25130 29792 25136 29804
rect 25188 29792 25194 29844
rect 25222 29792 25228 29844
rect 25280 29792 25286 29844
rect 25774 29792 25780 29844
rect 25832 29832 25838 29844
rect 26605 29835 26663 29841
rect 26605 29832 26617 29835
rect 25832 29804 26617 29832
rect 25832 29792 25838 29804
rect 26605 29801 26617 29804
rect 26651 29801 26663 29835
rect 26605 29795 26663 29801
rect 26786 29792 26792 29844
rect 26844 29832 26850 29844
rect 27430 29832 27436 29844
rect 26844 29804 27436 29832
rect 26844 29792 26850 29804
rect 27430 29792 27436 29804
rect 27488 29792 27494 29844
rect 27706 29792 27712 29844
rect 27764 29792 27770 29844
rect 27798 29792 27804 29844
rect 27856 29792 27862 29844
rect 28258 29792 28264 29844
rect 28316 29832 28322 29844
rect 28810 29832 28816 29844
rect 28316 29804 28816 29832
rect 28316 29792 28322 29804
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 29086 29792 29092 29844
rect 29144 29792 29150 29844
rect 30558 29792 30564 29844
rect 30616 29792 30622 29844
rect 30929 29835 30987 29841
rect 30929 29801 30941 29835
rect 30975 29832 30987 29835
rect 30975 29804 31754 29832
rect 30975 29801 30987 29804
rect 30929 29795 30987 29801
rect 6569 29736 6960 29764
rect 7024 29736 7788 29764
rect 5813 29699 5871 29705
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 7024 29696 7052 29736
rect 7285 29699 7343 29705
rect 7285 29696 7297 29699
rect 5859 29668 7052 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 5537 29631 5595 29637
rect 5537 29597 5549 29631
rect 5583 29597 5595 29631
rect 5537 29591 5595 29597
rect 5721 29631 5779 29637
rect 5721 29597 5733 29631
rect 5767 29597 5779 29631
rect 5721 29591 5779 29597
rect 5074 29520 5080 29572
rect 5132 29560 5138 29572
rect 5736 29560 5764 29591
rect 5132 29532 5764 29560
rect 5132 29520 5138 29532
rect 5828 29492 5856 29659
rect 6822 29588 6828 29640
rect 6880 29588 6886 29640
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29628 6975 29631
rect 7024 29628 7052 29668
rect 7116 29668 7297 29696
rect 7116 29637 7144 29668
rect 7285 29665 7297 29668
rect 7331 29665 7343 29699
rect 7285 29659 7343 29665
rect 7392 29668 7604 29696
rect 6963 29600 7052 29628
rect 7101 29631 7159 29637
rect 6963 29597 6975 29600
rect 6917 29591 6975 29597
rect 7101 29597 7113 29631
rect 7147 29597 7159 29631
rect 7101 29591 7159 29597
rect 7190 29588 7196 29640
rect 7248 29588 7254 29640
rect 7006 29520 7012 29572
rect 7064 29560 7070 29572
rect 7392 29560 7420 29668
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 7469 29591 7527 29597
rect 7064 29532 7420 29560
rect 7064 29520 7070 29532
rect 5000 29464 5856 29492
rect 6454 29452 6460 29504
rect 6512 29492 6518 29504
rect 7484 29492 7512 29591
rect 7576 29560 7604 29668
rect 7760 29637 7788 29736
rect 8021 29699 8079 29705
rect 8021 29665 8033 29699
rect 8067 29696 8079 29699
rect 8680 29696 8708 29792
rect 12621 29767 12679 29773
rect 12621 29733 12633 29767
rect 12667 29764 12679 29767
rect 12667 29733 12680 29764
rect 12621 29727 12680 29733
rect 8067 29668 8708 29696
rect 8067 29665 8079 29668
rect 8021 29659 8079 29665
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29628 7803 29631
rect 7834 29628 7840 29640
rect 7791 29600 7840 29628
rect 7791 29597 7803 29600
rect 7745 29591 7803 29597
rect 7834 29588 7840 29600
rect 7892 29588 7898 29640
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29597 7987 29631
rect 7929 29591 7987 29597
rect 7944 29560 7972 29591
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 8404 29637 8432 29668
rect 11238 29656 11244 29708
rect 11296 29696 11302 29708
rect 12161 29699 12219 29705
rect 11296 29668 11836 29696
rect 11296 29656 11302 29668
rect 8389 29631 8447 29637
rect 8389 29597 8401 29631
rect 8435 29597 8447 29631
rect 8389 29591 8447 29597
rect 8665 29631 8723 29637
rect 8665 29597 8677 29631
rect 8711 29597 8723 29631
rect 8665 29591 8723 29597
rect 7576 29532 7972 29560
rect 8680 29560 8708 29591
rect 9306 29588 9312 29640
rect 9364 29588 9370 29640
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29628 9551 29631
rect 9950 29628 9956 29640
rect 9539 29600 9956 29628
rect 9539 29597 9551 29600
rect 9493 29591 9551 29597
rect 9508 29560 9536 29591
rect 9950 29588 9956 29600
rect 10008 29588 10014 29640
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29628 10471 29631
rect 10778 29628 10784 29640
rect 10459 29600 10784 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 8680 29532 9536 29560
rect 10152 29560 10180 29591
rect 10778 29588 10784 29600
rect 10836 29588 10842 29640
rect 11808 29637 11836 29668
rect 12161 29665 12173 29699
rect 12207 29696 12219 29699
rect 12250 29696 12256 29708
rect 12207 29668 12256 29696
rect 12207 29665 12219 29668
rect 12161 29659 12219 29665
rect 12250 29656 12256 29668
rect 12308 29656 12314 29708
rect 12652 29685 12680 29727
rect 12802 29724 12808 29776
rect 12860 29764 12866 29776
rect 14553 29767 14611 29773
rect 14553 29764 14565 29767
rect 12860 29736 14565 29764
rect 12860 29724 12866 29736
rect 14553 29733 14565 29736
rect 14599 29733 14611 29767
rect 14553 29727 14611 29733
rect 14660 29736 15424 29764
rect 14660 29708 14688 29736
rect 12710 29685 12716 29708
rect 12652 29657 12716 29685
rect 12710 29656 12716 29657
rect 12768 29656 12774 29708
rect 13354 29656 13360 29708
rect 13412 29656 13418 29708
rect 14458 29696 14464 29708
rect 13556 29668 14464 29696
rect 11609 29631 11667 29637
rect 11609 29597 11621 29631
rect 11655 29597 11667 29631
rect 11609 29591 11667 29597
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29597 11851 29631
rect 11793 29591 11851 29597
rect 11146 29560 11152 29572
rect 10152 29532 11152 29560
rect 11146 29520 11152 29532
rect 11204 29520 11210 29572
rect 10226 29492 10232 29504
rect 6512 29464 10232 29492
rect 6512 29452 6518 29464
rect 10226 29452 10232 29464
rect 10284 29452 10290 29504
rect 10318 29452 10324 29504
rect 10376 29452 10382 29504
rect 11625 29492 11653 29591
rect 11882 29588 11888 29640
rect 11940 29588 11946 29640
rect 11974 29588 11980 29640
rect 12032 29588 12038 29640
rect 12986 29588 12992 29640
rect 13044 29628 13050 29640
rect 13081 29631 13139 29637
rect 13081 29628 13093 29631
rect 13044 29600 13093 29628
rect 13044 29588 13050 29600
rect 13081 29597 13093 29600
rect 13127 29597 13139 29631
rect 13081 29591 13139 29597
rect 13170 29588 13176 29640
rect 13228 29628 13234 29640
rect 13556 29637 13584 29668
rect 14458 29656 14464 29668
rect 14516 29656 14522 29708
rect 14642 29656 14648 29708
rect 14700 29656 14706 29708
rect 14737 29699 14795 29705
rect 14737 29665 14749 29699
rect 14783 29696 14795 29699
rect 14826 29696 14832 29708
rect 14783 29668 14832 29696
rect 14783 29665 14795 29668
rect 14737 29659 14795 29665
rect 14826 29656 14832 29668
rect 14884 29656 14890 29708
rect 13541 29631 13599 29637
rect 13541 29628 13553 29631
rect 13228 29600 13553 29628
rect 13228 29588 13234 29600
rect 13541 29597 13553 29600
rect 13587 29597 13599 29631
rect 13541 29591 13599 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29597 13783 29631
rect 13725 29591 13783 29597
rect 12158 29520 12164 29572
rect 12216 29520 12222 29572
rect 12342 29569 12348 29572
rect 12299 29563 12348 29569
rect 12299 29529 12311 29563
rect 12345 29529 12348 29563
rect 12299 29523 12348 29529
rect 12342 29520 12348 29523
rect 12400 29520 12406 29572
rect 12469 29563 12527 29569
rect 12469 29560 12481 29563
rect 12452 29529 12481 29560
rect 12515 29560 12527 29563
rect 13633 29563 13691 29569
rect 13633 29560 13645 29563
rect 12515 29532 13645 29560
rect 12515 29529 12527 29532
rect 12452 29523 12527 29529
rect 13633 29529 13645 29532
rect 13679 29529 13691 29563
rect 13633 29523 13691 29529
rect 13740 29560 13768 29591
rect 14274 29588 14280 29640
rect 14332 29588 14338 29640
rect 14369 29631 14427 29637
rect 14369 29597 14381 29631
rect 14415 29628 14427 29631
rect 14918 29628 14924 29640
rect 14415 29600 14924 29628
rect 14415 29597 14427 29600
rect 14369 29591 14427 29597
rect 14918 29588 14924 29600
rect 14976 29628 14982 29640
rect 15396 29637 15424 29736
rect 15470 29724 15476 29776
rect 15528 29764 15534 29776
rect 16025 29767 16083 29773
rect 16025 29764 16037 29767
rect 15528 29736 16037 29764
rect 15528 29724 15534 29736
rect 16025 29733 16037 29736
rect 16071 29733 16083 29767
rect 17236 29764 17264 29792
rect 22462 29764 22468 29776
rect 16025 29727 16083 29733
rect 16592 29736 17264 29764
rect 20548 29736 22468 29764
rect 16592 29705 16620 29736
rect 20548 29708 20576 29736
rect 16577 29699 16635 29705
rect 15764 29668 16068 29696
rect 15562 29637 15568 29640
rect 15381 29631 15439 29637
rect 14976 29600 15238 29628
rect 14976 29588 14982 29600
rect 15105 29563 15163 29569
rect 15105 29560 15117 29563
rect 13740 29532 15117 29560
rect 12452 29492 12480 29523
rect 11625 29464 12480 29492
rect 12710 29452 12716 29504
rect 12768 29452 12774 29504
rect 13538 29452 13544 29504
rect 13596 29492 13602 29504
rect 13740 29492 13768 29532
rect 15105 29529 15117 29532
rect 15151 29529 15163 29563
rect 15210 29560 15238 29600
rect 15381 29597 15393 29631
rect 15427 29597 15439 29631
rect 15381 29591 15439 29597
rect 15529 29631 15568 29637
rect 15529 29597 15541 29631
rect 15620 29628 15626 29640
rect 15764 29628 15792 29668
rect 15620 29600 15792 29628
rect 15529 29591 15568 29597
rect 15562 29588 15568 29591
rect 15620 29588 15626 29600
rect 15838 29588 15844 29640
rect 15896 29637 15902 29640
rect 15896 29628 15904 29637
rect 16040 29628 16068 29668
rect 16577 29665 16589 29699
rect 16623 29665 16635 29699
rect 16577 29659 16635 29665
rect 16758 29656 16764 29708
rect 16816 29696 16822 29708
rect 17681 29699 17739 29705
rect 17681 29696 17693 29699
rect 16816 29668 17693 29696
rect 16816 29656 16822 29668
rect 17681 29665 17693 29668
rect 17727 29665 17739 29699
rect 17681 29659 17739 29665
rect 20530 29656 20536 29708
rect 20588 29656 20594 29708
rect 20717 29699 20775 29705
rect 20717 29665 20729 29699
rect 20763 29696 20775 29699
rect 21453 29699 21511 29705
rect 21453 29696 21465 29699
rect 20763 29668 21465 29696
rect 20763 29665 20775 29668
rect 20717 29659 20775 29665
rect 21453 29665 21465 29668
rect 21499 29665 21511 29699
rect 21453 29659 21511 29665
rect 15896 29600 15941 29628
rect 16040 29600 17264 29628
rect 15896 29591 15904 29600
rect 15896 29588 15902 29591
rect 15657 29563 15715 29569
rect 15657 29560 15669 29563
rect 15210 29532 15669 29560
rect 15105 29523 15163 29529
rect 15657 29529 15669 29532
rect 15703 29529 15715 29563
rect 15657 29523 15715 29529
rect 15749 29563 15807 29569
rect 15749 29529 15761 29563
rect 15795 29560 15807 29563
rect 16114 29560 16120 29572
rect 15795 29532 16120 29560
rect 15795 29529 15807 29532
rect 15749 29523 15807 29529
rect 16114 29520 16120 29532
rect 16172 29520 16178 29572
rect 13596 29464 13768 29492
rect 13596 29452 13602 29464
rect 16482 29452 16488 29504
rect 16540 29492 16546 29504
rect 17129 29495 17187 29501
rect 17129 29492 17141 29495
rect 16540 29464 17141 29492
rect 16540 29452 16546 29464
rect 17129 29461 17141 29464
rect 17175 29461 17187 29495
rect 17236 29492 17264 29600
rect 17586 29588 17592 29640
rect 17644 29628 17650 29640
rect 19245 29631 19303 29637
rect 17644 29600 18644 29628
rect 17644 29588 17650 29600
rect 17497 29563 17555 29569
rect 17497 29529 17509 29563
rect 17543 29560 17555 29563
rect 17770 29560 17776 29572
rect 17543 29532 17776 29560
rect 17543 29529 17555 29532
rect 17497 29523 17555 29529
rect 17770 29520 17776 29532
rect 17828 29520 17834 29572
rect 17948 29563 18006 29569
rect 17948 29529 17960 29563
rect 17994 29560 18006 29563
rect 18506 29560 18512 29572
rect 17994 29532 18512 29560
rect 17994 29529 18006 29532
rect 17948 29523 18006 29529
rect 18506 29520 18512 29532
rect 18564 29520 18570 29572
rect 18616 29560 18644 29600
rect 19245 29597 19257 29631
rect 19291 29628 19303 29631
rect 19794 29628 19800 29640
rect 19291 29600 19800 29628
rect 19291 29597 19303 29600
rect 19245 29591 19303 29597
rect 19794 29588 19800 29600
rect 19852 29628 19858 29640
rect 19852 29600 20944 29628
rect 19852 29588 19858 29600
rect 19512 29563 19570 29569
rect 18616 29532 19472 29560
rect 18322 29492 18328 29504
rect 17236 29464 18328 29492
rect 17129 29455 17187 29461
rect 18322 29452 18328 29464
rect 18380 29492 18386 29504
rect 19061 29495 19119 29501
rect 19061 29492 19073 29495
rect 18380 29464 19073 29492
rect 18380 29452 18386 29464
rect 19061 29461 19073 29464
rect 19107 29461 19119 29495
rect 19444 29492 19472 29532
rect 19512 29529 19524 29563
rect 19558 29560 19570 29563
rect 20806 29560 20812 29572
rect 19558 29532 20812 29560
rect 19558 29529 19570 29532
rect 19512 29523 19570 29529
rect 20806 29520 20812 29532
rect 20864 29520 20870 29572
rect 20916 29560 20944 29600
rect 20990 29588 20996 29640
rect 21048 29588 21054 29640
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29597 21143 29631
rect 21085 29591 21143 29597
rect 21100 29560 21128 29591
rect 21174 29588 21180 29640
rect 21232 29588 21238 29640
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29628 21419 29631
rect 21560 29628 21588 29736
rect 22462 29724 22468 29736
rect 22520 29724 22526 29776
rect 24946 29764 24952 29776
rect 22940 29736 24952 29764
rect 22278 29656 22284 29708
rect 22336 29696 22342 29708
rect 22940 29696 22968 29736
rect 24946 29724 24952 29736
rect 25004 29764 25010 29776
rect 25041 29767 25099 29773
rect 25041 29764 25053 29767
rect 25004 29736 25053 29764
rect 25004 29724 25010 29736
rect 25041 29733 25053 29736
rect 25087 29733 25099 29767
rect 25240 29764 25268 29792
rect 25501 29767 25559 29773
rect 25501 29764 25513 29767
rect 25240 29736 25513 29764
rect 25041 29727 25099 29733
rect 25501 29733 25513 29736
rect 25547 29733 25559 29767
rect 25501 29727 25559 29733
rect 26694 29724 26700 29776
rect 26752 29764 26758 29776
rect 27249 29767 27307 29773
rect 27249 29764 27261 29767
rect 26752 29736 27261 29764
rect 26752 29724 26758 29736
rect 27249 29733 27261 29736
rect 27295 29733 27307 29767
rect 29104 29764 29132 29792
rect 30576 29764 30604 29792
rect 31726 29764 31754 29804
rect 31846 29792 31852 29844
rect 31904 29832 31910 29844
rect 32769 29835 32827 29841
rect 32769 29832 32781 29835
rect 31904 29804 32781 29832
rect 31904 29792 31910 29804
rect 32769 29801 32781 29804
rect 32815 29801 32827 29835
rect 32769 29795 32827 29801
rect 32214 29764 32220 29776
rect 27249 29727 27307 29733
rect 27586 29736 28028 29764
rect 29104 29736 29776 29764
rect 30576 29736 31616 29764
rect 31726 29736 32220 29764
rect 22336 29668 22416 29696
rect 22336 29656 22342 29668
rect 21407 29600 21588 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 22186 29588 22192 29640
rect 22244 29588 22250 29640
rect 22388 29637 22416 29668
rect 22848 29668 22968 29696
rect 22373 29631 22431 29637
rect 22373 29597 22385 29631
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 22738 29588 22744 29640
rect 22796 29588 22802 29640
rect 22848 29560 22876 29668
rect 23106 29656 23112 29708
rect 23164 29656 23170 29708
rect 23566 29696 23572 29708
rect 23216 29668 23572 29696
rect 22922 29588 22928 29640
rect 22980 29588 22986 29640
rect 23216 29637 23244 29668
rect 23566 29656 23572 29668
rect 23624 29696 23630 29708
rect 23624 29668 26944 29696
rect 23624 29656 23630 29668
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29597 23075 29631
rect 23017 29591 23075 29597
rect 23201 29631 23259 29637
rect 23201 29597 23213 29631
rect 23247 29597 23259 29631
rect 23385 29631 23443 29637
rect 23385 29628 23397 29631
rect 23201 29591 23259 29597
rect 23308 29600 23397 29628
rect 20916 29532 21036 29560
rect 21100 29532 22876 29560
rect 20898 29492 20904 29504
rect 19444 29464 20904 29492
rect 19061 29455 19119 29461
rect 20898 29452 20904 29464
rect 20956 29452 20962 29504
rect 21008 29492 21036 29532
rect 22462 29492 22468 29504
rect 21008 29464 22468 29492
rect 22462 29452 22468 29464
rect 22520 29452 22526 29504
rect 22554 29452 22560 29504
rect 22612 29492 22618 29504
rect 23032 29492 23060 29591
rect 22612 29464 23060 29492
rect 22612 29452 22618 29464
rect 23106 29452 23112 29504
rect 23164 29492 23170 29504
rect 23308 29492 23336 29600
rect 23385 29597 23397 29600
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 23753 29631 23811 29637
rect 23753 29628 23765 29631
rect 23532 29600 23765 29628
rect 23532 29588 23538 29600
rect 23753 29597 23765 29600
rect 23799 29597 23811 29631
rect 23753 29591 23811 29597
rect 24578 29588 24584 29640
rect 24636 29588 24642 29640
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 24857 29631 24915 29637
rect 24857 29628 24869 29631
rect 24820 29600 24869 29628
rect 24820 29588 24826 29600
rect 24857 29597 24869 29600
rect 24903 29597 24915 29631
rect 24857 29591 24915 29597
rect 25041 29631 25099 29637
rect 25041 29597 25053 29631
rect 25087 29597 25099 29631
rect 25041 29591 25099 29597
rect 23566 29520 23572 29572
rect 23624 29520 23630 29572
rect 23658 29520 23664 29572
rect 23716 29520 23722 29572
rect 25056 29560 25084 29591
rect 25222 29588 25228 29640
rect 25280 29588 25286 29640
rect 26237 29631 26295 29637
rect 26237 29597 26249 29631
rect 26283 29628 26295 29631
rect 26916 29628 26944 29668
rect 27430 29656 27436 29708
rect 27488 29696 27494 29708
rect 27586 29696 27614 29736
rect 27488 29668 27614 29696
rect 27488 29656 27494 29668
rect 26283 29600 26556 29628
rect 26916 29600 27197 29628
rect 26283 29597 26295 29600
rect 26237 29591 26295 29597
rect 26528 29572 26556 29600
rect 25130 29560 25136 29572
rect 25056 29532 25136 29560
rect 25130 29520 25136 29532
rect 25188 29520 25194 29572
rect 26326 29520 26332 29572
rect 26384 29560 26390 29572
rect 26421 29563 26479 29569
rect 26421 29560 26433 29563
rect 26384 29532 26433 29560
rect 26384 29520 26390 29532
rect 26421 29529 26433 29532
rect 26467 29529 26479 29563
rect 26421 29523 26479 29529
rect 26510 29520 26516 29572
rect 26568 29520 26574 29572
rect 26878 29520 26884 29572
rect 26936 29520 26942 29572
rect 27065 29563 27123 29569
rect 27065 29529 27077 29563
rect 27111 29529 27123 29563
rect 27065 29523 27123 29529
rect 23164 29464 23336 29492
rect 23937 29495 23995 29501
rect 23164 29452 23170 29464
rect 23937 29461 23949 29495
rect 23983 29492 23995 29495
rect 24118 29492 24124 29504
rect 23983 29464 24124 29492
rect 23983 29461 23995 29464
rect 23937 29455 23995 29461
rect 24118 29452 24124 29464
rect 24176 29452 24182 29504
rect 24854 29452 24860 29504
rect 24912 29492 24918 29504
rect 25682 29492 25688 29504
rect 24912 29464 25688 29492
rect 24912 29452 24918 29464
rect 25682 29452 25688 29464
rect 25740 29452 25746 29504
rect 26050 29452 26056 29504
rect 26108 29492 26114 29504
rect 27080 29492 27108 29523
rect 26108 29464 27108 29492
rect 27169 29492 27197 29600
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 28000 29637 28028 29736
rect 28460 29668 29408 29696
rect 28460 29640 28488 29668
rect 27341 29631 27399 29637
rect 27341 29628 27353 29631
rect 27304 29600 27353 29628
rect 27304 29588 27310 29600
rect 27341 29597 27353 29600
rect 27387 29628 27399 29631
rect 27801 29631 27859 29637
rect 27801 29628 27813 29631
rect 27387 29600 27813 29628
rect 27387 29597 27399 29600
rect 27341 29591 27399 29597
rect 27801 29597 27813 29600
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 27985 29631 28043 29637
rect 27985 29597 27997 29631
rect 28031 29597 28043 29631
rect 27985 29591 28043 29597
rect 27430 29520 27436 29572
rect 27488 29560 27494 29572
rect 27525 29563 27583 29569
rect 27525 29560 27537 29563
rect 27488 29532 27537 29560
rect 27488 29520 27494 29532
rect 27525 29529 27537 29532
rect 27571 29529 27583 29563
rect 27816 29560 27844 29591
rect 28442 29588 28448 29640
rect 28500 29588 28506 29640
rect 28626 29588 28632 29640
rect 28684 29628 28690 29640
rect 29380 29637 29408 29668
rect 29181 29631 29239 29637
rect 29181 29628 29193 29631
rect 28684 29600 29193 29628
rect 28684 29588 28690 29600
rect 29181 29597 29193 29600
rect 29227 29597 29239 29631
rect 29181 29591 29239 29597
rect 29365 29631 29423 29637
rect 29365 29597 29377 29631
rect 29411 29628 29423 29631
rect 29546 29628 29552 29640
rect 29411 29600 29552 29628
rect 29411 29597 29423 29600
rect 29365 29591 29423 29597
rect 29546 29588 29552 29600
rect 29604 29588 29610 29640
rect 29748 29628 29776 29736
rect 30561 29699 30619 29705
rect 30561 29665 30573 29699
rect 30607 29696 30619 29699
rect 30650 29696 30656 29708
rect 30607 29668 30656 29696
rect 30607 29665 30619 29668
rect 30561 29659 30619 29665
rect 30650 29656 30656 29668
rect 30708 29656 30714 29708
rect 31588 29696 31616 29736
rect 32214 29724 32220 29736
rect 32272 29724 32278 29776
rect 31757 29699 31815 29705
rect 31757 29696 31769 29699
rect 30760 29668 31524 29696
rect 31588 29668 31769 29696
rect 30282 29628 30288 29640
rect 29748 29600 30288 29628
rect 30282 29588 30288 29600
rect 30340 29588 30346 29640
rect 30466 29588 30472 29640
rect 30524 29588 30530 29640
rect 30760 29637 30788 29668
rect 30745 29631 30803 29637
rect 30745 29597 30757 29631
rect 30791 29597 30803 29631
rect 30745 29591 30803 29597
rect 31021 29631 31079 29637
rect 31021 29597 31033 29631
rect 31067 29628 31079 29631
rect 31110 29628 31116 29640
rect 31067 29600 31116 29628
rect 31067 29597 31079 29600
rect 31021 29591 31079 29597
rect 31110 29588 31116 29600
rect 31168 29588 31174 29640
rect 31386 29588 31392 29640
rect 31444 29588 31450 29640
rect 31496 29630 31524 29668
rect 31757 29665 31769 29668
rect 31803 29665 31815 29699
rect 31757 29659 31815 29665
rect 32401 29631 32459 29637
rect 31496 29628 31616 29630
rect 32401 29628 32413 29631
rect 31496 29602 32413 29628
rect 31588 29600 32413 29602
rect 32401 29597 32413 29600
rect 32447 29597 32459 29631
rect 32784 29628 32812 29795
rect 32953 29631 33011 29637
rect 32953 29628 32965 29631
rect 32784 29600 32965 29628
rect 32401 29591 32459 29597
rect 32953 29597 32965 29600
rect 32999 29628 33011 29631
rect 35253 29631 35311 29637
rect 35253 29628 35265 29631
rect 32999 29600 35265 29628
rect 32999 29597 33011 29600
rect 32953 29591 33011 29597
rect 35253 29597 35265 29600
rect 35299 29628 35311 29631
rect 35437 29631 35495 29637
rect 35437 29628 35449 29631
rect 35299 29600 35449 29628
rect 35299 29597 35311 29600
rect 35253 29591 35311 29597
rect 35437 29597 35449 29600
rect 35483 29597 35495 29631
rect 35437 29591 35495 29597
rect 29086 29560 29092 29572
rect 27816 29532 29092 29560
rect 27525 29523 27583 29529
rect 29086 29520 29092 29532
rect 29144 29520 29150 29572
rect 30006 29560 30012 29572
rect 29196 29532 30012 29560
rect 29196 29492 29224 29532
rect 30006 29520 30012 29532
rect 30064 29520 30070 29572
rect 30558 29520 30564 29572
rect 30616 29560 30622 29572
rect 30834 29560 30840 29572
rect 30616 29532 30840 29560
rect 30616 29520 30622 29532
rect 30834 29520 30840 29532
rect 30892 29560 30898 29572
rect 31205 29563 31263 29569
rect 31205 29560 31217 29563
rect 30892 29532 31217 29560
rect 30892 29520 30898 29532
rect 31205 29529 31217 29532
rect 31251 29529 31263 29563
rect 31205 29523 31263 29529
rect 31294 29520 31300 29572
rect 31352 29520 31358 29572
rect 32030 29520 32036 29572
rect 32088 29560 32094 29572
rect 33689 29563 33747 29569
rect 33689 29560 33701 29563
rect 32088 29532 33701 29560
rect 32088 29520 32094 29532
rect 33689 29529 33701 29532
rect 33735 29529 33747 29563
rect 33689 29523 33747 29529
rect 36262 29520 36268 29572
rect 36320 29520 36326 29572
rect 27169 29464 29224 29492
rect 29273 29495 29331 29501
rect 26108 29452 26114 29464
rect 29273 29461 29285 29495
rect 29319 29492 29331 29495
rect 30282 29492 30288 29504
rect 29319 29464 30288 29492
rect 29319 29461 29331 29464
rect 29273 29455 29331 29461
rect 30282 29452 30288 29464
rect 30340 29452 30346 29504
rect 30377 29495 30435 29501
rect 30377 29461 30389 29495
rect 30423 29492 30435 29495
rect 31478 29492 31484 29504
rect 30423 29464 31484 29492
rect 30423 29461 30435 29464
rect 30377 29455 30435 29461
rect 31478 29452 31484 29464
rect 31536 29452 31542 29504
rect 31570 29452 31576 29504
rect 31628 29452 31634 29504
rect 1104 29402 43884 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 43884 29402
rect 1104 29328 43884 29350
rect 2682 29288 2688 29300
rect 2148 29260 2688 29288
rect 1854 29180 1860 29232
rect 1912 29180 1918 29232
rect 2148 29161 2176 29260
rect 2682 29248 2688 29260
rect 2740 29288 2746 29300
rect 3437 29291 3495 29297
rect 3437 29288 3449 29291
rect 2740 29260 3449 29288
rect 2740 29248 2746 29260
rect 3437 29257 3449 29260
rect 3483 29257 3495 29291
rect 3437 29251 3495 29257
rect 3602 29248 3608 29300
rect 3660 29248 3666 29300
rect 3789 29291 3847 29297
rect 3789 29257 3801 29291
rect 3835 29288 3847 29291
rect 4062 29288 4068 29300
rect 3835 29260 4068 29288
rect 3835 29257 3847 29260
rect 3789 29251 3847 29257
rect 4062 29248 4068 29260
rect 4120 29248 4126 29300
rect 4614 29248 4620 29300
rect 4672 29248 4678 29300
rect 4807 29291 4865 29297
rect 4807 29257 4819 29291
rect 4853 29288 4865 29291
rect 5074 29288 5080 29300
rect 4853 29260 5080 29288
rect 4853 29257 4865 29260
rect 4807 29251 4865 29257
rect 5074 29248 5080 29260
rect 5132 29248 5138 29300
rect 5169 29291 5227 29297
rect 5169 29257 5181 29291
rect 5215 29288 5227 29291
rect 5258 29288 5264 29300
rect 5215 29260 5264 29288
rect 5215 29257 5227 29260
rect 5169 29251 5227 29257
rect 5258 29248 5264 29260
rect 5316 29248 5322 29300
rect 7006 29288 7012 29300
rect 6748 29260 7012 29288
rect 2593 29223 2651 29229
rect 2593 29189 2605 29223
rect 2639 29220 2651 29223
rect 3237 29223 3295 29229
rect 2639 29192 2912 29220
rect 2639 29189 2651 29192
rect 2593 29183 2651 29189
rect 2884 29161 2912 29192
rect 3237 29189 3249 29223
rect 3283 29220 3295 29223
rect 3326 29220 3332 29232
rect 3283 29192 3332 29220
rect 3283 29189 3295 29192
rect 3237 29183 3295 29189
rect 3326 29180 3332 29192
rect 3384 29180 3390 29232
rect 3620 29220 3648 29248
rect 4632 29220 4660 29248
rect 4893 29223 4951 29229
rect 4893 29220 4905 29223
rect 3620 29192 3924 29220
rect 4632 29192 4905 29220
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29121 2099 29155
rect 2041 29115 2099 29121
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29121 2191 29155
rect 2133 29115 2191 29121
rect 2409 29155 2467 29161
rect 2409 29121 2421 29155
rect 2455 29152 2467 29155
rect 2685 29155 2743 29161
rect 2455 29124 2636 29152
rect 2455 29121 2467 29124
rect 2409 29115 2467 29121
rect 2056 29084 2084 29115
rect 2608 29096 2636 29124
rect 2685 29121 2697 29155
rect 2731 29121 2743 29155
rect 2685 29115 2743 29121
rect 2869 29155 2927 29161
rect 2869 29121 2881 29155
rect 2915 29121 2927 29155
rect 2869 29115 2927 29121
rect 2498 29084 2504 29096
rect 2056 29056 2504 29084
rect 2498 29044 2504 29056
rect 2556 29044 2562 29096
rect 2590 29044 2596 29096
rect 2648 29044 2654 29096
rect 1486 28976 1492 29028
rect 1544 29016 1550 29028
rect 1673 29019 1731 29025
rect 1673 29016 1685 29019
rect 1544 28988 1685 29016
rect 1544 28976 1550 28988
rect 1673 28985 1685 28988
rect 1719 28985 1731 29019
rect 1673 28979 1731 28985
rect 1857 29019 1915 29025
rect 1857 28985 1869 29019
rect 1903 29016 1915 29019
rect 2314 29016 2320 29028
rect 1903 28988 2320 29016
rect 1903 28985 1915 28988
rect 1857 28979 1915 28985
rect 2314 28976 2320 28988
rect 2372 28976 2378 29028
rect 2700 29016 2728 29115
rect 2884 29084 2912 29115
rect 3050 29112 3056 29164
rect 3108 29112 3114 29164
rect 3896 29161 3924 29192
rect 4893 29189 4905 29192
rect 4939 29220 4951 29223
rect 6638 29220 6644 29232
rect 4939 29192 6644 29220
rect 4939 29189 4951 29192
rect 4893 29183 4951 29189
rect 6638 29180 6644 29192
rect 6696 29180 6702 29232
rect 3697 29155 3755 29161
rect 3697 29121 3709 29155
rect 3743 29121 3755 29155
rect 3697 29115 3755 29121
rect 3881 29155 3939 29161
rect 3881 29121 3893 29155
rect 3927 29121 3939 29155
rect 3881 29115 3939 29121
rect 3234 29084 3240 29096
rect 2884 29056 3240 29084
rect 3234 29044 3240 29056
rect 3292 29044 3298 29096
rect 3418 29044 3424 29096
rect 3476 29084 3482 29096
rect 3712 29084 3740 29115
rect 4522 29112 4528 29164
rect 4580 29112 4586 29164
rect 4706 29112 4712 29164
rect 4764 29112 4770 29164
rect 4982 29112 4988 29164
rect 5040 29112 5046 29164
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 5273 29158 5331 29161
rect 5273 29155 5393 29158
rect 5273 29121 5285 29155
rect 5319 29152 5393 29155
rect 5442 29152 5448 29164
rect 5319 29130 5448 29152
rect 5319 29121 5331 29130
rect 5365 29124 5448 29130
rect 5273 29115 5331 29121
rect 3476 29056 3740 29084
rect 3476 29044 3482 29056
rect 2608 28988 2728 29016
rect 2869 29019 2927 29025
rect 1762 28908 1768 28960
rect 1820 28948 1826 28960
rect 2222 28948 2228 28960
rect 1820 28920 2228 28948
rect 1820 28908 1826 28920
rect 2222 28908 2228 28920
rect 2280 28908 2286 28960
rect 2406 28908 2412 28960
rect 2464 28948 2470 28960
rect 2608 28948 2636 28988
rect 2869 28985 2881 29019
rect 2915 29016 2927 29019
rect 3142 29016 3148 29028
rect 2915 28988 3148 29016
rect 2915 28985 2927 28988
rect 2869 28979 2927 28985
rect 3142 28976 3148 28988
rect 3200 29016 3206 29028
rect 5092 29016 5120 29115
rect 5442 29112 5448 29124
rect 5500 29112 5506 29164
rect 6748 29084 6776 29260
rect 7006 29248 7012 29260
rect 7064 29248 7070 29300
rect 7834 29288 7840 29300
rect 7116 29260 7840 29288
rect 6825 29155 6883 29161
rect 6825 29121 6837 29155
rect 6871 29152 6883 29155
rect 6871 29124 6960 29152
rect 6871 29121 6883 29124
rect 6825 29115 6883 29121
rect 6932 29084 6960 29124
rect 7006 29112 7012 29164
rect 7064 29112 7070 29164
rect 7116 29161 7144 29260
rect 7834 29248 7840 29260
rect 7892 29288 7898 29300
rect 7945 29291 8003 29297
rect 7945 29288 7957 29291
rect 7892 29260 7957 29288
rect 7892 29248 7898 29260
rect 7945 29257 7957 29260
rect 7991 29257 8003 29291
rect 7945 29251 8003 29257
rect 8110 29248 8116 29300
rect 8168 29248 8174 29300
rect 9039 29291 9097 29297
rect 9039 29257 9051 29291
rect 9085 29288 9097 29291
rect 9306 29288 9312 29300
rect 9085 29260 9312 29288
rect 9085 29257 9097 29260
rect 9039 29251 9097 29257
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 9490 29248 9496 29300
rect 9548 29288 9554 29300
rect 9548 29260 10088 29288
rect 9548 29248 9554 29260
rect 7745 29223 7803 29229
rect 7745 29220 7757 29223
rect 7208 29192 7757 29220
rect 7101 29155 7159 29161
rect 7101 29121 7113 29155
rect 7147 29121 7159 29155
rect 7101 29115 7159 29121
rect 7208 29084 7236 29192
rect 7282 29112 7288 29164
rect 7340 29152 7346 29164
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 7340 29124 7389 29152
rect 7340 29112 7346 29124
rect 7377 29121 7389 29124
rect 7423 29121 7435 29155
rect 7377 29115 7435 29121
rect 6748 29056 6868 29084
rect 6932 29056 7236 29084
rect 6840 29025 6868 29056
rect 6825 29019 6883 29025
rect 3200 28988 5856 29016
rect 3200 28976 3206 28988
rect 5828 28960 5856 28988
rect 6825 28985 6837 29019
rect 6871 28985 6883 29019
rect 7392 29016 7420 29115
rect 7558 29112 7564 29164
rect 7616 29112 7622 29164
rect 7668 29161 7696 29192
rect 7745 29189 7757 29192
rect 7791 29220 7803 29223
rect 8386 29220 8392 29232
rect 7791 29192 8392 29220
rect 7791 29189 7803 29192
rect 7745 29183 7803 29189
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 10060 29229 10088 29260
rect 10318 29248 10324 29300
rect 10376 29288 10382 29300
rect 10689 29291 10747 29297
rect 10689 29288 10701 29291
rect 10376 29260 10701 29288
rect 10376 29248 10382 29260
rect 10689 29257 10701 29260
rect 10735 29257 10747 29291
rect 10689 29251 10747 29257
rect 11238 29248 11244 29300
rect 11296 29288 11302 29300
rect 11606 29288 11612 29300
rect 11296 29260 11612 29288
rect 11296 29248 11302 29260
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 12526 29288 12532 29300
rect 12216 29260 12532 29288
rect 12216 29248 12222 29260
rect 12526 29248 12532 29260
rect 12584 29248 12590 29300
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 12805 29291 12863 29297
rect 12805 29257 12817 29291
rect 12851 29288 12863 29291
rect 12851 29260 12940 29288
rect 12851 29257 12863 29260
rect 12805 29251 12863 29257
rect 12912 29232 12940 29260
rect 13078 29248 13084 29300
rect 13136 29288 13142 29300
rect 14737 29291 14795 29297
rect 14737 29288 14749 29291
rect 13136 29260 14749 29288
rect 13136 29248 13142 29260
rect 14737 29257 14749 29260
rect 14783 29257 14795 29291
rect 14737 29251 14795 29257
rect 16942 29248 16948 29300
rect 17000 29288 17006 29300
rect 17865 29291 17923 29297
rect 17865 29288 17877 29291
rect 17000 29260 17877 29288
rect 17000 29248 17006 29260
rect 17865 29257 17877 29260
rect 17911 29257 17923 29291
rect 17865 29251 17923 29257
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18325 29291 18383 29297
rect 18325 29288 18337 29291
rect 18196 29260 18337 29288
rect 18196 29248 18202 29260
rect 18325 29257 18337 29260
rect 18371 29257 18383 29291
rect 18325 29251 18383 29257
rect 18506 29248 18512 29300
rect 18564 29248 18570 29300
rect 18874 29248 18880 29300
rect 18932 29248 18938 29300
rect 19242 29248 19248 29300
rect 19300 29248 19306 29300
rect 19429 29291 19487 29297
rect 19429 29257 19441 29291
rect 19475 29288 19487 29291
rect 19610 29288 19616 29300
rect 19475 29260 19616 29288
rect 19475 29257 19487 29260
rect 19429 29251 19487 29257
rect 19610 29248 19616 29260
rect 19668 29248 19674 29300
rect 20714 29288 20720 29300
rect 19812 29260 20720 29288
rect 8941 29223 8999 29229
rect 8941 29189 8953 29223
rect 8987 29189 8999 29223
rect 8941 29183 8999 29189
rect 9677 29223 9735 29229
rect 9677 29189 9689 29223
rect 9723 29189 9735 29223
rect 9677 29183 9735 29189
rect 10045 29223 10103 29229
rect 10045 29189 10057 29223
rect 10091 29189 10103 29223
rect 10045 29183 10103 29189
rect 7653 29155 7711 29161
rect 7653 29121 7665 29155
rect 7699 29121 7711 29155
rect 7653 29115 7711 29121
rect 8956 29096 8984 29183
rect 9125 29155 9183 29161
rect 9125 29121 9137 29155
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 8938 29044 8944 29096
rect 8996 29044 9002 29096
rect 9140 29084 9168 29115
rect 9214 29112 9220 29164
rect 9272 29112 9278 29164
rect 9490 29112 9496 29164
rect 9548 29161 9554 29164
rect 9548 29155 9570 29161
rect 9558 29121 9570 29155
rect 9692 29152 9720 29183
rect 10410 29180 10416 29232
rect 10468 29180 10474 29232
rect 10502 29180 10508 29232
rect 10560 29183 10566 29232
rect 10796 29192 11008 29220
rect 10560 29180 10573 29183
rect 10515 29177 10573 29180
rect 9548 29115 9570 29121
rect 9646 29124 9720 29152
rect 9548 29112 9554 29115
rect 9306 29084 9312 29096
rect 9140 29056 9312 29084
rect 9306 29044 9312 29056
rect 9364 29044 9370 29096
rect 9646 29095 9674 29124
rect 9766 29112 9772 29164
rect 9824 29112 9830 29164
rect 10229 29155 10287 29161
rect 10229 29121 10241 29155
rect 10275 29121 10287 29155
rect 10515 29143 10527 29177
rect 10561 29143 10573 29177
rect 10515 29137 10573 29143
rect 10229 29115 10287 29121
rect 9600 29067 9674 29095
rect 10244 29084 10272 29115
rect 10796 29084 10824 29192
rect 10870 29112 10876 29164
rect 10928 29112 10934 29164
rect 9122 29016 9128 29028
rect 7392 28988 9128 29016
rect 6825 28979 6883 28985
rect 9122 28976 9128 28988
rect 9180 28976 9186 29028
rect 2464 28920 2636 28948
rect 2464 28908 2470 28920
rect 2774 28908 2780 28960
rect 2832 28948 2838 28960
rect 3326 28948 3332 28960
rect 2832 28920 3332 28948
rect 2832 28908 2838 28920
rect 3326 28908 3332 28920
rect 3384 28908 3390 28960
rect 3418 28908 3424 28960
rect 3476 28908 3482 28960
rect 4249 28951 4307 28957
rect 4249 28917 4261 28951
rect 4295 28948 4307 28951
rect 4798 28948 4804 28960
rect 4295 28920 4804 28948
rect 4295 28917 4307 28920
rect 4249 28911 4307 28917
rect 4798 28908 4804 28920
rect 4856 28908 4862 28960
rect 5810 28908 5816 28960
rect 5868 28908 5874 28960
rect 7006 28908 7012 28960
rect 7064 28948 7070 28960
rect 7193 28951 7251 28957
rect 7193 28948 7205 28951
rect 7064 28920 7205 28948
rect 7064 28908 7070 28920
rect 7193 28917 7205 28920
rect 7239 28948 7251 28951
rect 7929 28951 7987 28957
rect 7929 28948 7941 28951
rect 7239 28920 7941 28948
rect 7239 28917 7251 28920
rect 7193 28911 7251 28917
rect 7929 28917 7941 28920
rect 7975 28917 7987 28951
rect 7929 28911 7987 28917
rect 8294 28908 8300 28960
rect 8352 28948 8358 28960
rect 9600 28948 9628 29067
rect 10244 29056 10824 29084
rect 10888 29016 10916 29112
rect 10980 29084 11008 29192
rect 11330 29180 11336 29232
rect 11388 29220 11394 29232
rect 11388 29192 11652 29220
rect 11388 29180 11394 29192
rect 11054 29112 11060 29164
rect 11112 29112 11118 29164
rect 11146 29112 11152 29164
rect 11204 29112 11210 29164
rect 11514 29112 11520 29164
rect 11572 29112 11578 29164
rect 11624 29152 11652 29192
rect 12894 29180 12900 29232
rect 12952 29180 12958 29232
rect 14461 29223 14519 29229
rect 14461 29220 14473 29223
rect 13001 29192 14473 29220
rect 11974 29152 11980 29164
rect 11624 29124 11980 29152
rect 11974 29112 11980 29124
rect 12032 29152 12038 29164
rect 12253 29155 12311 29161
rect 12253 29152 12265 29155
rect 12032 29124 12265 29152
rect 12032 29112 12038 29124
rect 12253 29121 12265 29124
rect 12299 29121 12311 29155
rect 12802 29152 12808 29164
rect 12253 29115 12311 29121
rect 12360 29124 12664 29152
rect 12763 29124 12808 29152
rect 11532 29084 11560 29112
rect 10980 29056 11560 29084
rect 12360 29016 12388 29124
rect 12526 29044 12532 29096
rect 12584 29044 12590 29096
rect 12636 29084 12664 29124
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 13001 29084 13029 29192
rect 14461 29189 14473 29192
rect 14507 29189 14519 29223
rect 14461 29183 14519 29189
rect 15930 29180 15936 29232
rect 15988 29220 15994 29232
rect 15988 29192 16344 29220
rect 15988 29180 15994 29192
rect 13446 29112 13452 29164
rect 13504 29112 13510 29164
rect 13630 29112 13636 29164
rect 13688 29112 13694 29164
rect 14185 29155 14243 29161
rect 14185 29121 14197 29155
rect 14231 29121 14243 29155
rect 14185 29115 14243 29121
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 12636 29056 13029 29084
rect 13262 29044 13268 29096
rect 13320 29044 13326 29096
rect 13464 29084 13492 29112
rect 13722 29084 13728 29096
rect 13464 29056 13728 29084
rect 13722 29044 13728 29056
rect 13780 29084 13786 29096
rect 13909 29087 13967 29093
rect 13909 29084 13921 29087
rect 13780 29056 13921 29084
rect 13780 29044 13786 29056
rect 13909 29053 13921 29056
rect 13955 29053 13967 29087
rect 13909 29047 13967 29053
rect 13173 29019 13231 29025
rect 13173 29016 13185 29019
rect 10888 28988 12388 29016
rect 12452 28988 13185 29016
rect 10594 28948 10600 28960
rect 8352 28920 10600 28948
rect 8352 28908 8358 28920
rect 10594 28908 10600 28920
rect 10652 28948 10658 28960
rect 11054 28948 11060 28960
rect 10652 28920 11060 28948
rect 10652 28908 10658 28920
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 11606 28908 11612 28960
rect 11664 28948 11670 28960
rect 12066 28948 12072 28960
rect 11664 28920 12072 28948
rect 11664 28908 11670 28920
rect 12066 28908 12072 28920
rect 12124 28908 12130 28960
rect 12342 28908 12348 28960
rect 12400 28908 12406 28960
rect 12452 28957 12480 28988
rect 13173 28985 13185 28988
rect 13219 28985 13231 29019
rect 13817 29019 13875 29025
rect 13817 29016 13829 29019
rect 13173 28979 13231 28985
rect 13556 28988 13829 29016
rect 13556 28960 13584 28988
rect 13817 28985 13829 28988
rect 13863 28985 13875 29019
rect 14200 29016 14228 29115
rect 14384 29084 14412 29115
rect 14642 29112 14648 29164
rect 14700 29112 14706 29164
rect 14734 29112 14740 29164
rect 14792 29152 14798 29164
rect 14918 29152 14924 29164
rect 14792 29124 14924 29152
rect 14792 29112 14798 29124
rect 14918 29112 14924 29124
rect 14976 29152 14982 29164
rect 15473 29155 15531 29161
rect 15473 29152 15485 29155
rect 14976 29124 15485 29152
rect 14976 29112 14982 29124
rect 15473 29121 15485 29124
rect 15519 29121 15531 29155
rect 15473 29115 15531 29121
rect 15562 29112 15568 29164
rect 15620 29112 15626 29164
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 16316 29152 16344 29192
rect 17034 29180 17040 29232
rect 17092 29220 17098 29232
rect 18414 29220 18420 29232
rect 17092 29192 18420 29220
rect 17092 29180 17098 29192
rect 18414 29180 18420 29192
rect 18472 29180 18478 29232
rect 18892 29220 18920 29248
rect 19260 29220 19288 29248
rect 19812 29220 19840 29260
rect 20714 29248 20720 29260
rect 20772 29248 20778 29300
rect 20806 29248 20812 29300
rect 20864 29248 20870 29300
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 21048 29260 21128 29288
rect 21048 29248 21054 29260
rect 18800 29192 18920 29220
rect 18984 29192 19288 29220
rect 19444 29192 19840 29220
rect 17402 29152 17408 29164
rect 16316 29124 17408 29152
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 17494 29112 17500 29164
rect 17552 29152 17558 29164
rect 18138 29152 18144 29164
rect 17552 29124 18144 29152
rect 17552 29112 17558 29124
rect 18138 29112 18144 29124
rect 18196 29112 18202 29164
rect 18800 29161 18828 29192
rect 18984 29161 19012 29192
rect 18785 29155 18843 29161
rect 18785 29121 18797 29155
rect 18831 29121 18843 29155
rect 18785 29115 18843 29121
rect 18877 29155 18935 29161
rect 18877 29121 18889 29155
rect 18923 29121 18935 29155
rect 18877 29115 18935 29121
rect 18969 29155 19027 29161
rect 18969 29121 18981 29155
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 14826 29084 14832 29096
rect 14384 29056 14832 29084
rect 14826 29044 14832 29056
rect 14884 29084 14890 29096
rect 15580 29084 15608 29112
rect 15657 29087 15715 29093
rect 15657 29084 15669 29087
rect 14884 29056 14964 29084
rect 15580 29056 15669 29084
rect 14884 29044 14890 29056
rect 14734 29016 14740 29028
rect 14200 28988 14740 29016
rect 13817 28979 13875 28985
rect 14734 28976 14740 28988
rect 14792 28976 14798 29028
rect 14936 29016 14964 29056
rect 15657 29053 15669 29056
rect 15703 29053 15715 29087
rect 15657 29047 15715 29053
rect 15838 29044 15844 29096
rect 15896 29044 15902 29096
rect 17310 29044 17316 29096
rect 17368 29084 17374 29096
rect 17770 29084 17776 29096
rect 17368 29056 17776 29084
rect 17368 29044 17374 29056
rect 17770 29044 17776 29056
rect 17828 29044 17834 29096
rect 18892 29084 18920 29115
rect 19150 29112 19156 29164
rect 19208 29112 19214 29164
rect 19444 29152 19472 29192
rect 19812 29161 19840 29192
rect 19904 29192 21036 29220
rect 19904 29161 19932 29192
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 19260 29124 19472 29152
rect 19511 29124 19717 29152
rect 19260 29084 19288 29124
rect 18892 29056 19288 29084
rect 19334 29044 19340 29096
rect 19392 29084 19398 29096
rect 19511 29084 19539 29124
rect 19705 29121 19717 29124
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19797 29155 19855 29161
rect 19797 29121 19809 29155
rect 19843 29121 19855 29155
rect 19797 29115 19855 29121
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29121 19947 29155
rect 19889 29115 19947 29121
rect 19978 29112 19984 29164
rect 20036 29152 20042 29164
rect 20073 29155 20131 29161
rect 20073 29152 20085 29155
rect 20036 29124 20085 29152
rect 20036 29112 20042 29124
rect 20073 29121 20085 29124
rect 20119 29152 20131 29155
rect 20530 29152 20536 29164
rect 20119 29124 20536 29152
rect 20119 29121 20131 29124
rect 20073 29115 20131 29121
rect 19392 29056 19539 29084
rect 19392 29044 19398 29056
rect 19610 29044 19616 29096
rect 19668 29084 19674 29096
rect 20165 29087 20223 29093
rect 20165 29084 20177 29087
rect 19668 29056 20177 29084
rect 19668 29044 19674 29056
rect 20165 29053 20177 29056
rect 20211 29053 20223 29087
rect 20165 29047 20223 29053
rect 19352 29016 19380 29044
rect 20263 29016 20291 29124
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 14936 28988 19380 29016
rect 19444 28988 20291 29016
rect 21008 29016 21036 29192
rect 21100 29161 21128 29260
rect 21174 29248 21180 29300
rect 21232 29248 21238 29300
rect 22738 29288 22744 29300
rect 21376 29260 22744 29288
rect 21192 29220 21220 29248
rect 21192 29192 21312 29220
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21174 29112 21180 29164
rect 21232 29112 21238 29164
rect 21284 29084 21312 29192
rect 21376 29161 21404 29260
rect 22738 29248 22744 29260
rect 22796 29248 22802 29300
rect 23658 29288 23664 29300
rect 22848 29260 23664 29288
rect 22848 29220 22876 29260
rect 23658 29248 23664 29260
rect 23716 29248 23722 29300
rect 23750 29248 23756 29300
rect 23808 29248 23814 29300
rect 23842 29248 23848 29300
rect 23900 29248 23906 29300
rect 24394 29248 24400 29300
rect 24452 29288 24458 29300
rect 24452 29260 25183 29288
rect 24452 29248 24458 29260
rect 22756 29192 22876 29220
rect 22756 29164 22784 29192
rect 23290 29180 23296 29232
rect 23348 29220 23354 29232
rect 23348 29192 23612 29220
rect 23348 29180 23354 29192
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 21450 29112 21456 29164
rect 21508 29161 21514 29164
rect 21508 29155 21521 29161
rect 21509 29152 21521 29155
rect 21509 29124 21553 29152
rect 21509 29121 21521 29124
rect 21508 29115 21521 29121
rect 21508 29112 21514 29115
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 21913 29155 21971 29161
rect 21913 29152 21925 29155
rect 21784 29124 21925 29152
rect 21784 29112 21790 29124
rect 21913 29121 21925 29124
rect 21959 29121 21971 29155
rect 21913 29115 21971 29121
rect 22020 29084 22048 29138
rect 22738 29112 22744 29164
rect 22796 29112 22802 29164
rect 23014 29112 23020 29164
rect 23072 29112 23078 29164
rect 23198 29112 23204 29164
rect 23256 29112 23262 29164
rect 23584 29161 23612 29192
rect 23569 29155 23627 29161
rect 23569 29121 23581 29155
rect 23615 29121 23627 29155
rect 23569 29115 23627 29121
rect 23658 29112 23664 29164
rect 23716 29112 23722 29164
rect 21284 29056 22048 29084
rect 22922 29044 22928 29096
rect 22980 29044 22986 29096
rect 23768 29016 23796 29248
rect 23860 29220 23888 29248
rect 23860 29192 23980 29220
rect 23952 29161 23980 29192
rect 24210 29180 24216 29232
rect 24268 29220 24274 29232
rect 24857 29223 24915 29229
rect 24268 29192 24532 29220
rect 24268 29180 24274 29192
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29152 23995 29155
rect 24302 29152 24308 29164
rect 23983 29124 24308 29152
rect 23983 29121 23995 29124
rect 23937 29115 23995 29121
rect 23860 29084 23888 29115
rect 24302 29112 24308 29124
rect 24360 29112 24366 29164
rect 24504 29161 24532 29192
rect 24857 29189 24869 29223
rect 24903 29220 24915 29223
rect 24946 29220 24952 29232
rect 24903 29192 24952 29220
rect 24903 29189 24915 29192
rect 24857 29183 24915 29189
rect 24946 29180 24952 29192
rect 25004 29180 25010 29232
rect 25155 29220 25183 29260
rect 25222 29248 25228 29300
rect 25280 29288 25286 29300
rect 25498 29288 25504 29300
rect 25280 29260 25504 29288
rect 25280 29248 25286 29260
rect 25498 29248 25504 29260
rect 25556 29288 25562 29300
rect 25685 29291 25743 29297
rect 25685 29288 25697 29291
rect 25556 29260 25697 29288
rect 25556 29248 25562 29260
rect 25685 29257 25697 29260
rect 25731 29257 25743 29291
rect 25685 29251 25743 29257
rect 26970 29248 26976 29300
rect 27028 29248 27034 29300
rect 27522 29288 27528 29300
rect 27172 29260 27528 29288
rect 27062 29220 27068 29232
rect 25155 29192 25360 29220
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24397 29115 24455 29121
rect 24489 29155 24547 29161
rect 24489 29121 24501 29155
rect 24535 29121 24547 29155
rect 24489 29115 24547 29121
rect 24213 29087 24271 29093
rect 24213 29084 24225 29087
rect 23860 29056 24225 29084
rect 24213 29053 24225 29056
rect 24259 29053 24271 29087
rect 24213 29047 24271 29053
rect 21008 28988 23796 29016
rect 24320 29016 24348 29112
rect 24412 29084 24440 29115
rect 24578 29112 24584 29164
rect 24636 29112 24642 29164
rect 24670 29112 24676 29164
rect 24728 29112 24734 29164
rect 25038 29112 25044 29164
rect 25096 29152 25102 29164
rect 25332 29161 25360 29192
rect 25700 29192 27068 29220
rect 25700 29164 25728 29192
rect 27062 29180 27068 29192
rect 27120 29180 27126 29232
rect 25317 29155 25375 29161
rect 25096 29124 25273 29152
rect 25096 29112 25102 29124
rect 24762 29084 24768 29096
rect 24412 29056 24768 29084
rect 24762 29044 24768 29056
rect 24820 29084 24826 29096
rect 25245 29084 25273 29124
rect 25317 29121 25329 29155
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25406 29112 25412 29164
rect 25464 29152 25470 29164
rect 25464 29124 25509 29152
rect 25464 29112 25470 29124
rect 25682 29112 25688 29164
rect 25740 29112 25746 29164
rect 26418 29112 26424 29164
rect 26476 29112 26482 29164
rect 27172 29161 27200 29260
rect 27522 29248 27528 29260
rect 27580 29288 27586 29300
rect 27706 29288 27712 29300
rect 27580 29260 27712 29288
rect 27580 29248 27586 29260
rect 27706 29248 27712 29260
rect 27764 29248 27770 29300
rect 28718 29248 28724 29300
rect 28776 29248 28782 29300
rect 29086 29288 29092 29300
rect 28920 29260 29092 29288
rect 27430 29180 27436 29232
rect 27488 29220 27494 29232
rect 27488 29192 27752 29220
rect 27488 29180 27494 29192
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 27338 29112 27344 29164
rect 27396 29112 27402 29164
rect 27522 29112 27528 29164
rect 27580 29152 27586 29164
rect 27724 29161 27752 29192
rect 27890 29180 27896 29232
rect 27948 29180 27954 29232
rect 27985 29223 28043 29229
rect 27985 29189 27997 29223
rect 28031 29220 28043 29223
rect 28534 29220 28540 29232
rect 28031 29192 28540 29220
rect 28031 29189 28043 29192
rect 27985 29183 28043 29189
rect 27617 29155 27675 29161
rect 27617 29152 27629 29155
rect 27580 29124 27629 29152
rect 27580 29112 27586 29124
rect 27617 29121 27629 29124
rect 27663 29121 27675 29155
rect 27617 29115 27675 29121
rect 27709 29155 27767 29161
rect 27709 29121 27721 29155
rect 27755 29121 27767 29155
rect 27908 29152 27936 29180
rect 28169 29155 28227 29161
rect 28169 29152 28181 29155
rect 27908 29124 28181 29152
rect 27709 29115 27767 29121
rect 28169 29121 28181 29124
rect 28215 29121 28227 29155
rect 28169 29115 28227 29121
rect 26234 29084 26240 29096
rect 24820 29056 25176 29084
rect 25245 29056 26240 29084
rect 24820 29044 24826 29056
rect 25148 29016 25176 29056
rect 26234 29044 26240 29056
rect 26292 29044 26298 29096
rect 26436 29084 26464 29112
rect 27249 29087 27307 29093
rect 27249 29084 27261 29087
rect 26436 29056 27261 29084
rect 27249 29053 27261 29056
rect 27295 29053 27307 29087
rect 27249 29047 27307 29053
rect 27433 29087 27491 29093
rect 27433 29053 27445 29087
rect 27479 29053 27491 29087
rect 28276 29084 28304 29192
rect 28534 29180 28540 29192
rect 28592 29180 28598 29232
rect 28736 29152 28764 29248
rect 28920 29161 28948 29260
rect 29086 29248 29092 29260
rect 29144 29248 29150 29300
rect 29178 29248 29184 29300
rect 29236 29288 29242 29300
rect 29236 29260 29776 29288
rect 29236 29248 29242 29260
rect 29196 29220 29224 29248
rect 29012 29192 29224 29220
rect 29273 29223 29331 29229
rect 29012 29161 29040 29192
rect 29273 29189 29285 29223
rect 29319 29220 29331 29223
rect 29319 29192 29500 29220
rect 29319 29189 29331 29192
rect 29273 29183 29331 29189
rect 29472 29164 29500 29192
rect 28813 29155 28871 29161
rect 28813 29152 28825 29155
rect 28736 29124 28825 29152
rect 28813 29121 28825 29124
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 28905 29155 28963 29161
rect 28905 29121 28917 29155
rect 28951 29121 28963 29155
rect 28905 29115 28963 29121
rect 28997 29155 29055 29161
rect 28997 29121 29009 29155
rect 29043 29121 29055 29155
rect 28997 29115 29055 29121
rect 29086 29112 29092 29164
rect 29144 29152 29150 29164
rect 29181 29155 29239 29161
rect 29181 29152 29193 29155
rect 29144 29124 29193 29152
rect 29144 29112 29150 29124
rect 29181 29121 29193 29124
rect 29227 29121 29239 29155
rect 29181 29115 29239 29121
rect 29362 29112 29368 29164
rect 29420 29112 29426 29164
rect 29454 29112 29460 29164
rect 29512 29112 29518 29164
rect 29546 29112 29552 29164
rect 29604 29152 29610 29164
rect 29748 29161 29776 29260
rect 30374 29248 30380 29300
rect 30432 29288 30438 29300
rect 30469 29291 30527 29297
rect 30469 29288 30481 29291
rect 30432 29260 30481 29288
rect 30432 29248 30438 29260
rect 30469 29257 30481 29260
rect 30515 29257 30527 29291
rect 30469 29251 30527 29257
rect 31570 29248 31576 29300
rect 31628 29248 31634 29300
rect 33226 29248 33232 29300
rect 33284 29288 33290 29300
rect 33597 29291 33655 29297
rect 33597 29288 33609 29291
rect 33284 29260 33609 29288
rect 33284 29248 33290 29260
rect 33597 29257 33609 29260
rect 33643 29288 33655 29291
rect 34517 29291 34575 29297
rect 34517 29288 34529 29291
rect 33643 29260 34529 29288
rect 33643 29257 33655 29260
rect 33597 29251 33655 29257
rect 34517 29257 34529 29260
rect 34563 29257 34575 29291
rect 34517 29251 34575 29257
rect 30834 29180 30840 29232
rect 30892 29180 30898 29232
rect 30929 29223 30987 29229
rect 30929 29189 30941 29223
rect 30975 29220 30987 29223
rect 30975 29192 31432 29220
rect 30975 29189 30987 29192
rect 30929 29183 30987 29189
rect 31404 29164 31432 29192
rect 29641 29155 29699 29161
rect 29641 29152 29653 29155
rect 29604 29124 29653 29152
rect 29604 29112 29610 29124
rect 29641 29121 29653 29124
rect 29687 29121 29699 29155
rect 29641 29115 29699 29121
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 29917 29155 29975 29161
rect 29917 29121 29929 29155
rect 29963 29121 29975 29155
rect 29917 29115 29975 29121
rect 27433 29047 27491 29053
rect 28000 29056 28304 29084
rect 28721 29087 28779 29093
rect 25225 29019 25283 29025
rect 25225 29016 25237 29019
rect 24320 28988 24532 29016
rect 25148 28988 25237 29016
rect 12437 28951 12495 28957
rect 12437 28917 12449 28951
rect 12483 28917 12495 28951
rect 12437 28911 12495 28917
rect 12526 28908 12532 28960
rect 12584 28948 12590 28960
rect 12986 28948 12992 28960
rect 12584 28920 12992 28948
rect 12584 28908 12590 28920
rect 12986 28908 12992 28920
rect 13044 28908 13050 28960
rect 13446 28908 13452 28960
rect 13504 28908 13510 28960
rect 13538 28908 13544 28960
rect 13596 28908 13602 28960
rect 17678 28908 17684 28960
rect 17736 28948 17742 28960
rect 19058 28948 19064 28960
rect 17736 28920 19064 28948
rect 17736 28908 17742 28920
rect 19058 28908 19064 28920
rect 19116 28908 19122 28960
rect 19150 28908 19156 28960
rect 19208 28948 19214 28960
rect 19444 28948 19472 28988
rect 19208 28920 19472 28948
rect 19208 28908 19214 28920
rect 20530 28908 20536 28960
rect 20588 28948 20594 28960
rect 20901 28951 20959 28957
rect 20901 28948 20913 28951
rect 20588 28920 20913 28948
rect 20588 28908 20594 28920
rect 20901 28917 20913 28920
rect 20947 28917 20959 28951
rect 20901 28911 20959 28917
rect 22646 28908 22652 28960
rect 22704 28948 22710 28960
rect 23017 28951 23075 28957
rect 23017 28948 23029 28951
rect 22704 28920 23029 28948
rect 22704 28908 22710 28920
rect 23017 28917 23029 28920
rect 23063 28917 23075 28951
rect 23017 28911 23075 28917
rect 23385 28951 23443 28957
rect 23385 28917 23397 28951
rect 23431 28948 23443 28951
rect 24394 28948 24400 28960
rect 23431 28920 24400 28948
rect 23431 28917 23443 28920
rect 23385 28911 23443 28917
rect 24394 28908 24400 28920
rect 24452 28908 24458 28960
rect 24504 28948 24532 28988
rect 25225 28985 25237 28988
rect 25271 29016 25283 29019
rect 27448 29016 27476 29047
rect 27801 29019 27859 29025
rect 27801 29016 27813 29019
rect 25271 28988 27384 29016
rect 27448 28988 27813 29016
rect 25271 28985 25283 28988
rect 25225 28979 25283 28985
rect 25961 28951 26019 28957
rect 25961 28948 25973 28951
rect 24504 28920 25973 28948
rect 25961 28917 25973 28920
rect 26007 28917 26019 28951
rect 27356 28948 27384 28988
rect 27801 28985 27813 28988
rect 27847 29016 27859 29019
rect 27890 29016 27896 29028
rect 27847 28988 27896 29016
rect 27847 28985 27859 28988
rect 27801 28979 27859 28985
rect 27890 28976 27896 28988
rect 27948 28976 27954 29028
rect 28000 28948 28028 29056
rect 28721 29053 28733 29087
rect 28767 29053 28779 29087
rect 28721 29047 28779 29053
rect 28074 28976 28080 29028
rect 28132 29016 28138 29028
rect 28353 29019 28411 29025
rect 28353 29016 28365 29019
rect 28132 28988 28365 29016
rect 28132 28976 28138 28988
rect 28353 28985 28365 28988
rect 28399 29016 28411 29019
rect 28399 28988 28488 29016
rect 28399 28985 28411 28988
rect 28353 28979 28411 28985
rect 27356 28920 28028 28948
rect 28460 28948 28488 28988
rect 28534 28976 28540 29028
rect 28592 28976 28598 29028
rect 28626 28976 28632 29028
rect 28684 29016 28690 29028
rect 28736 29016 28764 29047
rect 29270 29044 29276 29096
rect 29328 29084 29334 29096
rect 29932 29084 29960 29115
rect 30282 29112 30288 29164
rect 30340 29112 30346 29164
rect 30558 29112 30564 29164
rect 30616 29152 30622 29164
rect 30653 29155 30711 29161
rect 30653 29152 30665 29155
rect 30616 29124 30665 29152
rect 30616 29112 30622 29124
rect 30653 29121 30665 29124
rect 30699 29121 30711 29155
rect 30653 29115 30711 29121
rect 31018 29112 31024 29164
rect 31076 29112 31082 29164
rect 31110 29112 31116 29164
rect 31168 29112 31174 29164
rect 31297 29155 31355 29161
rect 31297 29121 31309 29155
rect 31343 29121 31355 29155
rect 31297 29115 31355 29121
rect 29328 29056 29960 29084
rect 29328 29044 29334 29056
rect 30098 29044 30104 29096
rect 30156 29044 30162 29096
rect 30300 29084 30328 29112
rect 31128 29084 31156 29112
rect 30300 29056 31156 29084
rect 31312 29084 31340 29115
rect 31386 29112 31392 29164
rect 31444 29112 31450 29164
rect 31588 29152 31616 29248
rect 31662 29180 31668 29232
rect 31720 29220 31726 29232
rect 31941 29223 31999 29229
rect 31941 29220 31953 29223
rect 31720 29192 31953 29220
rect 31720 29180 31726 29192
rect 31941 29189 31953 29192
rect 31987 29189 31999 29223
rect 31941 29183 31999 29189
rect 32953 29223 33011 29229
rect 32953 29189 32965 29223
rect 32999 29220 33011 29223
rect 33244 29220 33272 29248
rect 32999 29192 33272 29220
rect 32999 29189 33011 29192
rect 32953 29183 33011 29189
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31588 29124 32137 29152
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 33410 29152 33416 29164
rect 32125 29115 32183 29121
rect 32600 29124 33416 29152
rect 32600 29084 32628 29124
rect 33410 29112 33416 29124
rect 33468 29112 33474 29164
rect 33505 29155 33563 29161
rect 33505 29121 33517 29155
rect 33551 29152 33563 29155
rect 33551 29124 34100 29152
rect 33551 29121 33563 29124
rect 33505 29115 33563 29121
rect 33042 29084 33048 29096
rect 31312 29056 32628 29084
rect 32692 29056 33048 29084
rect 28684 28988 28764 29016
rect 28684 28976 28690 28988
rect 29638 28976 29644 29028
rect 29696 29016 29702 29028
rect 29733 29019 29791 29025
rect 29733 29016 29745 29019
rect 29696 28988 29745 29016
rect 29696 28976 29702 28988
rect 29733 28985 29745 28988
rect 29779 28985 29791 29019
rect 29733 28979 29791 28985
rect 30650 28976 30656 29028
rect 30708 28976 30714 29028
rect 31205 29019 31263 29025
rect 31205 28985 31217 29019
rect 31251 29016 31263 29019
rect 32692 29016 32720 29056
rect 33042 29044 33048 29056
rect 33100 29044 33106 29096
rect 34072 29028 34100 29124
rect 31251 28988 32720 29016
rect 32769 29019 32827 29025
rect 31251 28985 31263 28988
rect 31205 28979 31263 28985
rect 32769 28985 32781 29019
rect 32815 29016 32827 29019
rect 33686 29016 33692 29028
rect 32815 28988 33692 29016
rect 32815 28985 32827 28988
rect 32769 28979 32827 28985
rect 33686 28976 33692 28988
rect 33744 28976 33750 29028
rect 34054 28976 34060 29028
rect 34112 29016 34118 29028
rect 34149 29019 34207 29025
rect 34149 29016 34161 29019
rect 34112 28988 34161 29016
rect 34112 28976 34118 28988
rect 34149 28985 34161 28988
rect 34195 28985 34207 29019
rect 34149 28979 34207 28985
rect 28902 28948 28908 28960
rect 28460 28920 28908 28948
rect 25961 28911 26019 28917
rect 28902 28908 28908 28920
rect 28960 28908 28966 28960
rect 29457 28951 29515 28957
rect 29457 28917 29469 28951
rect 29503 28948 29515 28951
rect 30558 28948 30564 28960
rect 29503 28920 30564 28948
rect 29503 28917 29515 28920
rect 29457 28911 29515 28917
rect 30558 28908 30564 28920
rect 30616 28908 30622 28960
rect 30668 28948 30696 28976
rect 33045 28951 33103 28957
rect 33045 28948 33057 28951
rect 30668 28920 33057 28948
rect 33045 28917 33057 28920
rect 33091 28948 33103 28951
rect 33502 28948 33508 28960
rect 33091 28920 33508 28948
rect 33091 28917 33103 28920
rect 33045 28911 33103 28917
rect 33502 28908 33508 28920
rect 33560 28908 33566 28960
rect 1104 28858 43884 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 43884 28858
rect 1104 28784 43884 28806
rect 2498 28704 2504 28756
rect 2556 28744 2562 28756
rect 2869 28747 2927 28753
rect 2869 28744 2881 28747
rect 2556 28716 2881 28744
rect 2556 28704 2562 28716
rect 2869 28713 2881 28716
rect 2915 28744 2927 28747
rect 3418 28744 3424 28756
rect 2915 28716 3424 28744
rect 2915 28713 2927 28716
rect 2869 28707 2927 28713
rect 3418 28704 3424 28716
rect 3476 28704 3482 28756
rect 3694 28704 3700 28756
rect 3752 28704 3758 28756
rect 3970 28704 3976 28756
rect 4028 28704 4034 28756
rect 4985 28747 5043 28753
rect 4985 28744 4997 28747
rect 4172 28716 4997 28744
rect 3712 28676 3740 28704
rect 4172 28676 4200 28716
rect 4985 28713 4997 28716
rect 5031 28713 5043 28747
rect 4985 28707 5043 28713
rect 3712 28648 4200 28676
rect 5000 28676 5028 28707
rect 5074 28704 5080 28756
rect 5132 28744 5138 28756
rect 5442 28744 5448 28756
rect 5132 28716 5448 28744
rect 5132 28704 5138 28716
rect 5442 28704 5448 28716
rect 5500 28704 5506 28756
rect 5626 28704 5632 28756
rect 5684 28744 5690 28756
rect 6181 28747 6239 28753
rect 6181 28744 6193 28747
rect 5684 28716 6193 28744
rect 5684 28704 5690 28716
rect 6181 28713 6193 28716
rect 6227 28713 6239 28747
rect 6181 28707 6239 28713
rect 7101 28747 7159 28753
rect 7101 28713 7113 28747
rect 7147 28744 7159 28747
rect 7190 28744 7196 28756
rect 7147 28716 7196 28744
rect 7147 28713 7159 28716
rect 7101 28707 7159 28713
rect 7190 28704 7196 28716
rect 7248 28704 7254 28756
rect 7834 28704 7840 28756
rect 7892 28704 7898 28756
rect 9306 28704 9312 28756
rect 9364 28744 9370 28756
rect 9769 28747 9827 28753
rect 9769 28744 9781 28747
rect 9364 28716 9781 28744
rect 9364 28704 9370 28716
rect 9769 28713 9781 28716
rect 9815 28713 9827 28747
rect 9769 28707 9827 28713
rect 9950 28704 9956 28756
rect 10008 28704 10014 28756
rect 10318 28704 10324 28756
rect 10376 28744 10382 28756
rect 11057 28747 11115 28753
rect 11057 28744 11069 28747
rect 10376 28716 11069 28744
rect 10376 28704 10382 28716
rect 11057 28713 11069 28716
rect 11103 28713 11115 28747
rect 11057 28707 11115 28713
rect 11146 28704 11152 28756
rect 11204 28744 11210 28756
rect 11333 28747 11391 28753
rect 11333 28744 11345 28747
rect 11204 28716 11345 28744
rect 11204 28704 11210 28716
rect 11333 28713 11345 28716
rect 11379 28713 11391 28747
rect 11333 28707 11391 28713
rect 11514 28704 11520 28756
rect 11572 28704 11578 28756
rect 11974 28704 11980 28756
rect 12032 28704 12038 28756
rect 12342 28704 12348 28756
rect 12400 28744 12406 28756
rect 12710 28744 12716 28756
rect 12400 28716 12716 28744
rect 12400 28704 12406 28716
rect 12710 28704 12716 28716
rect 12768 28704 12774 28756
rect 12805 28747 12863 28753
rect 12805 28713 12817 28747
rect 12851 28744 12863 28747
rect 13262 28744 13268 28756
rect 12851 28716 13268 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 13262 28704 13268 28716
rect 13320 28704 13326 28756
rect 13354 28704 13360 28756
rect 13412 28704 13418 28756
rect 14182 28704 14188 28756
rect 14240 28744 14246 28756
rect 14369 28747 14427 28753
rect 14369 28744 14381 28747
rect 14240 28716 14381 28744
rect 14240 28704 14246 28716
rect 14369 28713 14381 28716
rect 14415 28744 14427 28747
rect 14826 28744 14832 28756
rect 14415 28716 14832 28744
rect 14415 28713 14427 28716
rect 14369 28707 14427 28713
rect 14826 28704 14832 28716
rect 14884 28704 14890 28756
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 17405 28747 17463 28753
rect 17405 28744 17417 28747
rect 17368 28716 17417 28744
rect 17368 28704 17374 28716
rect 17405 28713 17417 28716
rect 17451 28713 17463 28747
rect 17954 28744 17960 28756
rect 17405 28707 17463 28713
rect 17696 28716 17960 28744
rect 5000 28648 5672 28676
rect 1210 28568 1216 28620
rect 1268 28608 1274 28620
rect 1857 28611 1915 28617
rect 1857 28608 1869 28611
rect 1268 28580 1869 28608
rect 1268 28568 1274 28580
rect 1857 28577 1869 28580
rect 1903 28577 1915 28611
rect 1857 28571 1915 28577
rect 3786 28568 3792 28620
rect 3844 28568 3850 28620
rect 4338 28568 4344 28620
rect 4396 28608 4402 28620
rect 4396 28580 5396 28608
rect 4396 28568 4402 28580
rect 1578 28500 1584 28552
rect 1636 28500 1642 28552
rect 2590 28500 2596 28552
rect 2648 28540 2654 28552
rect 3050 28540 3056 28552
rect 2648 28512 3056 28540
rect 2648 28500 2654 28512
rect 3050 28500 3056 28512
rect 3108 28500 3114 28552
rect 3329 28543 3387 28549
rect 3329 28509 3341 28543
rect 3375 28540 3387 28543
rect 3804 28540 3832 28568
rect 3375 28512 3464 28540
rect 3804 28512 4032 28540
rect 3375 28509 3387 28512
rect 3329 28503 3387 28509
rect 3436 28484 3464 28512
rect 2746 28444 3372 28472
rect 1854 28364 1860 28416
rect 1912 28404 1918 28416
rect 2746 28404 2774 28444
rect 1912 28376 2774 28404
rect 1912 28364 1918 28376
rect 3234 28364 3240 28416
rect 3292 28364 3298 28416
rect 3344 28404 3372 28444
rect 3418 28432 3424 28484
rect 3476 28432 3482 28484
rect 3786 28432 3792 28484
rect 3844 28432 3850 28484
rect 4004 28472 4032 28512
rect 5031 28509 5089 28515
rect 4430 28472 4436 28484
rect 4004 28444 4436 28472
rect 4430 28432 4436 28444
rect 4488 28432 4494 28484
rect 4801 28475 4859 28481
rect 4801 28441 4813 28475
rect 4847 28472 4859 28475
rect 4890 28472 4896 28484
rect 4847 28444 4896 28472
rect 4847 28441 4859 28444
rect 4801 28435 4859 28441
rect 4890 28432 4896 28444
rect 4948 28432 4954 28484
rect 5031 28475 5043 28509
rect 5077 28475 5089 28509
rect 5031 28472 5089 28475
rect 5031 28469 5120 28472
rect 5046 28444 5120 28469
rect 5092 28416 5120 28444
rect 5258 28432 5264 28484
rect 5316 28432 5322 28484
rect 5368 28472 5396 28580
rect 5442 28500 5448 28552
rect 5500 28500 5506 28552
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5644 28540 5672 28648
rect 5810 28636 5816 28688
rect 5868 28676 5874 28688
rect 10502 28676 10508 28688
rect 5868 28648 10508 28676
rect 5868 28636 5874 28648
rect 6362 28568 6368 28620
rect 6420 28568 6426 28620
rect 6546 28568 6552 28620
rect 6604 28608 6610 28620
rect 6730 28608 6736 28620
rect 6604 28580 6736 28608
rect 6604 28568 6610 28580
rect 6730 28568 6736 28580
rect 6788 28568 6794 28620
rect 5592 28512 5672 28540
rect 5592 28500 5598 28512
rect 5810 28500 5816 28552
rect 5868 28540 5874 28552
rect 5905 28543 5963 28549
rect 5905 28540 5917 28543
rect 5868 28512 5917 28540
rect 5868 28500 5874 28512
rect 5905 28509 5917 28512
rect 5951 28540 5963 28543
rect 6380 28540 6408 28568
rect 7300 28549 7328 28648
rect 8220 28549 8248 28648
rect 10502 28636 10508 28648
rect 10560 28636 10566 28688
rect 11241 28679 11299 28685
rect 11241 28645 11253 28679
rect 11287 28676 11299 28679
rect 11532 28676 11560 28704
rect 11287 28648 11560 28676
rect 11992 28676 12020 28704
rect 14737 28679 14795 28685
rect 14737 28676 14749 28679
rect 11992 28648 12434 28676
rect 11287 28645 11299 28648
rect 11241 28639 11299 28645
rect 8294 28568 8300 28620
rect 8352 28568 8358 28620
rect 8481 28611 8539 28617
rect 8481 28577 8493 28611
rect 8527 28608 8539 28611
rect 8662 28608 8668 28620
rect 8527 28580 8668 28608
rect 8527 28577 8539 28580
rect 8481 28571 8539 28577
rect 8662 28568 8668 28580
rect 8720 28568 8726 28620
rect 9582 28568 9588 28620
rect 9640 28608 9646 28620
rect 11977 28611 12035 28617
rect 11977 28608 11989 28611
rect 9640 28580 11989 28608
rect 9640 28568 9646 28580
rect 11977 28577 11989 28580
rect 12023 28608 12035 28611
rect 12158 28608 12164 28620
rect 12023 28580 12164 28608
rect 12023 28577 12035 28580
rect 11977 28571 12035 28577
rect 12158 28568 12164 28580
rect 12216 28568 12222 28620
rect 5951 28512 6408 28540
rect 7101 28543 7159 28549
rect 5951 28509 5963 28512
rect 5905 28503 5963 28509
rect 7101 28509 7113 28543
rect 7147 28509 7159 28543
rect 7101 28503 7159 28509
rect 7285 28543 7343 28549
rect 7285 28509 7297 28543
rect 7331 28509 7343 28543
rect 7285 28503 7343 28509
rect 8205 28543 8263 28549
rect 8205 28509 8217 28543
rect 8251 28509 8263 28543
rect 8205 28503 8263 28509
rect 6086 28472 6092 28484
rect 5368 28444 6092 28472
rect 6086 28432 6092 28444
rect 6144 28472 6150 28484
rect 6730 28472 6736 28484
rect 6144 28444 6736 28472
rect 6144 28432 6150 28444
rect 6730 28432 6736 28444
rect 6788 28432 6794 28484
rect 7116 28472 7144 28503
rect 7190 28472 7196 28484
rect 7116 28444 7196 28472
rect 7190 28432 7196 28444
rect 7248 28432 7254 28484
rect 3989 28407 4047 28413
rect 3989 28404 4001 28407
rect 3344 28376 4001 28404
rect 3989 28373 4001 28376
rect 4035 28373 4047 28407
rect 3989 28367 4047 28373
rect 4154 28364 4160 28416
rect 4212 28404 4218 28416
rect 4982 28404 4988 28416
rect 4212 28376 4988 28404
rect 4212 28364 4218 28376
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 5074 28364 5080 28416
rect 5132 28364 5138 28416
rect 5166 28364 5172 28416
rect 5224 28364 5230 28416
rect 5350 28364 5356 28416
rect 5408 28413 5414 28416
rect 5408 28367 5417 28413
rect 5408 28364 5414 28367
rect 5626 28364 5632 28416
rect 5684 28404 5690 28416
rect 7558 28404 7564 28416
rect 5684 28376 7564 28404
rect 5684 28364 5690 28376
rect 7558 28364 7564 28376
rect 7616 28404 7622 28416
rect 8312 28404 8340 28568
rect 9214 28500 9220 28552
rect 9272 28540 9278 28552
rect 9272 28515 9858 28540
rect 9272 28512 9873 28515
rect 9272 28500 9278 28512
rect 9815 28509 9873 28512
rect 8938 28432 8944 28484
rect 8996 28472 9002 28484
rect 9585 28475 9643 28481
rect 9585 28472 9597 28475
rect 8996 28444 9597 28472
rect 8996 28432 9002 28444
rect 9585 28441 9597 28444
rect 9631 28472 9643 28475
rect 9674 28472 9680 28484
rect 9631 28444 9680 28472
rect 9631 28441 9643 28444
rect 9585 28435 9643 28441
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 9815 28475 9827 28509
rect 9861 28475 9873 28509
rect 10778 28500 10784 28552
rect 10836 28500 10842 28552
rect 12406 28540 12434 28648
rect 12636 28648 14749 28676
rect 12636 28620 12664 28648
rect 14737 28645 14749 28648
rect 14783 28676 14795 28679
rect 15105 28679 15163 28685
rect 15105 28676 15117 28679
rect 14783 28648 15117 28676
rect 14783 28645 14795 28648
rect 14737 28639 14795 28645
rect 15105 28645 15117 28648
rect 15151 28676 15163 28679
rect 15838 28676 15844 28688
rect 15151 28648 15844 28676
rect 15151 28645 15163 28648
rect 15105 28639 15163 28645
rect 15838 28636 15844 28648
rect 15896 28636 15902 28688
rect 12618 28568 12624 28620
rect 12676 28568 12682 28620
rect 12713 28611 12771 28617
rect 12713 28577 12725 28611
rect 12759 28608 12771 28611
rect 12759 28580 13400 28608
rect 12759 28577 12771 28580
rect 12713 28571 12771 28577
rect 12986 28543 13044 28549
rect 12986 28540 12998 28543
rect 12406 28512 12998 28540
rect 12986 28509 12998 28512
rect 13032 28540 13044 28543
rect 13372 28540 13400 28580
rect 13446 28568 13452 28620
rect 13504 28568 13510 28620
rect 13032 28512 13124 28540
rect 13372 28512 13676 28540
rect 13032 28509 13044 28512
rect 12986 28503 13044 28509
rect 9815 28469 9873 28475
rect 7616 28376 8340 28404
rect 10796 28404 10824 28500
rect 10873 28475 10931 28481
rect 10873 28441 10885 28475
rect 10919 28472 10931 28475
rect 11238 28472 11244 28484
rect 10919 28444 11244 28472
rect 10919 28441 10931 28444
rect 10873 28435 10931 28441
rect 11238 28432 11244 28444
rect 11296 28432 11302 28484
rect 11882 28432 11888 28484
rect 11940 28472 11946 28484
rect 12526 28472 12532 28484
rect 11940 28444 12532 28472
rect 11940 28432 11946 28444
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 11073 28407 11131 28413
rect 11073 28404 11085 28407
rect 10796 28376 11085 28404
rect 7616 28364 7622 28376
rect 11073 28373 11085 28376
rect 11119 28373 11131 28407
rect 11073 28367 11131 28373
rect 11606 28364 11612 28416
rect 11664 28404 11670 28416
rect 11701 28407 11759 28413
rect 11701 28404 11713 28407
rect 11664 28376 11713 28404
rect 11664 28364 11670 28376
rect 11701 28373 11713 28376
rect 11747 28373 11759 28407
rect 11701 28367 11759 28373
rect 11790 28364 11796 28416
rect 11848 28364 11854 28416
rect 12986 28364 12992 28416
rect 13044 28364 13050 28416
rect 13096 28404 13124 28512
rect 13446 28432 13452 28484
rect 13504 28472 13510 28484
rect 13541 28475 13599 28481
rect 13541 28472 13553 28475
rect 13504 28444 13553 28472
rect 13504 28432 13510 28444
rect 13541 28441 13553 28444
rect 13587 28441 13599 28475
rect 13648 28472 13676 28512
rect 13722 28500 13728 28552
rect 13780 28500 13786 28552
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16758 28540 16764 28552
rect 16071 28512 16764 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 17310 28500 17316 28552
rect 17368 28540 17374 28552
rect 17589 28543 17647 28549
rect 17589 28540 17601 28543
rect 17368 28512 17601 28540
rect 17368 28500 17374 28512
rect 17589 28509 17601 28512
rect 17635 28509 17647 28543
rect 17696 28540 17724 28716
rect 17954 28704 17960 28716
rect 18012 28704 18018 28756
rect 18141 28747 18199 28753
rect 18141 28713 18153 28747
rect 18187 28744 18199 28747
rect 19705 28747 19763 28753
rect 18187 28716 18258 28744
rect 18187 28713 18199 28716
rect 18141 28707 18199 28713
rect 17862 28636 17868 28688
rect 17920 28636 17926 28688
rect 18230 28676 18258 28716
rect 19705 28713 19717 28747
rect 19751 28744 19763 28747
rect 20162 28744 20168 28756
rect 19751 28716 20168 28744
rect 19751 28713 19763 28716
rect 19705 28707 19763 28713
rect 20162 28704 20168 28716
rect 20220 28704 20226 28756
rect 20257 28747 20315 28753
rect 20257 28713 20269 28747
rect 20303 28744 20315 28747
rect 20303 28716 23060 28744
rect 20303 28713 20315 28716
rect 20257 28707 20315 28713
rect 18598 28676 18604 28688
rect 18230 28648 18604 28676
rect 18598 28636 18604 28648
rect 18656 28636 18662 28688
rect 18966 28636 18972 28688
rect 19024 28676 19030 28688
rect 19613 28679 19671 28685
rect 19613 28676 19625 28679
rect 19024 28648 19625 28676
rect 19024 28636 19030 28648
rect 19613 28645 19625 28648
rect 19659 28645 19671 28679
rect 19613 28639 19671 28645
rect 19794 28636 19800 28688
rect 19852 28636 19858 28688
rect 19886 28636 19892 28688
rect 19944 28676 19950 28688
rect 23032 28676 23060 28716
rect 23198 28704 23204 28756
rect 23256 28704 23262 28756
rect 23658 28704 23664 28756
rect 23716 28744 23722 28756
rect 23937 28747 23995 28753
rect 23937 28744 23949 28747
rect 23716 28716 23949 28744
rect 23716 28704 23722 28716
rect 23937 28713 23949 28716
rect 23983 28713 23995 28747
rect 23937 28707 23995 28713
rect 24118 28704 24124 28756
rect 24176 28704 24182 28756
rect 24394 28704 24400 28756
rect 24452 28704 24458 28756
rect 26418 28704 26424 28756
rect 26476 28704 26482 28756
rect 26878 28704 26884 28756
rect 26936 28744 26942 28756
rect 27065 28747 27123 28753
rect 27065 28744 27077 28747
rect 26936 28716 27077 28744
rect 26936 28704 26942 28716
rect 27065 28713 27077 28716
rect 27111 28744 27123 28747
rect 27154 28744 27160 28756
rect 27111 28716 27160 28744
rect 27111 28713 27123 28716
rect 27065 28707 27123 28713
rect 27154 28704 27160 28716
rect 27212 28704 27218 28756
rect 27249 28747 27307 28753
rect 27249 28713 27261 28747
rect 27295 28744 27307 28747
rect 27522 28744 27528 28756
rect 27295 28716 27528 28744
rect 27295 28713 27307 28716
rect 27249 28707 27307 28713
rect 27522 28704 27528 28716
rect 27580 28704 27586 28756
rect 28718 28744 28724 28756
rect 27632 28716 28724 28744
rect 24136 28676 24164 28704
rect 19944 28648 20668 28676
rect 23032 28648 24164 28676
rect 19944 28636 19950 28648
rect 17880 28608 17908 28636
rect 20640 28617 20668 28648
rect 18877 28611 18935 28617
rect 18877 28608 18889 28611
rect 17880 28580 18889 28608
rect 18877 28577 18889 28580
rect 18923 28577 18935 28611
rect 20625 28611 20683 28617
rect 18877 28571 18935 28577
rect 18984 28580 20024 28608
rect 18984 28552 19012 28580
rect 17773 28543 17831 28549
rect 17773 28540 17785 28543
rect 17696 28512 17785 28540
rect 17589 28503 17647 28509
rect 17773 28509 17785 28512
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 17957 28543 18015 28549
rect 17957 28509 17969 28543
rect 18003 28534 18015 28543
rect 18325 28543 18383 28549
rect 18003 28509 18024 28534
rect 17957 28503 18024 28509
rect 18325 28509 18337 28543
rect 18371 28540 18383 28543
rect 18598 28540 18604 28552
rect 18371 28512 18604 28540
rect 18371 28509 18383 28512
rect 18325 28503 18383 28509
rect 14366 28472 14372 28484
rect 13648 28444 14372 28472
rect 13541 28435 13599 28441
rect 14108 28416 14136 28444
rect 14366 28432 14372 28444
rect 14424 28432 14430 28484
rect 15473 28475 15531 28481
rect 15473 28472 15485 28475
rect 15304 28444 15485 28472
rect 15304 28416 15332 28444
rect 15473 28441 15485 28444
rect 15519 28441 15531 28475
rect 15473 28435 15531 28441
rect 16292 28475 16350 28481
rect 16292 28441 16304 28475
rect 16338 28472 16350 28475
rect 16482 28472 16488 28484
rect 16338 28444 16488 28472
rect 16338 28441 16350 28444
rect 16292 28435 16350 28441
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 17865 28475 17923 28481
rect 17865 28441 17877 28475
rect 17911 28441 17923 28475
rect 17996 28472 18024 28503
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 18966 28500 18972 28552
rect 19024 28500 19030 28552
rect 19058 28500 19064 28552
rect 19116 28500 19122 28552
rect 19150 28500 19156 28552
rect 19208 28540 19214 28552
rect 19996 28549 20024 28580
rect 20625 28577 20637 28611
rect 20671 28577 20683 28611
rect 20625 28571 20683 28577
rect 20806 28568 20812 28620
rect 20864 28608 20870 28620
rect 24412 28617 24440 28704
rect 26602 28676 26608 28688
rect 25976 28648 26608 28676
rect 24397 28611 24455 28617
rect 20864 28580 21404 28608
rect 20864 28568 20870 28580
rect 19521 28543 19579 28549
rect 19521 28540 19533 28543
rect 19208 28512 19533 28540
rect 19208 28500 19214 28512
rect 19521 28509 19533 28512
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28509 20039 28543
rect 19981 28503 20039 28509
rect 18138 28472 18144 28484
rect 17996 28444 18144 28472
rect 17865 28435 17923 28441
rect 13909 28407 13967 28413
rect 13909 28404 13921 28407
rect 13096 28376 13921 28404
rect 13909 28373 13921 28376
rect 13955 28373 13967 28407
rect 13909 28367 13967 28373
rect 14090 28364 14096 28416
rect 14148 28364 14154 28416
rect 15286 28364 15292 28416
rect 15344 28364 15350 28416
rect 15930 28364 15936 28416
rect 15988 28404 15994 28416
rect 16942 28404 16948 28416
rect 15988 28376 16948 28404
rect 15988 28364 15994 28376
rect 16942 28364 16948 28376
rect 17000 28404 17006 28416
rect 17494 28404 17500 28416
rect 17000 28376 17500 28404
rect 17000 28364 17006 28376
rect 17494 28364 17500 28376
rect 17552 28364 17558 28416
rect 17880 28404 17908 28435
rect 18138 28432 18144 28444
rect 18196 28472 18202 28484
rect 19076 28472 19104 28500
rect 18196 28444 19104 28472
rect 19536 28472 19564 28503
rect 20070 28500 20076 28552
rect 20128 28500 20134 28552
rect 20162 28500 20168 28552
rect 20220 28500 20226 28552
rect 20346 28500 20352 28552
rect 20404 28500 20410 28552
rect 21269 28543 21327 28549
rect 21269 28540 21281 28543
rect 20916 28512 21281 28540
rect 20364 28472 20392 28500
rect 19536 28444 20392 28472
rect 18196 28432 18202 28444
rect 20916 28416 20944 28512
rect 21269 28509 21281 28512
rect 21315 28509 21327 28543
rect 21376 28540 21404 28580
rect 24397 28577 24409 28611
rect 24443 28577 24455 28611
rect 24397 28571 24455 28577
rect 25976 28549 26004 28648
rect 26602 28636 26608 28648
rect 26660 28636 26666 28688
rect 27338 28636 27344 28688
rect 27396 28636 27402 28688
rect 26234 28568 26240 28620
rect 26292 28608 26298 28620
rect 26878 28608 26884 28620
rect 26292 28580 26884 28608
rect 26292 28568 26298 28580
rect 26878 28568 26884 28580
rect 26936 28568 26942 28620
rect 23385 28543 23443 28549
rect 23385 28540 23397 28543
rect 21376 28512 23397 28540
rect 21269 28503 21327 28509
rect 23385 28509 23397 28512
rect 23431 28540 23443 28543
rect 25961 28543 26019 28549
rect 23431 28512 24348 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 21514 28475 21572 28481
rect 21514 28472 21526 28475
rect 21376 28444 21526 28472
rect 19150 28404 19156 28416
rect 17880 28376 19156 28404
rect 19150 28364 19156 28376
rect 19208 28364 19214 28416
rect 19245 28407 19303 28413
rect 19245 28373 19257 28407
rect 19291 28404 19303 28407
rect 19417 28404 19423 28416
rect 19291 28376 19423 28404
rect 19291 28373 19303 28376
rect 19245 28367 19303 28373
rect 19417 28364 19423 28376
rect 19475 28364 19481 28416
rect 20438 28364 20444 28416
rect 20496 28364 20502 28416
rect 20898 28364 20904 28416
rect 20956 28364 20962 28416
rect 21177 28407 21235 28413
rect 21177 28373 21189 28407
rect 21223 28404 21235 28407
rect 21376 28404 21404 28444
rect 21514 28441 21526 28444
rect 21560 28441 21572 28475
rect 21514 28435 21572 28441
rect 24320 28416 24348 28512
rect 25961 28509 25973 28543
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 26145 28543 26203 28549
rect 26145 28509 26157 28543
rect 26191 28509 26203 28543
rect 26145 28503 26203 28509
rect 25682 28432 25688 28484
rect 25740 28472 25746 28484
rect 26160 28472 26188 28503
rect 26694 28500 26700 28552
rect 26752 28540 26758 28552
rect 27356 28549 27384 28636
rect 27430 28568 27436 28620
rect 27488 28608 27494 28620
rect 27488 28580 27568 28608
rect 27488 28568 27494 28580
rect 27540 28549 27568 28580
rect 27632 28549 27660 28716
rect 28718 28704 28724 28716
rect 28776 28704 28782 28756
rect 28810 28704 28816 28756
rect 28868 28744 28874 28756
rect 28868 28716 29868 28744
rect 28868 28704 28874 28716
rect 28258 28636 28264 28688
rect 28316 28676 28322 28688
rect 28353 28679 28411 28685
rect 28353 28676 28365 28679
rect 28316 28648 28365 28676
rect 28316 28636 28322 28648
rect 28353 28645 28365 28648
rect 28399 28676 28411 28679
rect 28994 28676 29000 28688
rect 28399 28648 29000 28676
rect 28399 28645 28411 28648
rect 28353 28639 28411 28645
rect 28994 28636 29000 28648
rect 29052 28636 29058 28688
rect 29840 28685 29868 28716
rect 31110 28704 31116 28756
rect 31168 28744 31174 28756
rect 32950 28744 32956 28756
rect 31168 28716 32956 28744
rect 31168 28704 31174 28716
rect 32950 28704 32956 28716
rect 33008 28704 33014 28756
rect 33410 28704 33416 28756
rect 33468 28704 33474 28756
rect 43530 28704 43536 28756
rect 43588 28704 43594 28756
rect 29825 28679 29883 28685
rect 29825 28645 29837 28679
rect 29871 28645 29883 28679
rect 29825 28639 29883 28645
rect 42150 28636 42156 28688
rect 42208 28636 42214 28688
rect 43548 28676 43576 28704
rect 42812 28648 43576 28676
rect 28534 28568 28540 28620
rect 28592 28608 28598 28620
rect 29178 28608 29184 28620
rect 28592 28580 29184 28608
rect 28592 28568 28598 28580
rect 29178 28568 29184 28580
rect 29236 28568 29242 28620
rect 29549 28611 29607 28617
rect 29549 28577 29561 28611
rect 29595 28608 29607 28611
rect 29730 28608 29736 28620
rect 29595 28580 29736 28608
rect 29595 28577 29607 28580
rect 29549 28571 29607 28577
rect 29730 28568 29736 28580
rect 29788 28568 29794 28620
rect 30009 28611 30067 28617
rect 30009 28577 30021 28611
rect 30055 28577 30067 28611
rect 30009 28571 30067 28577
rect 27065 28543 27123 28549
rect 26752 28512 27016 28540
rect 26752 28500 26758 28512
rect 25740 28444 26188 28472
rect 25740 28432 25746 28444
rect 26234 28432 26240 28484
rect 26292 28432 26298 28484
rect 26326 28432 26332 28484
rect 26384 28472 26390 28484
rect 26789 28475 26847 28481
rect 26789 28472 26801 28475
rect 26384 28444 26801 28472
rect 26384 28432 26390 28444
rect 26789 28441 26801 28444
rect 26835 28441 26847 28475
rect 26988 28472 27016 28512
rect 27065 28509 27077 28543
rect 27111 28540 27123 28543
rect 27341 28543 27399 28549
rect 27341 28540 27353 28543
rect 27111 28512 27353 28540
rect 27111 28509 27123 28512
rect 27065 28503 27123 28509
rect 27341 28509 27353 28512
rect 27387 28509 27399 28543
rect 27341 28503 27399 28509
rect 27525 28543 27583 28549
rect 27525 28509 27537 28543
rect 27571 28509 27583 28543
rect 27525 28503 27583 28509
rect 27617 28543 27675 28549
rect 27617 28509 27629 28543
rect 27663 28509 27675 28543
rect 27617 28503 27675 28509
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 27801 28543 27859 28549
rect 27801 28540 27813 28543
rect 27764 28512 27813 28540
rect 27764 28500 27770 28512
rect 27801 28509 27813 28512
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 28077 28543 28135 28549
rect 28077 28509 28089 28543
rect 28123 28540 28135 28543
rect 28353 28543 28411 28549
rect 28123 28512 28157 28540
rect 28123 28509 28135 28512
rect 28077 28503 28135 28509
rect 28353 28509 28365 28543
rect 28399 28509 28411 28543
rect 28353 28503 28411 28509
rect 28092 28472 28120 28503
rect 28258 28472 28264 28484
rect 26988 28444 28264 28472
rect 26789 28435 26847 28441
rect 28258 28432 28264 28444
rect 28316 28432 28322 28484
rect 28368 28472 28396 28503
rect 28718 28500 28724 28552
rect 28776 28500 28782 28552
rect 29086 28500 29092 28552
rect 29144 28500 29150 28552
rect 30024 28540 30052 28571
rect 32030 28568 32036 28620
rect 32088 28568 32094 28620
rect 33042 28568 33048 28620
rect 33100 28608 33106 28620
rect 33100 28580 33732 28608
rect 33100 28568 33106 28580
rect 30282 28540 30288 28552
rect 30024 28512 30288 28540
rect 30282 28500 30288 28512
rect 30340 28540 30346 28552
rect 30469 28543 30527 28549
rect 30469 28540 30481 28543
rect 30340 28512 30481 28540
rect 30340 28500 30346 28512
rect 30469 28509 30481 28512
rect 30515 28509 30527 28543
rect 30469 28503 30527 28509
rect 30837 28543 30895 28549
rect 30837 28509 30849 28543
rect 30883 28540 30895 28543
rect 31018 28540 31024 28552
rect 30883 28512 31024 28540
rect 30883 28509 30895 28512
rect 30837 28503 30895 28509
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 31113 28543 31171 28549
rect 31113 28509 31125 28543
rect 31159 28509 31171 28543
rect 31113 28503 31171 28509
rect 28534 28472 28540 28484
rect 28368 28444 28540 28472
rect 28534 28432 28540 28444
rect 28592 28472 28598 28484
rect 29104 28472 29132 28500
rect 28592 28444 29132 28472
rect 28592 28432 28598 28444
rect 30374 28432 30380 28484
rect 30432 28472 30438 28484
rect 30653 28475 30711 28481
rect 30653 28472 30665 28475
rect 30432 28444 30665 28472
rect 30432 28432 30438 28444
rect 30653 28441 30665 28444
rect 30699 28441 30711 28475
rect 30653 28435 30711 28441
rect 30742 28432 30748 28484
rect 30800 28432 30806 28484
rect 31128 28472 31156 28503
rect 31386 28500 31392 28552
rect 31444 28500 31450 28552
rect 33502 28500 33508 28552
rect 33560 28500 33566 28552
rect 33704 28549 33732 28580
rect 42812 28552 42840 28648
rect 42889 28611 42947 28617
rect 42889 28577 42901 28611
rect 42935 28608 42947 28611
rect 43257 28611 43315 28617
rect 43257 28608 43269 28611
rect 42935 28580 43269 28608
rect 42935 28577 42947 28580
rect 42889 28571 42947 28577
rect 43257 28577 43269 28580
rect 43303 28577 43315 28611
rect 43257 28571 43315 28577
rect 33689 28543 33747 28549
rect 33689 28509 33701 28543
rect 33735 28509 33747 28543
rect 33689 28503 33747 28509
rect 41874 28500 41880 28552
rect 41932 28540 41938 28552
rect 42061 28543 42119 28549
rect 42061 28540 42073 28543
rect 41932 28512 42073 28540
rect 41932 28500 41938 28512
rect 42061 28509 42073 28512
rect 42107 28509 42119 28543
rect 42061 28503 42119 28509
rect 42334 28500 42340 28552
rect 42392 28500 42398 28552
rect 42613 28543 42671 28549
rect 42613 28509 42625 28543
rect 42659 28540 42671 28543
rect 42794 28540 42800 28552
rect 42659 28512 42800 28540
rect 42659 28509 42671 28512
rect 42613 28503 42671 28509
rect 42794 28500 42800 28512
rect 42852 28500 42858 28552
rect 43073 28543 43131 28549
rect 43073 28509 43085 28543
rect 43119 28509 43131 28543
rect 43073 28503 43131 28509
rect 43165 28543 43223 28549
rect 43165 28509 43177 28543
rect 43211 28540 43223 28543
rect 43211 28512 43300 28540
rect 43211 28509 43223 28512
rect 43165 28503 43223 28509
rect 32122 28472 32128 28484
rect 31128 28444 32128 28472
rect 32122 28432 32128 28444
rect 32180 28432 32186 28484
rect 32300 28475 32358 28481
rect 32300 28441 32312 28475
rect 32346 28472 32358 28475
rect 33962 28472 33968 28484
rect 32346 28444 33968 28472
rect 32346 28441 32358 28444
rect 32300 28435 32358 28441
rect 33962 28432 33968 28444
rect 34020 28432 34026 28484
rect 36262 28432 36268 28484
rect 36320 28472 36326 28484
rect 42978 28472 42984 28484
rect 36320 28444 42984 28472
rect 36320 28432 36326 28444
rect 42978 28432 42984 28444
rect 43036 28472 43042 28484
rect 43088 28472 43116 28503
rect 43036 28444 43116 28472
rect 43036 28432 43042 28444
rect 21223 28376 21404 28404
rect 21223 28373 21235 28376
rect 21177 28367 21235 28373
rect 21910 28364 21916 28416
rect 21968 28404 21974 28416
rect 22649 28407 22707 28413
rect 22649 28404 22661 28407
rect 21968 28376 22661 28404
rect 21968 28364 21974 28376
rect 22649 28373 22661 28376
rect 22695 28373 22707 28407
rect 22649 28367 22707 28373
rect 24302 28364 24308 28416
rect 24360 28364 24366 28416
rect 25038 28364 25044 28416
rect 25096 28364 25102 28416
rect 26142 28364 26148 28416
rect 26200 28404 26206 28416
rect 26349 28404 26377 28432
rect 43272 28416 43300 28512
rect 26200 28376 26377 28404
rect 26200 28364 26206 28376
rect 26418 28364 26424 28416
rect 26476 28413 26482 28416
rect 26476 28407 26495 28413
rect 26483 28373 26495 28407
rect 26476 28367 26495 28373
rect 26476 28364 26482 28367
rect 26602 28364 26608 28416
rect 26660 28364 26666 28416
rect 27246 28364 27252 28416
rect 27304 28404 27310 28416
rect 27433 28407 27491 28413
rect 27433 28404 27445 28407
rect 27304 28376 27445 28404
rect 27304 28364 27310 28376
rect 27433 28373 27445 28376
rect 27479 28373 27491 28407
rect 27433 28367 27491 28373
rect 27522 28364 27528 28416
rect 27580 28404 27586 28416
rect 27709 28407 27767 28413
rect 27709 28404 27721 28407
rect 27580 28376 27721 28404
rect 27580 28364 27586 28376
rect 27709 28373 27721 28376
rect 27755 28373 27767 28407
rect 27709 28367 27767 28373
rect 28626 28364 28632 28416
rect 28684 28404 28690 28416
rect 29273 28407 29331 28413
rect 29273 28404 29285 28407
rect 28684 28376 29285 28404
rect 28684 28364 28690 28376
rect 29273 28373 29285 28376
rect 29319 28373 29331 28407
rect 29273 28367 29331 28373
rect 31021 28407 31079 28413
rect 31021 28373 31033 28407
rect 31067 28404 31079 28407
rect 33226 28404 33232 28416
rect 31067 28376 33232 28404
rect 31067 28373 31079 28376
rect 31021 28367 31079 28373
rect 33226 28364 33232 28376
rect 33284 28364 33290 28416
rect 33502 28364 33508 28416
rect 33560 28404 33566 28416
rect 33873 28407 33931 28413
rect 33873 28404 33885 28407
rect 33560 28376 33885 28404
rect 33560 28364 33566 28376
rect 33873 28373 33885 28376
rect 33919 28373 33931 28407
rect 33873 28367 33931 28373
rect 41874 28364 41880 28416
rect 41932 28364 41938 28416
rect 43254 28364 43260 28416
rect 43312 28364 43318 28416
rect 1104 28314 43884 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 43884 28314
rect 1104 28240 43884 28262
rect 1673 28203 1731 28209
rect 1673 28169 1685 28203
rect 1719 28200 1731 28203
rect 1762 28200 1768 28212
rect 1719 28172 1768 28200
rect 1719 28169 1731 28172
rect 1673 28163 1731 28169
rect 1762 28160 1768 28172
rect 1820 28160 1826 28212
rect 1854 28160 1860 28212
rect 1912 28160 1918 28212
rect 2406 28200 2412 28212
rect 2148 28172 2412 28200
rect 1489 28135 1547 28141
rect 1489 28101 1501 28135
rect 1535 28132 1547 28135
rect 2148 28132 2176 28172
rect 2406 28160 2412 28172
rect 2464 28200 2470 28212
rect 3786 28200 3792 28212
rect 2464 28172 3792 28200
rect 2464 28160 2470 28172
rect 3786 28160 3792 28172
rect 3844 28160 3850 28212
rect 4062 28160 4068 28212
rect 4120 28200 4126 28212
rect 4338 28200 4344 28212
rect 4120 28172 4344 28200
rect 4120 28160 4126 28172
rect 4338 28160 4344 28172
rect 4396 28160 4402 28212
rect 4706 28160 4712 28212
rect 4764 28200 4770 28212
rect 4801 28203 4859 28209
rect 4801 28200 4813 28203
rect 4764 28172 4813 28200
rect 4764 28160 4770 28172
rect 4801 28169 4813 28172
rect 4847 28169 4859 28203
rect 4801 28163 4859 28169
rect 5166 28160 5172 28212
rect 5224 28160 5230 28212
rect 5442 28160 5448 28212
rect 5500 28200 5506 28212
rect 5905 28203 5963 28209
rect 5905 28200 5917 28203
rect 5500 28172 5917 28200
rect 5500 28160 5506 28172
rect 5905 28169 5917 28172
rect 5951 28169 5963 28203
rect 5905 28163 5963 28169
rect 6730 28160 6736 28212
rect 6788 28200 6794 28212
rect 7653 28203 7711 28209
rect 7653 28200 7665 28203
rect 6788 28172 7665 28200
rect 6788 28160 6794 28172
rect 7653 28169 7665 28172
rect 7699 28200 7711 28203
rect 9122 28200 9128 28212
rect 7699 28172 9128 28200
rect 7699 28169 7711 28172
rect 7653 28163 7711 28169
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 9214 28160 9220 28212
rect 9272 28200 9278 28212
rect 10137 28203 10195 28209
rect 10137 28200 10149 28203
rect 9272 28172 10149 28200
rect 9272 28160 9278 28172
rect 10137 28169 10149 28172
rect 10183 28169 10195 28203
rect 10137 28163 10195 28169
rect 10594 28160 10600 28212
rect 10652 28160 10658 28212
rect 10778 28160 10784 28212
rect 10836 28200 10842 28212
rect 12069 28203 12127 28209
rect 12069 28200 12081 28203
rect 10836 28172 12081 28200
rect 10836 28160 10842 28172
rect 12069 28169 12081 28172
rect 12115 28169 12127 28203
rect 12069 28163 12127 28169
rect 12897 28203 12955 28209
rect 12897 28169 12909 28203
rect 12943 28200 12955 28203
rect 12986 28200 12992 28212
rect 12943 28172 12992 28200
rect 12943 28169 12955 28172
rect 12897 28163 12955 28169
rect 12986 28160 12992 28172
rect 13044 28160 13050 28212
rect 13078 28160 13084 28212
rect 13136 28160 13142 28212
rect 13170 28160 13176 28212
rect 13228 28200 13234 28212
rect 13265 28203 13323 28209
rect 13265 28200 13277 28203
rect 13228 28172 13277 28200
rect 13228 28160 13234 28172
rect 13265 28169 13277 28172
rect 13311 28169 13323 28203
rect 13265 28163 13323 28169
rect 1535 28104 2176 28132
rect 2225 28135 2283 28141
rect 1535 28101 1547 28104
rect 1489 28095 1547 28101
rect 2225 28101 2237 28135
rect 2271 28132 2283 28135
rect 3050 28132 3056 28144
rect 2271 28104 3056 28132
rect 2271 28101 2283 28104
rect 2225 28095 2283 28101
rect 3050 28092 3056 28104
rect 3108 28092 3114 28144
rect 3145 28135 3203 28141
rect 3145 28101 3157 28135
rect 3191 28132 3203 28135
rect 3234 28132 3240 28144
rect 3191 28104 3240 28132
rect 3191 28101 3203 28104
rect 3145 28095 3203 28101
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28064 1823 28067
rect 1854 28064 1860 28076
rect 1811 28036 1860 28064
rect 1811 28033 1823 28036
rect 1765 28027 1823 28033
rect 1854 28024 1860 28036
rect 1912 28024 1918 28076
rect 2317 28067 2375 28073
rect 2317 28033 2329 28067
rect 2363 28064 2375 28067
rect 3160 28064 3188 28095
rect 3234 28092 3240 28104
rect 3292 28092 3298 28144
rect 3620 28104 4476 28132
rect 2363 28036 3188 28064
rect 2363 28033 2375 28036
rect 2317 28027 2375 28033
rect 3510 28024 3516 28076
rect 3568 28024 3574 28076
rect 2130 27996 2136 28008
rect 1504 27968 2136 27996
rect 1504 27937 1532 27968
rect 2130 27956 2136 27968
rect 2188 27956 2194 28008
rect 2498 27956 2504 28008
rect 2556 27956 2562 28008
rect 3329 27999 3387 28005
rect 3329 27965 3341 27999
rect 3375 27996 3387 27999
rect 3620 27996 3648 28104
rect 4448 28073 4476 28104
rect 3697 28067 3755 28073
rect 3697 28033 3709 28067
rect 3743 28033 3755 28067
rect 3697 28027 3755 28033
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28033 4215 28067
rect 4157 28027 4215 28033
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28064 4491 28067
rect 4985 28067 5043 28073
rect 4479 28036 4752 28064
rect 4479 28033 4491 28036
rect 4433 28027 4491 28033
rect 3375 27968 3648 27996
rect 3375 27965 3387 27968
rect 3329 27959 3387 27965
rect 1489 27931 1547 27937
rect 1489 27897 1501 27931
rect 1535 27897 1547 27931
rect 3712 27928 3740 28027
rect 4172 27996 4200 28027
rect 4172 27968 4660 27996
rect 4632 27940 4660 27968
rect 3878 27928 3884 27940
rect 3712 27900 3884 27928
rect 1489 27891 1547 27897
rect 3878 27888 3884 27900
rect 3936 27928 3942 27940
rect 4522 27928 4528 27940
rect 3936 27900 4528 27928
rect 3936 27888 3942 27900
rect 4522 27888 4528 27900
rect 4580 27888 4586 27940
rect 4614 27888 4620 27940
rect 4672 27888 4678 27940
rect 4724 27928 4752 28036
rect 4985 28033 4997 28067
rect 5031 28033 5043 28067
rect 4985 28027 5043 28033
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5184 28064 5212 28160
rect 5537 28135 5595 28141
rect 5537 28132 5549 28135
rect 5276 28104 5549 28132
rect 5276 28073 5304 28104
rect 5537 28101 5549 28104
rect 5583 28101 5595 28135
rect 6086 28132 6092 28144
rect 5537 28095 5595 28101
rect 6012 28104 6092 28132
rect 5123 28036 5212 28064
rect 5261 28067 5319 28073
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 5261 28033 5273 28067
rect 5307 28033 5319 28067
rect 5261 28027 5319 28033
rect 4798 27956 4804 28008
rect 4856 27996 4862 28008
rect 5000 27996 5028 28027
rect 5350 28024 5356 28076
rect 5408 28024 5414 28076
rect 5626 28064 5632 28076
rect 5465 28063 5632 28064
rect 5449 28057 5632 28063
rect 4856 27968 5028 27996
rect 5169 27999 5227 28005
rect 4856 27956 4862 27968
rect 5169 27965 5181 27999
rect 5215 27996 5227 27999
rect 5368 27996 5396 28024
rect 5449 28023 5461 28057
rect 5495 28036 5632 28057
rect 5495 28023 5507 28036
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 6012 28073 6040 28104
rect 6086 28092 6092 28104
rect 6144 28092 6150 28144
rect 6457 28135 6515 28141
rect 6457 28132 6469 28135
rect 6380 28104 6469 28132
rect 5721 28067 5779 28073
rect 5721 28033 5733 28067
rect 5767 28033 5779 28067
rect 5721 28027 5779 28033
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 5997 28027 6055 28033
rect 5449 28017 5507 28023
rect 5215 27968 5396 27996
rect 5215 27965 5227 27968
rect 5169 27959 5227 27965
rect 5534 27956 5540 28008
rect 5592 27996 5598 28008
rect 5736 27996 5764 28027
rect 5592 27968 5764 27996
rect 6380 27996 6408 28104
rect 6457 28101 6469 28104
rect 6503 28101 6515 28135
rect 7098 28132 7104 28144
rect 6457 28095 6515 28101
rect 6886 28104 7104 28132
rect 6886 28098 6914 28104
rect 6840 28076 6914 28098
rect 7098 28092 7104 28104
rect 7156 28092 7162 28144
rect 9309 28135 9367 28141
rect 9309 28132 9321 28135
rect 8864 28104 9321 28132
rect 6638 28024 6644 28076
rect 6696 28024 6702 28076
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 6822 28024 6828 28076
rect 6880 28070 6914 28076
rect 6880 28024 6886 28070
rect 7190 28024 7196 28076
rect 7248 28064 7254 28076
rect 7469 28067 7527 28073
rect 7469 28064 7481 28067
rect 7248 28036 7481 28064
rect 7248 28024 7254 28036
rect 7469 28033 7481 28036
rect 7515 28033 7527 28067
rect 7469 28027 7527 28033
rect 7745 28067 7803 28073
rect 7745 28033 7757 28067
rect 7791 28064 7803 28067
rect 7791 28036 8064 28064
rect 7791 28033 7803 28036
rect 7745 28027 7803 28033
rect 6656 27996 6684 28024
rect 8036 28008 8064 28036
rect 8294 28024 8300 28076
rect 8352 28064 8358 28076
rect 8864 28073 8892 28104
rect 9309 28101 9321 28104
rect 9355 28132 9367 28135
rect 9677 28135 9735 28141
rect 9677 28132 9689 28135
rect 9355 28104 9689 28132
rect 9355 28101 9367 28104
rect 9309 28095 9367 28101
rect 9677 28101 9689 28104
rect 9723 28101 9735 28135
rect 9677 28095 9735 28101
rect 10502 28092 10508 28144
rect 10560 28132 10566 28144
rect 10560 28104 11192 28132
rect 10560 28092 10566 28104
rect 8573 28067 8631 28073
rect 8573 28064 8585 28067
rect 8352 28036 8585 28064
rect 8352 28024 8358 28036
rect 8573 28033 8585 28036
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28033 8907 28067
rect 8849 28027 8907 28033
rect 9217 28067 9275 28073
rect 9217 28033 9229 28067
rect 9263 28064 9275 28067
rect 9401 28067 9459 28073
rect 9263 28036 9352 28064
rect 9263 28033 9275 28036
rect 9217 28027 9275 28033
rect 9324 28008 9352 28036
rect 9401 28033 9413 28067
rect 9447 28033 9459 28067
rect 9401 28027 9459 28033
rect 9493 28067 9551 28073
rect 9493 28033 9505 28067
rect 9539 28064 9551 28067
rect 9769 28067 9827 28073
rect 9539 28036 9619 28064
rect 9539 28033 9551 28036
rect 9493 28027 9551 28033
rect 6380 27968 6597 27996
rect 6656 27968 6914 27996
rect 5592 27956 5598 27968
rect 4724 27900 5488 27928
rect 5460 27872 5488 27900
rect 6178 27888 6184 27940
rect 6236 27928 6242 27940
rect 6457 27931 6515 27937
rect 6457 27928 6469 27931
rect 6236 27900 6469 27928
rect 6236 27888 6242 27900
rect 6457 27897 6469 27900
rect 6503 27897 6515 27931
rect 6457 27891 6515 27897
rect 2682 27820 2688 27872
rect 2740 27820 2746 27872
rect 3142 27820 3148 27872
rect 3200 27860 3206 27872
rect 3513 27863 3571 27869
rect 3513 27860 3525 27863
rect 3200 27832 3525 27860
rect 3200 27820 3206 27832
rect 3513 27829 3525 27832
rect 3559 27829 3571 27863
rect 3513 27823 3571 27829
rect 3973 27863 4031 27869
rect 3973 27829 3985 27863
rect 4019 27860 4031 27863
rect 5258 27860 5264 27872
rect 4019 27832 5264 27860
rect 4019 27829 4031 27832
rect 3973 27823 4031 27829
rect 5258 27820 5264 27832
rect 5316 27820 5322 27872
rect 5442 27820 5448 27872
rect 5500 27820 5506 27872
rect 6569 27860 6597 27968
rect 6886 27928 6914 27968
rect 8018 27956 8024 28008
rect 8076 27956 8082 28008
rect 9306 27956 9312 28008
rect 9364 27956 9370 28008
rect 9416 27996 9444 28027
rect 9416 27968 9536 27996
rect 9508 27940 9536 27968
rect 8202 27928 8208 27940
rect 6886 27900 8208 27928
rect 8202 27888 8208 27900
rect 8260 27928 8266 27940
rect 8260 27900 8892 27928
rect 8260 27888 8266 27900
rect 6822 27860 6828 27872
rect 6569 27832 6828 27860
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 7285 27863 7343 27869
rect 7285 27829 7297 27863
rect 7331 27860 7343 27863
rect 7558 27860 7564 27872
rect 7331 27832 7564 27860
rect 7331 27829 7343 27832
rect 7285 27823 7343 27829
rect 7558 27820 7564 27832
rect 7616 27820 7622 27872
rect 7926 27820 7932 27872
rect 7984 27860 7990 27872
rect 8389 27863 8447 27869
rect 8389 27860 8401 27863
rect 7984 27832 8401 27860
rect 7984 27820 7990 27832
rect 8389 27829 8401 27832
rect 8435 27829 8447 27863
rect 8389 27823 8447 27829
rect 8754 27820 8760 27872
rect 8812 27820 8818 27872
rect 8864 27860 8892 27900
rect 8938 27888 8944 27940
rect 8996 27928 9002 27940
rect 9490 27928 9496 27940
rect 8996 27900 9496 27928
rect 8996 27888 9002 27900
rect 9490 27888 9496 27900
rect 9548 27888 9554 27940
rect 9591 27860 9619 28036
rect 9769 28033 9781 28067
rect 9815 28033 9827 28067
rect 9769 28027 9827 28033
rect 9784 27996 9812 28027
rect 9858 28024 9864 28076
rect 9916 28024 9922 28076
rect 10965 28067 11023 28073
rect 10965 28064 10977 28067
rect 10796 28036 10977 28064
rect 10318 27996 10324 28008
rect 9784 27968 10324 27996
rect 10318 27956 10324 27968
rect 10376 27956 10382 28008
rect 10410 27956 10416 28008
rect 10468 27996 10474 28008
rect 10796 28005 10824 28036
rect 10965 28033 10977 28036
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 10781 27999 10839 28005
rect 10781 27996 10793 27999
rect 10468 27968 10793 27996
rect 10468 27956 10474 27968
rect 10781 27965 10793 27968
rect 10827 27965 10839 27999
rect 10781 27959 10839 27965
rect 11054 27956 11060 28008
rect 11112 27956 11118 28008
rect 11164 27996 11192 28104
rect 11238 28092 11244 28144
rect 11296 28132 11302 28144
rect 11882 28132 11888 28144
rect 11296 28104 11888 28132
rect 11296 28092 11302 28104
rect 11330 28024 11336 28076
rect 11388 28064 11394 28076
rect 11716 28073 11744 28104
rect 11882 28092 11888 28104
rect 11940 28092 11946 28144
rect 12437 28135 12495 28141
rect 12437 28101 12449 28135
rect 12483 28132 12495 28135
rect 13096 28132 13124 28160
rect 12483 28104 13124 28132
rect 13280 28132 13308 28163
rect 13354 28160 13360 28212
rect 13412 28200 13418 28212
rect 13814 28200 13820 28212
rect 13412 28172 13820 28200
rect 13412 28160 13418 28172
rect 13814 28160 13820 28172
rect 13872 28160 13878 28212
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 15010 28200 15016 28212
rect 14240 28172 15016 28200
rect 14240 28160 14246 28172
rect 15010 28160 15016 28172
rect 15068 28160 15074 28212
rect 15378 28160 15384 28212
rect 15436 28200 15442 28212
rect 15473 28203 15531 28209
rect 15473 28200 15485 28203
rect 15436 28172 15485 28200
rect 15436 28160 15442 28172
rect 15473 28169 15485 28172
rect 15519 28200 15531 28203
rect 15930 28200 15936 28212
rect 15519 28172 15936 28200
rect 15519 28169 15531 28172
rect 15473 28163 15531 28169
rect 15930 28160 15936 28172
rect 15988 28160 15994 28212
rect 16758 28160 16764 28212
rect 16816 28200 16822 28212
rect 16816 28172 20668 28200
rect 16816 28160 16822 28172
rect 13280 28104 13676 28132
rect 12483 28101 12495 28104
rect 12437 28095 12495 28101
rect 11517 28067 11575 28073
rect 11517 28064 11529 28067
rect 11388 28036 11529 28064
rect 11388 28024 11394 28036
rect 11517 28033 11529 28036
rect 11563 28033 11575 28067
rect 11517 28027 11575 28033
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 13078 28024 13084 28076
rect 13136 28073 13142 28076
rect 13136 28067 13158 28073
rect 13146 28033 13158 28067
rect 13136 28027 13158 28033
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 13136 28024 13142 28027
rect 12066 27996 12072 28008
rect 11164 27968 12072 27996
rect 12066 27956 12072 27968
rect 12124 27996 12130 28008
rect 12529 27999 12587 28005
rect 12529 27996 12541 27999
rect 12124 27968 12541 27996
rect 12124 27956 12130 27968
rect 12529 27965 12541 27968
rect 12575 27965 12587 27999
rect 12529 27959 12587 27965
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27996 12771 27999
rect 12986 27996 12992 28008
rect 12759 27968 12992 27996
rect 12759 27965 12771 27968
rect 12713 27959 12771 27965
rect 12986 27956 12992 27968
rect 13044 27956 13050 28008
rect 13372 27996 13400 28027
rect 13538 28024 13544 28076
rect 13596 28024 13602 28076
rect 13648 28073 13676 28104
rect 13722 28092 13728 28144
rect 13780 28132 13786 28144
rect 14645 28135 14703 28141
rect 14645 28132 14657 28135
rect 13780 28104 14657 28132
rect 13780 28092 13786 28104
rect 14645 28101 14657 28104
rect 14691 28101 14703 28135
rect 14645 28095 14703 28101
rect 15286 28092 15292 28144
rect 15344 28132 15350 28144
rect 16390 28132 16396 28144
rect 15344 28104 16396 28132
rect 15344 28092 15350 28104
rect 16390 28092 16396 28104
rect 16448 28132 16454 28144
rect 16448 28104 16896 28132
rect 16448 28092 16454 28104
rect 13633 28067 13691 28073
rect 13633 28033 13645 28067
rect 13679 28033 13691 28067
rect 13633 28027 13691 28033
rect 13814 28024 13820 28076
rect 13872 28024 13878 28076
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28064 14611 28067
rect 14737 28067 14795 28073
rect 14599 28036 14688 28064
rect 14599 28033 14611 28036
rect 14553 28027 14611 28033
rect 14660 28008 14688 28036
rect 14737 28033 14749 28067
rect 14783 28064 14795 28067
rect 16482 28064 16488 28076
rect 14783 28036 16488 28064
rect 14783 28033 14795 28036
rect 14737 28027 14795 28033
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 14182 27996 14188 28008
rect 13372 27968 14188 27996
rect 9674 27888 9680 27940
rect 9732 27928 9738 27940
rect 10045 27931 10103 27937
rect 10045 27928 10057 27931
rect 9732 27900 10057 27928
rect 9732 27888 9738 27900
rect 10045 27897 10057 27900
rect 10091 27897 10103 27931
rect 10045 27891 10103 27897
rect 10226 27888 10232 27940
rect 10284 27928 10290 27940
rect 11606 27928 11612 27940
rect 10284 27900 11612 27928
rect 10284 27888 10290 27900
rect 11606 27888 11612 27900
rect 11664 27888 11670 27940
rect 12342 27928 12348 27940
rect 11716 27900 12348 27928
rect 11716 27860 11744 27900
rect 12342 27888 12348 27900
rect 12400 27888 12406 27940
rect 12434 27888 12440 27940
rect 12492 27928 12498 27940
rect 13372 27928 13400 27968
rect 13648 27940 13676 27968
rect 14182 27956 14188 27968
rect 14240 27956 14246 28008
rect 14642 27956 14648 28008
rect 14700 27956 14706 28008
rect 15562 27956 15568 28008
rect 15620 27956 15626 28008
rect 16669 27999 16727 28005
rect 16669 27965 16681 27999
rect 16715 27996 16727 27999
rect 16758 27996 16764 28008
rect 16715 27968 16764 27996
rect 16715 27965 16727 27968
rect 16669 27959 16727 27965
rect 16758 27956 16764 27968
rect 16816 27956 16822 28008
rect 16868 28005 16896 28104
rect 18414 28092 18420 28144
rect 18472 28092 18478 28144
rect 18969 28135 19027 28141
rect 18969 28101 18981 28135
rect 19015 28132 19027 28135
rect 19521 28135 19579 28141
rect 19521 28132 19533 28135
rect 19015 28104 19533 28132
rect 19015 28101 19027 28104
rect 18969 28095 19027 28101
rect 19521 28101 19533 28104
rect 19567 28101 19579 28135
rect 19521 28095 19579 28101
rect 17586 28024 17592 28076
rect 17644 28024 17650 28076
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28033 17923 28067
rect 18432 28064 18460 28092
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18432 28036 19073 28064
rect 17865 28027 17923 28033
rect 19061 28033 19073 28036
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 16853 27999 16911 28005
rect 16853 27965 16865 27999
rect 16899 27965 16911 27999
rect 16853 27959 16911 27965
rect 17678 27956 17684 28008
rect 17736 28005 17742 28008
rect 17736 27999 17785 28005
rect 17736 27965 17739 27999
rect 17773 27965 17785 27999
rect 17880 27996 17908 28027
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19720 28073 19748 28172
rect 19794 28092 19800 28144
rect 19852 28132 19858 28144
rect 20640 28132 20668 28172
rect 24302 28160 24308 28212
rect 24360 28160 24366 28212
rect 24394 28160 24400 28212
rect 24452 28200 24458 28212
rect 24581 28203 24639 28209
rect 24581 28200 24593 28203
rect 24452 28172 24593 28200
rect 24452 28160 24458 28172
rect 24581 28169 24593 28172
rect 24627 28169 24639 28203
rect 24581 28163 24639 28169
rect 26234 28160 26240 28212
rect 26292 28200 26298 28212
rect 27706 28200 27712 28212
rect 26292 28172 27712 28200
rect 26292 28160 26298 28172
rect 27706 28160 27712 28172
rect 27764 28160 27770 28212
rect 28629 28203 28687 28209
rect 28629 28169 28641 28203
rect 28675 28200 28687 28203
rect 28675 28172 28856 28200
rect 28675 28169 28687 28172
rect 28629 28163 28687 28169
rect 20898 28132 20904 28144
rect 19852 28104 20567 28132
rect 20640 28104 20904 28132
rect 19852 28092 19858 28104
rect 19429 28067 19487 28073
rect 19429 28064 19441 28067
rect 19392 28036 19441 28064
rect 19392 28024 19398 28036
rect 19429 28033 19441 28036
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 19972 28067 20030 28073
rect 19972 28033 19984 28067
rect 20018 28064 20030 28067
rect 20438 28064 20444 28076
rect 20018 28036 20444 28064
rect 20018 28033 20030 28036
rect 19972 28027 20030 28033
rect 20438 28024 20444 28036
rect 20496 28024 20502 28076
rect 20539 28064 20567 28104
rect 20898 28092 20904 28104
rect 20956 28092 20962 28144
rect 27798 28132 27804 28144
rect 22480 28104 27804 28132
rect 22480 28076 22508 28104
rect 20539 28036 20760 28064
rect 17880 27968 18267 27996
rect 17736 27959 17785 27965
rect 17736 27956 17742 27959
rect 12492 27900 13400 27928
rect 12492 27888 12498 27900
rect 13630 27888 13636 27940
rect 13688 27888 13694 27940
rect 15194 27928 15200 27940
rect 14384 27900 15200 27928
rect 14384 27872 14412 27900
rect 15194 27888 15200 27900
rect 15252 27888 15258 27940
rect 16132 27900 16335 27928
rect 8864 27832 11744 27860
rect 12158 27820 12164 27872
rect 12216 27860 12222 27872
rect 13538 27860 13544 27872
rect 12216 27832 13544 27860
rect 12216 27820 12222 27832
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 14366 27820 14372 27872
rect 14424 27820 14430 27872
rect 15010 27820 15016 27872
rect 15068 27860 15074 27872
rect 16132 27860 16160 27900
rect 15068 27832 16160 27860
rect 15068 27820 15074 27832
rect 16206 27820 16212 27872
rect 16264 27820 16270 27872
rect 16307 27860 16335 27900
rect 17034 27888 17040 27940
rect 17092 27928 17098 27940
rect 17313 27931 17371 27937
rect 17313 27928 17325 27931
rect 17092 27900 17325 27928
rect 17092 27888 17098 27900
rect 17313 27897 17325 27900
rect 17359 27897 17371 27931
rect 17313 27891 17371 27897
rect 17586 27860 17592 27872
rect 16307 27832 17592 27860
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 17770 27820 17776 27872
rect 17828 27860 17834 27872
rect 18239 27860 18267 27968
rect 18966 27956 18972 28008
rect 19024 27996 19030 28008
rect 19153 27999 19211 28005
rect 19153 27996 19165 27999
rect 19024 27968 19165 27996
rect 19024 27956 19030 27968
rect 19153 27965 19165 27968
rect 19199 27965 19211 27999
rect 20732 27996 20760 28036
rect 21910 28024 21916 28076
rect 21968 28024 21974 28076
rect 22462 28024 22468 28076
rect 22520 28024 22526 28076
rect 22557 28067 22615 28073
rect 22557 28033 22569 28067
rect 22603 28064 22615 28067
rect 22646 28064 22652 28076
rect 22603 28036 22652 28064
rect 22603 28033 22615 28036
rect 22557 28027 22615 28033
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 22940 28073 22968 28104
rect 27798 28092 27804 28104
rect 27856 28132 27862 28144
rect 28828 28132 28856 28172
rect 30742 28160 30748 28212
rect 30800 28200 30806 28212
rect 31941 28203 31999 28209
rect 31941 28200 31953 28203
rect 30800 28172 31953 28200
rect 30800 28160 30806 28172
rect 31941 28169 31953 28172
rect 31987 28169 31999 28203
rect 31941 28163 31999 28169
rect 32122 28160 32128 28212
rect 32180 28200 32186 28212
rect 33505 28203 33563 28209
rect 33505 28200 33517 28203
rect 32180 28172 33517 28200
rect 32180 28160 32186 28172
rect 33505 28169 33517 28172
rect 33551 28169 33563 28203
rect 33505 28163 33563 28169
rect 33962 28160 33968 28212
rect 34020 28160 34026 28212
rect 41874 28200 41880 28212
rect 41386 28172 41880 28200
rect 28966 28135 29024 28141
rect 28966 28132 28978 28135
rect 27856 28104 28764 28132
rect 28828 28104 28978 28132
rect 27856 28092 27862 28104
rect 22925 28067 22983 28073
rect 22925 28033 22937 28067
rect 22971 28033 22983 28067
rect 22925 28027 22983 28033
rect 23192 28067 23250 28073
rect 23192 28033 23204 28067
rect 23238 28064 23250 28067
rect 25038 28064 25044 28076
rect 23238 28036 25044 28064
rect 23238 28033 23250 28036
rect 23192 28027 23250 28033
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25866 28024 25872 28076
rect 25924 28064 25930 28076
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 25924 28036 26065 28064
rect 25924 28024 25930 28036
rect 26053 28033 26065 28036
rect 26099 28033 26111 28067
rect 26053 28027 26111 28033
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 26786 28064 26792 28076
rect 26283 28036 26792 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 26786 28024 26792 28036
rect 26844 28024 26850 28076
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28064 27215 28067
rect 27246 28064 27252 28076
rect 27203 28036 27252 28064
rect 27203 28033 27215 28036
rect 27157 28027 27215 28033
rect 27246 28024 27252 28036
rect 27304 28024 27310 28076
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 27522 28064 27528 28076
rect 27387 28036 27528 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27522 28024 27528 28036
rect 27580 28024 27586 28076
rect 27614 28024 27620 28076
rect 27672 28024 27678 28076
rect 27706 28024 27712 28076
rect 27764 28024 27770 28076
rect 27893 28067 27951 28073
rect 27893 28033 27905 28067
rect 27939 28064 27951 28067
rect 28074 28064 28080 28076
rect 27939 28036 28080 28064
rect 27939 28033 27951 28036
rect 27893 28027 27951 28033
rect 28074 28024 28080 28036
rect 28132 28024 28138 28076
rect 28445 28067 28503 28073
rect 28445 28033 28457 28067
rect 28491 28064 28503 28067
rect 28626 28064 28632 28076
rect 28491 28036 28632 28064
rect 28491 28033 28503 28036
rect 28445 28027 28503 28033
rect 28626 28024 28632 28036
rect 28684 28024 28690 28076
rect 28736 28073 28764 28104
rect 28966 28101 28978 28104
rect 29012 28101 29024 28135
rect 28966 28095 29024 28101
rect 29270 28092 29276 28144
rect 29328 28132 29334 28144
rect 29328 28104 31754 28132
rect 29328 28092 29334 28104
rect 28721 28067 28779 28073
rect 28721 28033 28733 28067
rect 28767 28033 28779 28067
rect 30650 28064 30656 28076
rect 28721 28027 28779 28033
rect 28828 28036 30656 28064
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 20732 27968 22784 27996
rect 19153 27959 19211 27965
rect 18509 27931 18567 27937
rect 18509 27897 18521 27931
rect 18555 27928 18567 27931
rect 21361 27931 21419 27937
rect 21361 27928 21373 27931
rect 18555 27900 19748 27928
rect 18555 27897 18567 27900
rect 18509 27891 18567 27897
rect 17828 27832 18267 27860
rect 17828 27820 17834 27832
rect 18414 27820 18420 27872
rect 18472 27860 18478 27872
rect 18601 27863 18659 27869
rect 18601 27860 18613 27863
rect 18472 27832 18613 27860
rect 18472 27820 18478 27832
rect 18601 27829 18613 27832
rect 18647 27829 18659 27863
rect 19720 27860 19748 27900
rect 20824 27900 21373 27928
rect 20824 27872 20852 27900
rect 21361 27897 21373 27900
rect 21407 27897 21419 27931
rect 21361 27891 21419 27897
rect 20714 27860 20720 27872
rect 19720 27832 20720 27860
rect 18601 27823 18659 27829
rect 20714 27820 20720 27832
rect 20772 27820 20778 27872
rect 20806 27820 20812 27872
rect 20864 27820 20870 27872
rect 21082 27820 21088 27872
rect 21140 27820 21146 27872
rect 21266 27820 21272 27872
rect 21324 27860 21330 27872
rect 22756 27869 22784 27968
rect 26252 27968 27445 27996
rect 26252 27940 26280 27968
rect 27433 27965 27445 27968
rect 27479 27996 27491 27999
rect 28261 27999 28319 28005
rect 27479 27968 28120 27996
rect 27479 27965 27491 27968
rect 27433 27959 27491 27965
rect 26234 27888 26240 27940
rect 26292 27888 26298 27940
rect 27249 27931 27307 27937
rect 27249 27897 27261 27931
rect 27295 27897 27307 27931
rect 27249 27891 27307 27897
rect 22465 27863 22523 27869
rect 22465 27860 22477 27863
rect 21324 27832 22477 27860
rect 21324 27820 21330 27832
rect 22465 27829 22477 27832
rect 22511 27829 22523 27863
rect 22465 27823 22523 27829
rect 22741 27863 22799 27869
rect 22741 27829 22753 27863
rect 22787 27860 22799 27863
rect 23658 27860 23664 27872
rect 22787 27832 23664 27860
rect 22787 27829 22799 27832
rect 22741 27823 22799 27829
rect 23658 27820 23664 27832
rect 23716 27820 23722 27872
rect 25682 27820 25688 27872
rect 25740 27860 25746 27872
rect 26326 27860 26332 27872
rect 25740 27832 26332 27860
rect 25740 27820 25746 27832
rect 26326 27820 26332 27832
rect 26384 27860 26390 27872
rect 26421 27863 26479 27869
rect 26421 27860 26433 27863
rect 26384 27832 26433 27860
rect 26384 27820 26390 27832
rect 26421 27829 26433 27832
rect 26467 27829 26479 27863
rect 26421 27823 26479 27829
rect 26694 27820 26700 27872
rect 26752 27860 26758 27872
rect 26973 27863 27031 27869
rect 26973 27860 26985 27863
rect 26752 27832 26985 27860
rect 26752 27820 26758 27832
rect 26973 27829 26985 27832
rect 27019 27829 27031 27863
rect 26973 27823 27031 27829
rect 27062 27820 27068 27872
rect 27120 27860 27126 27872
rect 27264 27860 27292 27891
rect 27338 27888 27344 27940
rect 27396 27928 27402 27940
rect 27522 27928 27528 27940
rect 27396 27900 27528 27928
rect 27396 27888 27402 27900
rect 27522 27888 27528 27900
rect 27580 27888 27586 27940
rect 28092 27937 28120 27968
rect 28261 27965 28273 27999
rect 28307 27996 28319 27999
rect 28828 27996 28856 28036
rect 30650 28024 30656 28036
rect 30708 28024 30714 28076
rect 30285 27999 30343 28005
rect 30285 27996 30297 27999
rect 28307 27968 28856 27996
rect 30116 27968 30297 27996
rect 28307 27965 28319 27968
rect 28261 27959 28319 27965
rect 28077 27931 28135 27937
rect 28077 27897 28089 27931
rect 28123 27928 28135 27931
rect 28350 27928 28356 27940
rect 28123 27900 28356 27928
rect 28123 27897 28135 27900
rect 28077 27891 28135 27897
rect 28350 27888 28356 27900
rect 28408 27888 28414 27940
rect 28534 27888 28540 27940
rect 28592 27888 28598 27940
rect 28552 27860 28580 27888
rect 30116 27872 30144 27968
rect 30285 27965 30297 27968
rect 30331 27965 30343 27999
rect 30285 27959 30343 27965
rect 30374 27956 30380 28008
rect 30432 27996 30438 28008
rect 31297 27999 31355 28005
rect 31297 27996 31309 27999
rect 30432 27968 31309 27996
rect 30432 27956 30438 27968
rect 31297 27965 31309 27968
rect 31343 27965 31355 27999
rect 31297 27959 31355 27965
rect 27120 27832 28580 27860
rect 27120 27820 27126 27832
rect 30098 27820 30104 27872
rect 30156 27820 30162 27872
rect 30190 27820 30196 27872
rect 30248 27860 30254 27872
rect 30929 27863 30987 27869
rect 30929 27860 30941 27863
rect 30248 27832 30941 27860
rect 30248 27820 30254 27832
rect 30929 27829 30941 27832
rect 30975 27829 30987 27863
rect 31726 27860 31754 28104
rect 32140 28104 36308 28132
rect 32140 28076 32168 28104
rect 36280 28076 36308 28104
rect 32122 28024 32128 28076
rect 32180 28024 32186 28076
rect 32392 28067 32450 28073
rect 32392 28033 32404 28067
rect 32438 28064 32450 28067
rect 33502 28064 33508 28076
rect 32438 28036 33508 28064
rect 32438 28033 32450 28036
rect 32392 28027 32450 28033
rect 33502 28024 33508 28036
rect 33560 28024 33566 28076
rect 33594 28024 33600 28076
rect 33652 28024 33658 28076
rect 33686 28024 33692 28076
rect 33744 28064 33750 28076
rect 33781 28067 33839 28073
rect 33781 28064 33793 28067
rect 33744 28036 33793 28064
rect 33744 28024 33750 28036
rect 33781 28033 33793 28036
rect 33827 28033 33839 28067
rect 33781 28027 33839 28033
rect 36262 28024 36268 28076
rect 36320 28024 36326 28076
rect 41386 27860 41414 28172
rect 41874 28160 41880 28172
rect 41932 28160 41938 28212
rect 42334 28160 42340 28212
rect 42392 28200 42398 28212
rect 42392 28172 43300 28200
rect 42392 28160 42398 28172
rect 42613 28135 42671 28141
rect 42613 28101 42625 28135
rect 42659 28132 42671 28135
rect 42794 28132 42800 28144
rect 42659 28104 42800 28132
rect 42659 28101 42671 28104
rect 42613 28095 42671 28101
rect 42794 28092 42800 28104
rect 42852 28092 42858 28144
rect 42978 28092 42984 28144
rect 43036 28141 43042 28144
rect 43036 28132 43048 28141
rect 43036 28104 43081 28132
rect 43036 28095 43048 28104
rect 43036 28092 43042 28095
rect 43272 28073 43300 28172
rect 43257 28067 43315 28073
rect 43257 28033 43269 28067
rect 43303 28033 43315 28067
rect 43257 28027 43315 28033
rect 43349 28067 43407 28073
rect 43349 28033 43361 28067
rect 43395 28064 43407 28067
rect 43806 28064 43812 28076
rect 43395 28036 43812 28064
rect 43395 28033 43407 28036
rect 43349 28027 43407 28033
rect 43806 28024 43812 28036
rect 43864 28024 43870 28076
rect 31726 27832 41414 27860
rect 42981 27863 43039 27869
rect 30929 27823 30987 27829
rect 42981 27829 42993 27863
rect 43027 27860 43039 27863
rect 43254 27860 43260 27872
rect 43027 27832 43260 27860
rect 43027 27829 43039 27832
rect 42981 27823 43039 27829
rect 43254 27820 43260 27832
rect 43312 27860 43318 27872
rect 43533 27863 43591 27869
rect 43533 27860 43545 27863
rect 43312 27832 43545 27860
rect 43312 27820 43318 27832
rect 43533 27829 43545 27832
rect 43579 27829 43591 27863
rect 43533 27823 43591 27829
rect 1104 27770 43884 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 43884 27770
rect 1104 27696 43884 27718
rect 3605 27659 3663 27665
rect 3605 27625 3617 27659
rect 3651 27656 3663 27659
rect 3786 27656 3792 27668
rect 3651 27628 3792 27656
rect 3651 27625 3663 27628
rect 3605 27619 3663 27625
rect 3786 27616 3792 27628
rect 3844 27616 3850 27668
rect 4154 27616 4160 27668
rect 4212 27656 4218 27668
rect 4709 27659 4767 27665
rect 4709 27656 4721 27659
rect 4212 27628 4721 27656
rect 4212 27616 4218 27628
rect 4709 27625 4721 27628
rect 4755 27625 4767 27659
rect 5074 27656 5080 27668
rect 4709 27619 4767 27625
rect 4913 27628 5080 27656
rect 2038 27548 2044 27600
rect 2096 27588 2102 27600
rect 3326 27588 3332 27600
rect 2096 27560 3332 27588
rect 2096 27548 2102 27560
rect 3326 27548 3332 27560
rect 3384 27548 3390 27600
rect 3973 27591 4031 27597
rect 3973 27557 3985 27591
rect 4019 27557 4031 27591
rect 4913 27588 4941 27628
rect 5074 27616 5080 27628
rect 5132 27616 5138 27668
rect 5368 27628 5580 27656
rect 5368 27600 5396 27628
rect 3973 27551 4031 27557
rect 4356 27560 4941 27588
rect 4992 27560 5301 27588
rect 1210 27480 1216 27532
rect 1268 27520 1274 27532
rect 1857 27523 1915 27529
rect 1857 27520 1869 27523
rect 1268 27492 1869 27520
rect 1268 27480 1274 27492
rect 1857 27489 1869 27492
rect 1903 27489 1915 27523
rect 3988 27520 4016 27551
rect 4356 27532 4384 27560
rect 1857 27483 1915 27489
rect 3252 27492 4016 27520
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27421 1639 27455
rect 1581 27415 1639 27421
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27452 3111 27455
rect 3142 27452 3148 27464
rect 3099 27424 3148 27452
rect 3099 27421 3111 27424
rect 3053 27415 3111 27421
rect 1596 27328 1624 27415
rect 3142 27412 3148 27424
rect 3200 27412 3206 27464
rect 3252 27461 3280 27492
rect 4338 27480 4344 27532
rect 4396 27480 4402 27532
rect 4992 27520 5020 27560
rect 4540 27492 5020 27520
rect 5273 27520 5301 27560
rect 5350 27548 5356 27600
rect 5408 27548 5414 27600
rect 5445 27591 5503 27597
rect 5445 27557 5457 27591
rect 5491 27557 5503 27591
rect 5445 27551 5503 27557
rect 5460 27520 5488 27551
rect 5273 27492 5488 27520
rect 5552 27520 5580 27628
rect 5626 27616 5632 27668
rect 5684 27656 5690 27668
rect 5684 27628 7053 27656
rect 5684 27616 5690 27628
rect 6178 27548 6184 27600
rect 6236 27588 6242 27600
rect 6362 27588 6368 27600
rect 6236 27560 6368 27588
rect 6236 27548 6242 27560
rect 6362 27548 6368 27560
rect 6420 27548 6426 27600
rect 6733 27591 6791 27597
rect 6733 27557 6745 27591
rect 6779 27557 6791 27591
rect 7025 27588 7053 27628
rect 7098 27616 7104 27668
rect 7156 27616 7162 27668
rect 8294 27656 8300 27668
rect 7760 27628 8300 27656
rect 7760 27588 7788 27628
rect 8294 27616 8300 27628
rect 8352 27616 8358 27668
rect 8573 27659 8631 27665
rect 8573 27625 8585 27659
rect 8619 27656 8631 27659
rect 8754 27656 8760 27668
rect 8619 27628 8760 27656
rect 8619 27625 8631 27628
rect 8573 27619 8631 27625
rect 8754 27616 8760 27628
rect 8812 27616 8818 27668
rect 9769 27659 9827 27665
rect 9769 27625 9781 27659
rect 9815 27656 9827 27659
rect 9858 27656 9864 27668
rect 9815 27628 9864 27656
rect 9815 27625 9827 27628
rect 9769 27619 9827 27625
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 10318 27616 10324 27668
rect 10376 27616 10382 27668
rect 11146 27616 11152 27668
rect 11204 27656 11210 27668
rect 11241 27659 11299 27665
rect 11241 27656 11253 27659
rect 11204 27628 11253 27656
rect 11204 27616 11210 27628
rect 11241 27625 11253 27628
rect 11287 27625 11299 27659
rect 11241 27619 11299 27625
rect 11609 27659 11667 27665
rect 11609 27625 11621 27659
rect 11655 27656 11667 27659
rect 11790 27656 11796 27668
rect 11655 27628 11796 27656
rect 11655 27625 11667 27628
rect 11609 27619 11667 27625
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 12342 27616 12348 27668
rect 12400 27656 12406 27668
rect 13170 27656 13176 27668
rect 12400 27628 13176 27656
rect 12400 27616 12406 27628
rect 13170 27616 13176 27628
rect 13228 27656 13234 27668
rect 13817 27659 13875 27665
rect 13817 27656 13829 27659
rect 13228 27628 13829 27656
rect 13228 27616 13234 27628
rect 13817 27625 13829 27628
rect 13863 27625 13875 27659
rect 13817 27619 13875 27625
rect 16577 27659 16635 27665
rect 16577 27625 16589 27659
rect 16623 27656 16635 27659
rect 16942 27656 16948 27668
rect 16623 27628 16948 27656
rect 16623 27625 16635 27628
rect 16577 27619 16635 27625
rect 16942 27616 16948 27628
rect 17000 27616 17006 27668
rect 17129 27659 17187 27665
rect 17129 27625 17141 27659
rect 17175 27656 17187 27659
rect 17954 27656 17960 27668
rect 17175 27628 17960 27656
rect 17175 27625 17187 27628
rect 17129 27619 17187 27625
rect 17954 27616 17960 27628
rect 18012 27656 18018 27668
rect 18966 27656 18972 27668
rect 18012 27628 18972 27656
rect 18012 27616 18018 27628
rect 18966 27616 18972 27628
rect 19024 27616 19030 27668
rect 19334 27616 19340 27668
rect 19392 27656 19398 27668
rect 20070 27656 20076 27668
rect 19392 27628 20076 27656
rect 19392 27616 19398 27628
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 20346 27616 20352 27668
rect 20404 27656 20410 27668
rect 21726 27656 21732 27668
rect 20404 27628 21732 27656
rect 20404 27616 20410 27628
rect 21726 27616 21732 27628
rect 21784 27616 21790 27668
rect 25155 27628 27292 27656
rect 7025 27560 7788 27588
rect 6733 27551 6791 27557
rect 6748 27520 6776 27551
rect 5552 27492 5764 27520
rect 6748 27492 7420 27520
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 3421 27455 3479 27461
rect 3421 27421 3433 27455
rect 3467 27452 3479 27455
rect 3694 27452 3700 27464
rect 3467 27424 3700 27452
rect 3467 27421 3479 27424
rect 3421 27415 3479 27421
rect 3694 27412 3700 27424
rect 3752 27412 3758 27464
rect 3878 27412 3884 27464
rect 3936 27412 3942 27464
rect 4540 27461 4568 27492
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27421 4215 27455
rect 4157 27415 4215 27421
rect 4249 27455 4307 27461
rect 4249 27421 4261 27455
rect 4295 27452 4307 27455
rect 4525 27455 4583 27461
rect 4295 27424 4476 27452
rect 4295 27421 4307 27424
rect 4249 27415 4307 27421
rect 3329 27387 3387 27393
rect 3329 27353 3341 27387
rect 3375 27384 3387 27387
rect 3896 27384 3924 27412
rect 3375 27356 3924 27384
rect 4172 27384 4200 27415
rect 4448 27396 4476 27424
rect 4525 27421 4537 27455
rect 4571 27421 4583 27455
rect 4525 27415 4583 27421
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27452 4675 27455
rect 4706 27452 4712 27464
rect 4663 27424 4712 27452
rect 4663 27421 4675 27424
rect 4617 27415 4675 27421
rect 4706 27412 4712 27424
rect 4764 27412 4770 27464
rect 4982 27412 4988 27464
rect 5040 27412 5046 27464
rect 5077 27455 5135 27461
rect 5077 27421 5089 27455
rect 5123 27421 5135 27455
rect 5077 27415 5135 27421
rect 5169 27455 5227 27461
rect 5169 27421 5181 27455
rect 5215 27452 5227 27455
rect 5258 27452 5264 27464
rect 5215 27424 5264 27452
rect 5215 27421 5227 27424
rect 5169 27415 5227 27421
rect 4172 27356 4292 27384
rect 3375 27353 3387 27356
rect 3329 27347 3387 27353
rect 4264 27328 4292 27356
rect 4338 27344 4344 27396
rect 4396 27344 4402 27396
rect 4430 27344 4436 27396
rect 4488 27384 4494 27396
rect 4488 27356 4752 27384
rect 4488 27344 4494 27356
rect 1578 27276 1584 27328
rect 1636 27276 1642 27328
rect 2498 27276 2504 27328
rect 2556 27316 2562 27328
rect 4246 27316 4252 27328
rect 2556 27288 4252 27316
rect 2556 27276 2562 27288
rect 4246 27276 4252 27288
rect 4304 27276 4310 27328
rect 4724 27316 4752 27356
rect 4798 27344 4804 27396
rect 4856 27384 4862 27396
rect 5092 27384 5120 27415
rect 5258 27412 5264 27424
rect 5316 27412 5322 27464
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5626 27452 5632 27464
rect 5399 27424 5632 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5626 27412 5632 27424
rect 5684 27412 5690 27464
rect 5736 27461 5764 27492
rect 5721 27455 5779 27461
rect 5721 27421 5733 27455
rect 5767 27421 5779 27455
rect 5721 27415 5779 27421
rect 6733 27455 6791 27461
rect 6733 27421 6745 27455
rect 6779 27421 6791 27455
rect 6733 27415 6791 27421
rect 7009 27455 7067 27461
rect 7009 27421 7021 27455
rect 7055 27452 7067 27455
rect 7282 27452 7288 27464
rect 7055 27424 7288 27452
rect 7055 27421 7067 27424
rect 7009 27415 7067 27421
rect 4856 27356 5120 27384
rect 5445 27387 5503 27393
rect 4856 27344 4862 27356
rect 5445 27353 5457 27387
rect 5491 27384 5503 27387
rect 5534 27384 5540 27396
rect 5491 27356 5540 27384
rect 5491 27353 5503 27356
rect 5445 27347 5503 27353
rect 5534 27344 5540 27356
rect 5592 27384 5598 27396
rect 6748 27384 6776 27415
rect 7282 27412 7288 27424
rect 7340 27412 7346 27464
rect 7392 27461 7420 27492
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27421 7435 27455
rect 7377 27415 7435 27421
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 7558 27412 7564 27464
rect 7616 27412 7622 27464
rect 7760 27461 7788 27560
rect 8202 27548 8208 27600
rect 8260 27548 8266 27600
rect 8386 27548 8392 27600
rect 8444 27548 8450 27600
rect 9214 27548 9220 27600
rect 9272 27588 9278 27600
rect 12158 27588 12164 27600
rect 9272 27560 12164 27588
rect 9272 27548 9278 27560
rect 8220 27520 8248 27548
rect 8941 27523 8999 27529
rect 8941 27520 8953 27523
rect 8128 27492 8248 27520
rect 8496 27492 8953 27520
rect 7745 27455 7803 27461
rect 7745 27421 7757 27455
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 7837 27455 7895 27461
rect 7837 27421 7849 27455
rect 7883 27452 7895 27455
rect 7926 27452 7932 27464
rect 7883 27424 7932 27452
rect 7883 27421 7895 27424
rect 7837 27415 7895 27421
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 8128 27461 8156 27492
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8113 27415 8171 27421
rect 8202 27412 8208 27464
rect 8260 27412 8266 27464
rect 8021 27387 8079 27393
rect 5592 27356 7880 27384
rect 5592 27344 5598 27356
rect 5626 27316 5632 27328
rect 4724 27288 5632 27316
rect 5626 27276 5632 27288
rect 5684 27276 5690 27328
rect 5994 27276 6000 27328
rect 6052 27276 6058 27328
rect 6086 27276 6092 27328
rect 6144 27316 6150 27328
rect 6822 27316 6828 27328
rect 6144 27288 6828 27316
rect 6144 27276 6150 27288
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 6917 27319 6975 27325
rect 6917 27285 6929 27319
rect 6963 27316 6975 27319
rect 7190 27316 7196 27328
rect 6963 27288 7196 27316
rect 6963 27285 6975 27288
rect 6917 27279 6975 27285
rect 7190 27276 7196 27288
rect 7248 27316 7254 27328
rect 7742 27316 7748 27328
rect 7248 27288 7748 27316
rect 7248 27276 7254 27288
rect 7742 27276 7748 27288
rect 7800 27276 7806 27328
rect 7852 27316 7880 27356
rect 8021 27353 8033 27387
rect 8067 27384 8079 27387
rect 8496 27384 8524 27492
rect 8941 27489 8953 27492
rect 8987 27489 8999 27523
rect 8941 27483 8999 27489
rect 9048 27492 10088 27520
rect 8570 27412 8576 27464
rect 8628 27412 8634 27464
rect 8757 27455 8815 27461
rect 8757 27421 8769 27455
rect 8803 27452 8815 27455
rect 9048 27452 9076 27492
rect 8803 27424 9076 27452
rect 8803 27421 8815 27424
rect 8757 27415 8815 27421
rect 8067 27356 8524 27384
rect 8067 27353 8079 27356
rect 8021 27347 8079 27353
rect 8772 27316 8800 27415
rect 9122 27412 9128 27464
rect 9180 27412 9186 27464
rect 9214 27412 9220 27464
rect 9272 27412 9278 27464
rect 9401 27455 9459 27461
rect 9401 27421 9413 27455
rect 9447 27421 9459 27455
rect 9401 27415 9459 27421
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9416 27384 9444 27415
rect 9232 27356 9444 27384
rect 9232 27328 9260 27356
rect 7852 27288 8800 27316
rect 9214 27276 9220 27328
rect 9272 27276 9278 27328
rect 9508 27316 9536 27415
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 9953 27455 10011 27461
rect 9953 27452 9965 27455
rect 9640 27424 9965 27452
rect 9640 27412 9646 27424
rect 9953 27421 9965 27424
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10060 27384 10088 27492
rect 10226 27480 10232 27532
rect 10284 27480 10290 27532
rect 10134 27412 10140 27464
rect 10192 27412 10198 27464
rect 10612 27461 10640 27560
rect 12158 27548 12164 27560
rect 12216 27548 12222 27600
rect 12802 27588 12808 27600
rect 12268 27560 12808 27588
rect 12268 27529 12296 27560
rect 12802 27548 12808 27560
rect 12860 27548 12866 27600
rect 12894 27548 12900 27600
rect 12952 27588 12958 27600
rect 13081 27591 13139 27597
rect 13081 27588 13093 27591
rect 12952 27560 13093 27588
rect 12952 27548 12958 27560
rect 13081 27557 13093 27560
rect 13127 27557 13139 27591
rect 13081 27551 13139 27557
rect 13722 27548 13728 27600
rect 13780 27548 13786 27600
rect 15010 27588 15016 27600
rect 14016 27560 15016 27588
rect 11425 27523 11483 27529
rect 11425 27520 11437 27523
rect 10796 27492 11437 27520
rect 10796 27461 10824 27492
rect 11425 27489 11437 27492
rect 11471 27489 11483 27523
rect 11425 27483 11483 27489
rect 12253 27523 12311 27529
rect 12253 27489 12265 27523
rect 12299 27489 12311 27523
rect 12912 27520 12940 27548
rect 12253 27483 12311 27489
rect 12452 27492 12940 27520
rect 12989 27523 13047 27529
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27421 10563 27455
rect 10505 27415 10563 27421
rect 10597 27455 10655 27461
rect 10597 27421 10609 27455
rect 10643 27421 10655 27455
rect 10597 27415 10655 27421
rect 10781 27455 10839 27461
rect 10781 27421 10793 27455
rect 10827 27421 10839 27455
rect 10781 27415 10839 27421
rect 10873 27455 10931 27461
rect 10873 27421 10885 27455
rect 10919 27452 10931 27455
rect 11054 27452 11060 27464
rect 10919 27424 11060 27452
rect 10919 27421 10931 27424
rect 10873 27415 10931 27421
rect 10410 27384 10416 27396
rect 10060 27356 10416 27384
rect 10410 27344 10416 27356
rect 10468 27344 10474 27396
rect 10520 27384 10548 27415
rect 10686 27384 10692 27396
rect 10520 27356 10692 27384
rect 10686 27344 10692 27356
rect 10744 27344 10750 27396
rect 9674 27316 9680 27328
rect 9508 27288 9680 27316
rect 9674 27276 9680 27288
rect 9732 27316 9738 27328
rect 10888 27316 10916 27415
rect 11054 27412 11060 27424
rect 11112 27412 11118 27464
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27452 11207 27455
rect 11238 27452 11244 27464
rect 11195 27424 11244 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 12452 27461 12480 27492
rect 12989 27489 13001 27523
rect 13035 27520 13047 27523
rect 13740 27520 13768 27548
rect 14016 27532 14044 27560
rect 15010 27548 15016 27560
rect 15068 27548 15074 27600
rect 18984 27588 19012 27616
rect 20990 27588 20996 27600
rect 18984 27560 20996 27588
rect 20990 27548 20996 27560
rect 21048 27548 21054 27600
rect 21174 27548 21180 27600
rect 21232 27588 21238 27600
rect 21453 27591 21511 27597
rect 21453 27588 21465 27591
rect 21232 27560 21465 27588
rect 21232 27548 21238 27560
rect 21453 27557 21465 27560
rect 21499 27557 21511 27591
rect 21453 27551 21511 27557
rect 22097 27591 22155 27597
rect 22097 27557 22109 27591
rect 22143 27557 22155 27591
rect 22097 27551 22155 27557
rect 13035 27492 13768 27520
rect 13035 27489 13047 27492
rect 12989 27483 13047 27489
rect 13998 27480 14004 27532
rect 14056 27480 14062 27532
rect 19426 27480 19432 27532
rect 19484 27520 19490 27532
rect 19797 27523 19855 27529
rect 19797 27520 19809 27523
rect 19484 27492 19809 27520
rect 19484 27480 19490 27492
rect 19797 27489 19809 27492
rect 19843 27489 19855 27523
rect 19797 27483 19855 27489
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 21637 27523 21695 27529
rect 21637 27520 21649 27523
rect 20772 27492 21649 27520
rect 20772 27480 20778 27492
rect 21637 27489 21649 27492
rect 21683 27489 21695 27523
rect 22112 27520 22140 27551
rect 23382 27548 23388 27600
rect 23440 27588 23446 27600
rect 23477 27591 23535 27597
rect 23477 27588 23489 27591
rect 23440 27560 23489 27588
rect 23440 27548 23446 27560
rect 23477 27557 23489 27560
rect 23523 27557 23535 27591
rect 23477 27551 23535 27557
rect 24486 27548 24492 27600
rect 24544 27588 24550 27600
rect 24765 27591 24823 27597
rect 24765 27588 24777 27591
rect 24544 27560 24777 27588
rect 24544 27548 24550 27560
rect 24765 27557 24777 27560
rect 24811 27557 24823 27591
rect 24765 27551 24823 27557
rect 23566 27520 23572 27532
rect 22112 27492 23572 27520
rect 21637 27483 21695 27489
rect 23566 27480 23572 27492
rect 23624 27480 23630 27532
rect 25041 27523 25099 27529
rect 25041 27520 25053 27523
rect 23768 27492 25053 27520
rect 23768 27464 23796 27492
rect 25041 27489 25053 27492
rect 25087 27489 25099 27523
rect 25041 27483 25099 27489
rect 11333 27455 11391 27461
rect 11333 27421 11345 27455
rect 11379 27452 11391 27455
rect 12437 27455 12495 27461
rect 11379 27424 11468 27452
rect 11379 27421 11391 27424
rect 11333 27415 11391 27421
rect 10965 27387 11023 27393
rect 10965 27353 10977 27387
rect 11011 27384 11023 27387
rect 11011 27356 11376 27384
rect 11011 27353 11023 27356
rect 10965 27347 11023 27353
rect 11348 27328 11376 27356
rect 11440 27328 11468 27424
rect 12437 27421 12449 27455
rect 12483 27421 12495 27455
rect 12437 27415 12495 27421
rect 12529 27455 12587 27461
rect 12529 27421 12541 27455
rect 12575 27421 12587 27455
rect 12529 27415 12587 27421
rect 11977 27387 12035 27393
rect 11977 27353 11989 27387
rect 12023 27384 12035 27387
rect 12544 27384 12572 27415
rect 12618 27412 12624 27464
rect 12676 27452 12682 27464
rect 12897 27455 12955 27461
rect 12897 27452 12909 27455
rect 12676 27424 12909 27452
rect 12676 27412 12682 27424
rect 12897 27421 12909 27424
rect 12943 27421 12955 27455
rect 12897 27415 12955 27421
rect 12023 27356 12572 27384
rect 12912 27384 12940 27415
rect 13170 27412 13176 27464
rect 13228 27412 13234 27464
rect 13262 27412 13268 27464
rect 13320 27452 13326 27464
rect 14185 27455 14243 27461
rect 14185 27452 14197 27455
rect 13320 27424 14197 27452
rect 13320 27412 13326 27424
rect 14185 27421 14197 27424
rect 14231 27421 14243 27455
rect 14185 27415 14243 27421
rect 14274 27412 14280 27464
rect 14332 27452 14338 27464
rect 14369 27455 14427 27461
rect 14369 27452 14381 27455
rect 14332 27424 14381 27452
rect 14332 27412 14338 27424
rect 14369 27421 14381 27424
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 14608 27424 14872 27452
rect 14608 27412 14614 27424
rect 13280 27384 13308 27412
rect 12912 27356 13308 27384
rect 13357 27387 13415 27393
rect 12023 27353 12035 27356
rect 11977 27347 12035 27353
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 14292 27384 14320 27412
rect 13403 27356 14320 27384
rect 14645 27387 14703 27393
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 14645 27353 14657 27387
rect 14691 27384 14703 27387
rect 14734 27384 14740 27396
rect 14691 27356 14740 27384
rect 14691 27353 14703 27356
rect 14645 27347 14703 27353
rect 14734 27344 14740 27356
rect 14792 27344 14798 27396
rect 14844 27384 14872 27424
rect 14918 27412 14924 27464
rect 14976 27452 14982 27464
rect 15197 27455 15255 27461
rect 15197 27452 15209 27455
rect 14976 27424 15209 27452
rect 14976 27412 14982 27424
rect 15197 27421 15209 27424
rect 15243 27452 15255 27455
rect 17218 27452 17224 27464
rect 15243 27424 17224 27452
rect 15243 27421 15255 27424
rect 15197 27415 15255 27421
rect 17218 27412 17224 27424
rect 17276 27412 17282 27464
rect 17488 27455 17546 27461
rect 17488 27421 17500 27455
rect 17534 27452 17546 27455
rect 17862 27452 17868 27464
rect 17534 27424 17868 27452
rect 17534 27421 17546 27424
rect 17488 27415 17546 27421
rect 17862 27412 17868 27424
rect 17920 27412 17926 27464
rect 17972 27424 19840 27452
rect 15464 27387 15522 27393
rect 14844 27356 15424 27384
rect 9732 27288 10916 27316
rect 9732 27276 9738 27288
rect 11330 27276 11336 27328
rect 11388 27276 11394 27328
rect 11422 27276 11428 27328
rect 11480 27276 11486 27328
rect 12069 27319 12127 27325
rect 12069 27285 12081 27319
rect 12115 27316 12127 27319
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 12115 27288 12725 27316
rect 12115 27285 12127 27288
rect 12069 27279 12127 27285
rect 12713 27285 12725 27288
rect 12759 27285 12771 27319
rect 12713 27279 12771 27285
rect 13262 27276 13268 27328
rect 13320 27316 13326 27328
rect 15286 27316 15292 27328
rect 13320 27288 15292 27316
rect 13320 27276 13326 27288
rect 15286 27276 15292 27288
rect 15344 27276 15350 27328
rect 15396 27316 15424 27356
rect 15464 27353 15476 27387
rect 15510 27384 15522 27387
rect 16206 27384 16212 27396
rect 15510 27356 16212 27384
rect 15510 27353 15522 27356
rect 15464 27347 15522 27353
rect 16206 27344 16212 27356
rect 16264 27344 16270 27396
rect 17972 27384 18000 27424
rect 16307 27356 18000 27384
rect 16307 27316 16335 27356
rect 18046 27344 18052 27396
rect 18104 27384 18110 27396
rect 19705 27387 19763 27393
rect 19705 27384 19717 27387
rect 18104 27356 19717 27384
rect 18104 27344 18110 27356
rect 19705 27353 19717 27356
rect 19751 27353 19763 27387
rect 19812 27384 19840 27424
rect 20070 27412 20076 27464
rect 20128 27412 20134 27464
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27452 20959 27455
rect 21082 27452 21088 27464
rect 20947 27424 21088 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 20916 27384 20944 27415
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 21729 27455 21787 27461
rect 21729 27452 21741 27455
rect 21324 27424 21741 27452
rect 21324 27412 21330 27424
rect 21729 27421 21741 27424
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 23750 27412 23756 27464
rect 23808 27412 23814 27464
rect 24026 27452 24032 27464
rect 23860 27424 24032 27452
rect 19812 27356 20944 27384
rect 19705 27347 19763 27353
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 22922 27344 22928 27396
rect 22980 27384 22986 27396
rect 23860 27384 23888 27424
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 24578 27412 24584 27464
rect 24636 27412 24642 27464
rect 24857 27455 24915 27461
rect 24857 27421 24869 27455
rect 24903 27452 24915 27455
rect 25155 27452 25183 27628
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 27264 27588 27292 27628
rect 27338 27616 27344 27668
rect 27396 27656 27402 27668
rect 28074 27656 28080 27668
rect 27396 27628 28080 27656
rect 27396 27616 27402 27628
rect 28074 27616 28080 27628
rect 28132 27616 28138 27668
rect 28718 27616 28724 27668
rect 28776 27616 28782 27668
rect 30190 27656 30196 27668
rect 30024 27628 30196 27656
rect 29822 27588 29828 27600
rect 26384 27560 27016 27588
rect 27264 27560 27660 27588
rect 26384 27548 26390 27560
rect 25314 27480 25320 27532
rect 25372 27480 25378 27532
rect 26418 27520 26424 27532
rect 25608 27492 26424 27520
rect 24903 27424 25183 27452
rect 25225 27455 25283 27461
rect 24903 27421 24915 27424
rect 24857 27415 24915 27421
rect 25225 27421 25237 27455
rect 25271 27452 25283 27455
rect 25332 27452 25360 27480
rect 25608 27464 25636 27492
rect 25271 27424 25360 27452
rect 25271 27421 25283 27424
rect 25225 27415 25283 27421
rect 25590 27412 25596 27464
rect 25648 27412 25654 27464
rect 26050 27412 26056 27464
rect 26108 27412 26114 27464
rect 26068 27384 26096 27412
rect 22980 27356 23888 27384
rect 23952 27356 26096 27384
rect 22980 27344 22986 27356
rect 15396 27288 16335 27316
rect 17402 27276 17408 27328
rect 17460 27316 17466 27328
rect 18601 27319 18659 27325
rect 18601 27316 18613 27319
rect 17460 27288 18613 27316
rect 17460 27276 17466 27288
rect 18601 27285 18613 27288
rect 18647 27285 18659 27319
rect 18601 27279 18659 27285
rect 19242 27276 19248 27328
rect 19300 27276 19306 27328
rect 19426 27276 19432 27328
rect 19484 27316 19490 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 19484 27288 19625 27316
rect 19484 27276 19490 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19613 27279 19671 27285
rect 20714 27276 20720 27328
rect 20772 27276 20778 27328
rect 21634 27276 21640 27328
rect 21692 27316 21698 27328
rect 23952 27316 23980 27356
rect 21692 27288 23980 27316
rect 21692 27276 21698 27288
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 25409 27319 25467 27325
rect 25409 27285 25421 27319
rect 25455 27316 25467 27319
rect 25590 27316 25596 27328
rect 25455 27288 25596 27316
rect 25455 27285 25467 27288
rect 25409 27279 25467 27285
rect 25590 27276 25596 27288
rect 25648 27276 25654 27328
rect 26050 27276 26056 27328
rect 26108 27276 26114 27328
rect 26160 27316 26188 27492
rect 26418 27480 26424 27492
rect 26476 27480 26482 27532
rect 26988 27520 27016 27560
rect 27632 27520 27660 27560
rect 28920 27560 29828 27588
rect 28718 27520 28724 27532
rect 26988 27492 27108 27520
rect 27632 27492 28724 27520
rect 26510 27412 26516 27464
rect 26568 27462 26574 27464
rect 26568 27461 26740 27462
rect 26568 27455 26755 27461
rect 26568 27434 26709 27455
rect 26568 27412 26574 27434
rect 26697 27421 26709 27434
rect 26743 27421 26755 27455
rect 26697 27415 26755 27421
rect 26786 27412 26792 27464
rect 26844 27412 26850 27464
rect 27080 27461 27108 27492
rect 28718 27480 28724 27492
rect 28776 27480 28782 27532
rect 26881 27455 26939 27461
rect 26881 27421 26893 27455
rect 26927 27449 26939 27455
rect 27065 27455 27123 27461
rect 26927 27446 26944 27449
rect 26927 27421 27016 27446
rect 26881 27418 27016 27421
rect 26881 27415 26939 27418
rect 26418 27344 26424 27396
rect 26476 27344 26482 27396
rect 26988 27316 27016 27418
rect 27065 27421 27077 27455
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 27338 27412 27344 27464
rect 27396 27412 27402 27464
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 27246 27344 27252 27396
rect 27304 27384 27310 27396
rect 27448 27384 27476 27415
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 27580 27424 27629 27452
rect 27580 27412 27586 27424
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 27709 27455 27767 27461
rect 27709 27421 27721 27455
rect 27755 27452 27767 27455
rect 27985 27455 28043 27461
rect 27755 27424 27936 27452
rect 27755 27421 27767 27424
rect 27709 27415 27767 27421
rect 27908 27396 27936 27424
rect 27985 27421 27997 27455
rect 28031 27452 28043 27455
rect 28074 27452 28080 27464
rect 28031 27424 28080 27452
rect 28031 27421 28043 27424
rect 27985 27415 28043 27421
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28166 27412 28172 27464
rect 28224 27412 28230 27464
rect 28920 27461 28948 27560
rect 29822 27548 29828 27560
rect 29880 27548 29886 27600
rect 29365 27523 29423 27529
rect 29365 27489 29377 27523
rect 29411 27520 29423 27523
rect 30024 27520 30052 27628
rect 30190 27616 30196 27628
rect 30248 27616 30254 27668
rect 31018 27656 31024 27668
rect 30300 27628 31024 27656
rect 30300 27520 30328 27628
rect 31018 27616 31024 27628
rect 31076 27656 31082 27668
rect 31076 27628 31156 27656
rect 31076 27616 31082 27628
rect 30558 27548 30564 27600
rect 30616 27548 30622 27600
rect 29411 27492 30052 27520
rect 30116 27492 30328 27520
rect 29411 27489 29423 27492
rect 29365 27483 29423 27489
rect 28905 27455 28963 27461
rect 28905 27421 28917 27455
rect 28951 27421 28963 27455
rect 28905 27415 28963 27421
rect 28994 27412 29000 27464
rect 29052 27412 29058 27464
rect 30116 27461 30144 27492
rect 29227 27455 29285 27461
rect 29227 27421 29239 27455
rect 29273 27452 29285 27455
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 29273 27424 30113 27452
rect 29273 27421 29285 27424
rect 29227 27415 29285 27421
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 30282 27412 30288 27464
rect 30340 27412 30346 27464
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27452 30435 27455
rect 30576 27452 30604 27548
rect 30423 27424 30604 27452
rect 30423 27421 30435 27424
rect 30377 27415 30435 27421
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30742 27412 30748 27464
rect 30800 27452 30806 27464
rect 30837 27455 30895 27461
rect 30837 27452 30849 27455
rect 30800 27424 30849 27452
rect 30800 27412 30806 27424
rect 30837 27421 30849 27424
rect 30883 27421 30895 27455
rect 30837 27415 30895 27421
rect 30926 27412 30932 27464
rect 30984 27412 30990 27464
rect 31021 27455 31079 27461
rect 31021 27421 31033 27455
rect 31067 27452 31079 27455
rect 31128 27452 31156 27628
rect 31202 27616 31208 27668
rect 31260 27656 31266 27668
rect 34054 27656 34060 27668
rect 31260 27628 34060 27656
rect 31260 27616 31266 27628
rect 34054 27616 34060 27628
rect 34112 27616 34118 27668
rect 31754 27588 31760 27600
rect 31404 27560 31760 27588
rect 31404 27529 31432 27560
rect 31754 27548 31760 27560
rect 31812 27548 31818 27600
rect 32677 27591 32735 27597
rect 32677 27588 32689 27591
rect 32140 27560 32689 27588
rect 31389 27523 31447 27529
rect 31389 27489 31401 27523
rect 31435 27489 31447 27523
rect 32140 27520 32168 27560
rect 32677 27557 32689 27560
rect 32723 27588 32735 27591
rect 32723 27560 32812 27588
rect 32723 27557 32735 27560
rect 32677 27551 32735 27557
rect 31389 27483 31447 27489
rect 31496 27492 32168 27520
rect 32784 27520 32812 27560
rect 33042 27548 33048 27600
rect 33100 27588 33106 27600
rect 33321 27591 33379 27597
rect 33321 27588 33333 27591
rect 33100 27560 33333 27588
rect 33100 27548 33106 27560
rect 33321 27557 33333 27560
rect 33367 27557 33379 27591
rect 33321 27551 33379 27557
rect 32784 27492 32996 27520
rect 31496 27464 31524 27492
rect 31067 27424 31156 27452
rect 31067 27421 31079 27424
rect 31021 27415 31079 27421
rect 27304 27356 27476 27384
rect 27801 27387 27859 27393
rect 27304 27344 27310 27356
rect 27801 27353 27813 27387
rect 27847 27353 27859 27387
rect 27801 27347 27859 27353
rect 26160 27288 27016 27316
rect 27154 27276 27160 27328
rect 27212 27276 27218 27328
rect 27816 27316 27844 27347
rect 27890 27344 27896 27396
rect 27948 27344 27954 27396
rect 28184 27384 28212 27412
rect 28000 27356 28212 27384
rect 29089 27387 29147 27393
rect 28000 27316 28028 27356
rect 29089 27353 29101 27387
rect 29135 27384 29147 27387
rect 29362 27384 29368 27396
rect 29135 27356 29368 27384
rect 29135 27353 29147 27356
rect 29089 27347 29147 27353
rect 29362 27344 29368 27356
rect 29420 27344 29426 27396
rect 29822 27344 29828 27396
rect 29880 27384 29886 27396
rect 30668 27384 30696 27412
rect 29880 27356 30696 27384
rect 31036 27384 31064 27415
rect 31478 27412 31484 27464
rect 31536 27412 31542 27464
rect 31938 27412 31944 27464
rect 31996 27412 32002 27464
rect 32125 27455 32183 27461
rect 32125 27421 32137 27455
rect 32171 27452 32183 27455
rect 32171 27424 32444 27452
rect 32171 27421 32183 27424
rect 32125 27415 32183 27421
rect 32416 27384 32444 27424
rect 32674 27412 32680 27464
rect 32732 27452 32738 27464
rect 32769 27455 32827 27461
rect 32769 27452 32781 27455
rect 32732 27424 32781 27452
rect 32732 27412 32738 27424
rect 32769 27421 32781 27424
rect 32815 27421 32827 27455
rect 32968 27452 32996 27492
rect 33226 27480 33232 27532
rect 33284 27520 33290 27532
rect 33284 27492 33640 27520
rect 33284 27480 33290 27492
rect 33612 27461 33640 27492
rect 33045 27455 33103 27461
rect 33045 27452 33057 27455
rect 32968 27424 33057 27452
rect 32769 27415 32827 27421
rect 33045 27421 33057 27424
rect 33091 27421 33103 27455
rect 33045 27415 33103 27421
rect 33137 27455 33195 27461
rect 33137 27421 33149 27455
rect 33183 27421 33195 27455
rect 33137 27415 33195 27421
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27421 33563 27455
rect 33505 27415 33563 27421
rect 33597 27455 33655 27461
rect 33597 27421 33609 27455
rect 33643 27421 33655 27455
rect 33597 27415 33655 27421
rect 32582 27384 32588 27396
rect 31036 27356 32343 27384
rect 32416 27356 32588 27384
rect 29880 27344 29886 27356
rect 27816 27288 28028 27316
rect 28166 27276 28172 27328
rect 28224 27276 28230 27328
rect 29730 27276 29736 27328
rect 29788 27276 29794 27328
rect 29917 27319 29975 27325
rect 29917 27285 29929 27319
rect 29963 27316 29975 27319
rect 31018 27316 31024 27328
rect 29963 27288 31024 27316
rect 29963 27285 29975 27288
rect 29917 27279 29975 27285
rect 31018 27276 31024 27288
rect 31076 27276 31082 27328
rect 31205 27319 31263 27325
rect 31205 27285 31217 27319
rect 31251 27316 31263 27319
rect 32214 27316 32220 27328
rect 31251 27288 32220 27316
rect 31251 27285 31263 27288
rect 31205 27279 31263 27285
rect 32214 27276 32220 27288
rect 32272 27276 32278 27328
rect 32315 27316 32343 27356
rect 32582 27344 32588 27356
rect 32640 27344 32646 27396
rect 32950 27344 32956 27396
rect 33008 27344 33014 27396
rect 33152 27316 33180 27415
rect 33520 27384 33548 27415
rect 34054 27384 34060 27396
rect 33520 27356 34060 27384
rect 34054 27344 34060 27356
rect 34112 27344 34118 27396
rect 32315 27288 33180 27316
rect 33778 27276 33784 27328
rect 33836 27276 33842 27328
rect 1104 27226 43884 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 43884 27226
rect 1104 27152 43884 27174
rect 2866 27072 2872 27124
rect 2924 27112 2930 27124
rect 3237 27115 3295 27121
rect 3237 27112 3249 27115
rect 2924 27084 3249 27112
rect 2924 27072 2930 27084
rect 3237 27081 3249 27084
rect 3283 27081 3295 27115
rect 3237 27075 3295 27081
rect 3418 27072 3424 27124
rect 3476 27072 3482 27124
rect 4154 27112 4160 27124
rect 3620 27084 4160 27112
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26976 1639 26979
rect 3418 26976 3424 26988
rect 1627 26948 3424 26976
rect 1627 26945 1639 26948
rect 1581 26939 1639 26945
rect 3418 26936 3424 26948
rect 3476 26936 3482 26988
rect 3620 26985 3648 27084
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 4798 27112 4804 27124
rect 4633 27084 4804 27112
rect 3973 27047 4031 27053
rect 3973 27013 3985 27047
rect 4019 27044 4031 27047
rect 4430 27044 4436 27056
rect 4019 27016 4436 27044
rect 4019 27013 4031 27016
rect 3973 27007 4031 27013
rect 3605 26979 3663 26985
rect 3605 26945 3617 26979
rect 3651 26945 3663 26979
rect 3605 26939 3663 26945
rect 3786 26936 3792 26988
rect 3844 26936 3850 26988
rect 3881 26979 3939 26985
rect 3881 26945 3893 26979
rect 3927 26976 3939 26979
rect 3988 26976 4016 27007
rect 4430 27004 4436 27016
rect 4488 27004 4494 27056
rect 3927 26948 4016 26976
rect 3927 26945 3939 26948
rect 3881 26939 3939 26945
rect 4062 26936 4068 26988
rect 4120 26976 4126 26988
rect 4157 26979 4215 26985
rect 4157 26976 4169 26979
rect 4120 26948 4169 26976
rect 4120 26936 4126 26948
rect 4157 26945 4169 26948
rect 4203 26945 4215 26979
rect 4157 26939 4215 26945
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 4633 26976 4661 27084
rect 4798 27072 4804 27084
rect 4856 27072 4862 27124
rect 4982 27072 4988 27124
rect 5040 27112 5046 27124
rect 5175 27115 5233 27121
rect 5175 27112 5187 27115
rect 5040 27084 5187 27112
rect 5040 27072 5046 27084
rect 5175 27081 5187 27084
rect 5221 27081 5233 27115
rect 6086 27112 6092 27124
rect 5175 27075 5233 27081
rect 5460 27084 6092 27112
rect 4706 27004 4712 27056
rect 4764 27044 4770 27056
rect 5460 27044 5488 27084
rect 6086 27072 6092 27084
rect 6144 27112 6150 27124
rect 6181 27115 6239 27121
rect 6181 27112 6193 27115
rect 6144 27084 6193 27112
rect 6144 27072 6150 27084
rect 6181 27081 6193 27084
rect 6227 27081 6239 27115
rect 6181 27075 6239 27081
rect 6270 27072 6276 27124
rect 6328 27112 6334 27124
rect 8202 27112 8208 27124
rect 6328 27084 8208 27112
rect 6328 27072 6334 27084
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 8294 27072 8300 27124
rect 8352 27072 8358 27124
rect 8570 27072 8576 27124
rect 8628 27072 8634 27124
rect 8849 27115 8907 27121
rect 8849 27081 8861 27115
rect 8895 27112 8907 27115
rect 8938 27112 8944 27124
rect 8895 27084 8944 27112
rect 8895 27081 8907 27084
rect 8849 27075 8907 27081
rect 8938 27072 8944 27084
rect 8996 27072 9002 27124
rect 9122 27072 9128 27124
rect 9180 27112 9186 27124
rect 9309 27115 9367 27121
rect 9309 27112 9321 27115
rect 9180 27084 9321 27112
rect 9180 27072 9186 27084
rect 9309 27081 9321 27084
rect 9355 27081 9367 27115
rect 9309 27075 9367 27081
rect 9490 27072 9496 27124
rect 9548 27112 9554 27124
rect 9677 27115 9735 27121
rect 9677 27112 9689 27115
rect 9548 27084 9689 27112
rect 9548 27072 9554 27084
rect 9677 27081 9689 27084
rect 9723 27081 9735 27115
rect 9677 27075 9735 27081
rect 10134 27072 10140 27124
rect 10192 27112 10198 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 10192 27084 10609 27112
rect 10192 27072 10198 27084
rect 10597 27081 10609 27084
rect 10643 27081 10655 27115
rect 10597 27075 10655 27081
rect 10686 27072 10692 27124
rect 10744 27112 10750 27124
rect 10781 27115 10839 27121
rect 10781 27112 10793 27115
rect 10744 27084 10793 27112
rect 10744 27072 10750 27084
rect 10781 27081 10793 27084
rect 10827 27081 10839 27115
rect 10781 27075 10839 27081
rect 11149 27115 11207 27121
rect 11149 27081 11161 27115
rect 11195 27112 11207 27115
rect 11238 27112 11244 27124
rect 11195 27084 11244 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 11514 27072 11520 27124
rect 11572 27112 11578 27124
rect 12345 27115 12403 27121
rect 11572 27084 11892 27112
rect 11572 27072 11578 27084
rect 4764 27016 5028 27044
rect 4764 27004 4770 27016
rect 4295 26948 4384 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 4356 26920 4384 26948
rect 4448 26948 4661 26976
rect 1854 26868 1860 26920
rect 1912 26868 1918 26920
rect 3510 26868 3516 26920
rect 3568 26908 3574 26920
rect 3568 26880 4016 26908
rect 3568 26868 3574 26880
rect 3988 26849 4016 26880
rect 4338 26868 4344 26920
rect 4396 26868 4402 26920
rect 4448 26917 4476 26948
rect 4798 26936 4804 26988
rect 4856 26936 4862 26988
rect 4899 26985 4927 27016
rect 4893 26979 4951 26985
rect 4893 26945 4905 26979
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 5000 26920 5028 27016
rect 5288 27016 5488 27044
rect 5813 27047 5871 27053
rect 5288 26988 5316 27016
rect 5813 27013 5825 27047
rect 5859 27044 5871 27047
rect 6641 27047 6699 27053
rect 6641 27044 6653 27047
rect 5859 27016 6653 27044
rect 5859 27013 5871 27016
rect 5813 27007 5871 27013
rect 6641 27013 6653 27016
rect 6687 27044 6699 27047
rect 6687 27016 7604 27044
rect 6687 27013 6699 27016
rect 6641 27007 6699 27013
rect 7576 26988 7604 27016
rect 7650 27004 7656 27056
rect 7708 27044 7714 27056
rect 8588 27044 8616 27072
rect 7708 27016 8432 27044
rect 8588 27016 9076 27044
rect 7708 27004 7714 27016
rect 5077 26979 5135 26985
rect 5077 26945 5089 26979
rect 5123 26976 5135 26979
rect 5166 26976 5172 26988
rect 5123 26948 5172 26976
rect 5123 26945 5135 26948
rect 5077 26939 5135 26945
rect 5166 26936 5172 26948
rect 5224 26936 5230 26988
rect 5258 26936 5264 26988
rect 5316 26936 5322 26988
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26976 5411 26979
rect 5399 26948 5488 26976
rect 5399 26945 5411 26948
rect 5353 26939 5411 26945
rect 5460 26920 5488 26948
rect 5534 26936 5540 26988
rect 5592 26936 5598 26988
rect 5718 26985 5724 26988
rect 5685 26979 5724 26985
rect 5685 26945 5697 26979
rect 5685 26939 5724 26945
rect 5718 26936 5724 26939
rect 5776 26936 5782 26988
rect 5902 26936 5908 26988
rect 5960 26936 5966 26988
rect 6043 26979 6101 26985
rect 6043 26945 6055 26979
rect 6089 26945 6101 26979
rect 6043 26939 6101 26945
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26877 4491 26911
rect 4433 26871 4491 26877
rect 4617 26911 4675 26917
rect 4617 26877 4629 26911
rect 4663 26877 4675 26911
rect 4617 26871 4675 26877
rect 4709 26911 4767 26917
rect 4709 26877 4721 26911
rect 4755 26877 4767 26911
rect 4709 26871 4767 26877
rect 3973 26843 4031 26849
rect 3973 26809 3985 26843
rect 4019 26809 4031 26843
rect 3973 26803 4031 26809
rect 4632 26772 4660 26871
rect 4724 26840 4752 26871
rect 4982 26868 4988 26920
rect 5040 26868 5046 26920
rect 5442 26868 5448 26920
rect 5500 26868 5506 26920
rect 6058 26908 6086 26939
rect 6362 26936 6368 26988
rect 6420 26936 6426 26988
rect 6454 26936 6460 26988
rect 6512 26976 6518 26988
rect 6512 26948 6557 26976
rect 6512 26936 6518 26948
rect 6730 26936 6736 26988
rect 6788 26936 6794 26988
rect 6822 26936 6828 26988
rect 6880 26985 6886 26988
rect 6880 26979 6929 26985
rect 6880 26945 6883 26979
rect 6917 26976 6929 26979
rect 6917 26948 6973 26976
rect 6917 26945 6929 26948
rect 6880 26939 6929 26945
rect 6880 26936 6886 26939
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 7852 26985 7880 27016
rect 8404 26988 8432 27016
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26945 7895 26979
rect 7837 26939 7895 26945
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26976 7987 26979
rect 7975 26948 8156 26976
rect 7975 26945 7987 26948
rect 7929 26939 7987 26945
rect 6840 26908 6868 26936
rect 6058 26880 6868 26908
rect 7282 26868 7288 26920
rect 7340 26908 7346 26920
rect 7653 26911 7711 26917
rect 7653 26908 7665 26911
rect 7340 26880 7665 26908
rect 7340 26868 7346 26880
rect 7653 26877 7665 26880
rect 7699 26908 7711 26911
rect 8018 26908 8024 26920
rect 7699 26880 8024 26908
rect 7699 26877 7711 26880
rect 7653 26871 7711 26877
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 4798 26840 4804 26852
rect 4724 26812 4804 26840
rect 4798 26800 4804 26812
rect 4856 26800 4862 26852
rect 5166 26800 5172 26852
rect 5224 26840 5230 26852
rect 8128 26840 8156 26948
rect 8386 26936 8392 26988
rect 8444 26936 8450 26988
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 8662 26976 8668 26988
rect 8527 26948 8668 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 8662 26936 8668 26948
rect 8720 26936 8726 26988
rect 8754 26936 8760 26988
rect 8812 26936 8818 26988
rect 8846 26936 8852 26988
rect 8904 26936 8910 26988
rect 9048 26985 9076 27016
rect 9214 27004 9220 27056
rect 9272 27004 9278 27056
rect 11422 27044 11428 27056
rect 9646 27016 11428 27044
rect 9033 26979 9091 26985
rect 9033 26945 9045 26979
rect 9079 26976 9091 26979
rect 9493 26979 9551 26985
rect 9493 26976 9505 26979
rect 9079 26948 9505 26976
rect 9079 26945 9091 26948
rect 9033 26939 9091 26945
rect 9493 26945 9505 26948
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 8864 26908 8892 26936
rect 8352 26880 8892 26908
rect 9125 26911 9183 26917
rect 8352 26868 8358 26880
rect 9125 26877 9137 26911
rect 9171 26908 9183 26911
rect 9646 26908 9674 27016
rect 11422 27004 11428 27016
rect 11480 27004 11486 27056
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26945 9827 26979
rect 9769 26939 9827 26945
rect 10505 26979 10563 26985
rect 10505 26945 10517 26979
rect 10551 26945 10563 26979
rect 10505 26939 10563 26945
rect 9171 26880 9674 26908
rect 9171 26877 9183 26880
rect 9125 26871 9183 26877
rect 5224 26812 8156 26840
rect 5224 26800 5230 26812
rect 5442 26772 5448 26784
rect 4632 26744 5448 26772
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 6178 26732 6184 26784
rect 6236 26772 6242 26784
rect 6454 26772 6460 26784
rect 6236 26744 6460 26772
rect 6236 26732 6242 26744
rect 6454 26732 6460 26744
rect 6512 26732 6518 26784
rect 7006 26732 7012 26784
rect 7064 26732 7070 26784
rect 7466 26732 7472 26784
rect 7524 26732 7530 26784
rect 8128 26772 8156 26812
rect 8754 26800 8760 26852
rect 8812 26840 8818 26852
rect 9306 26840 9312 26852
rect 8812 26812 9312 26840
rect 8812 26800 8818 26812
rect 9306 26800 9312 26812
rect 9364 26840 9370 26852
rect 9784 26840 9812 26939
rect 10520 26908 10548 26939
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 10689 26979 10747 26985
rect 10689 26976 10701 26979
rect 10652 26948 10701 26976
rect 10652 26936 10658 26948
rect 10689 26945 10701 26948
rect 10735 26945 10747 26979
rect 10689 26939 10747 26945
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26976 11023 26979
rect 11146 26976 11152 26988
rect 11011 26948 11152 26976
rect 11011 26945 11023 26948
rect 10965 26939 11023 26945
rect 10980 26908 11008 26939
rect 11146 26936 11152 26948
rect 11204 26936 11210 26988
rect 11241 26979 11299 26985
rect 11241 26945 11253 26979
rect 11287 26945 11299 26979
rect 11241 26939 11299 26945
rect 10520 26880 11008 26908
rect 11256 26908 11284 26939
rect 11330 26908 11336 26920
rect 11256 26880 11336 26908
rect 11330 26868 11336 26880
rect 11388 26868 11394 26920
rect 9364 26812 9812 26840
rect 9364 26800 9370 26812
rect 9674 26772 9680 26784
rect 8128 26744 9680 26772
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 11440 26772 11468 27004
rect 11698 26936 11704 26988
rect 11756 26936 11762 26988
rect 11864 26985 11892 27084
rect 12345 27081 12357 27115
rect 12391 27112 12403 27115
rect 12802 27112 12808 27124
rect 12391 27084 12808 27112
rect 12391 27081 12403 27084
rect 12345 27075 12403 27081
rect 12802 27072 12808 27084
rect 12860 27072 12866 27124
rect 13170 27072 13176 27124
rect 13228 27112 13234 27124
rect 13449 27115 13507 27121
rect 13449 27112 13461 27115
rect 13228 27084 13461 27112
rect 13228 27072 13234 27084
rect 13449 27081 13461 27084
rect 13495 27081 13507 27115
rect 13449 27075 13507 27081
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 13817 27115 13875 27121
rect 13817 27112 13829 27115
rect 13596 27084 13829 27112
rect 13596 27072 13602 27084
rect 13817 27081 13829 27084
rect 13863 27112 13875 27115
rect 14458 27112 14464 27124
rect 13863 27084 14464 27112
rect 13863 27081 13875 27084
rect 13817 27075 13875 27081
rect 14458 27072 14464 27084
rect 14516 27072 14522 27124
rect 15289 27115 15347 27121
rect 15289 27081 15301 27115
rect 15335 27112 15347 27115
rect 15562 27112 15568 27124
rect 15335 27084 15568 27112
rect 15335 27081 15347 27084
rect 15289 27075 15347 27081
rect 15562 27072 15568 27084
rect 15620 27072 15626 27124
rect 17126 27072 17132 27124
rect 17184 27072 17190 27124
rect 18046 27072 18052 27124
rect 18104 27072 18110 27124
rect 18322 27072 18328 27124
rect 18380 27112 18386 27124
rect 18509 27115 18567 27121
rect 18509 27112 18521 27115
rect 18380 27084 18521 27112
rect 18380 27072 18386 27084
rect 18509 27081 18521 27084
rect 18555 27081 18567 27115
rect 18509 27075 18567 27081
rect 18598 27072 18604 27124
rect 18656 27112 18662 27124
rect 20622 27112 20628 27124
rect 18656 27084 20628 27112
rect 18656 27072 18662 27084
rect 20622 27072 20628 27084
rect 20680 27072 20686 27124
rect 20714 27072 20720 27124
rect 20772 27072 20778 27124
rect 22922 27072 22928 27124
rect 22980 27072 22986 27124
rect 23017 27115 23075 27121
rect 23017 27081 23029 27115
rect 23063 27112 23075 27115
rect 24305 27115 24363 27121
rect 24305 27112 24317 27115
rect 23063 27084 24317 27112
rect 23063 27081 23075 27084
rect 23017 27075 23075 27081
rect 24305 27081 24317 27084
rect 24351 27081 24363 27115
rect 24305 27075 24363 27081
rect 26510 27072 26516 27124
rect 26568 27112 26574 27124
rect 26621 27115 26679 27121
rect 26621 27112 26633 27115
rect 26568 27084 26633 27112
rect 26568 27072 26574 27084
rect 26621 27081 26633 27084
rect 26667 27081 26679 27115
rect 27154 27112 27160 27124
rect 26621 27075 26679 27081
rect 26988 27084 27160 27112
rect 12069 27047 12127 27053
rect 12069 27013 12081 27047
rect 12115 27044 12127 27047
rect 15378 27044 15384 27056
rect 12115 27016 13032 27044
rect 12115 27013 12127 27016
rect 12069 27007 12127 27013
rect 11849 26979 11907 26985
rect 11849 26945 11861 26979
rect 11895 26945 11907 26979
rect 11849 26939 11907 26945
rect 11974 26936 11980 26988
rect 12032 26936 12038 26988
rect 11606 26868 11612 26920
rect 11664 26908 11670 26920
rect 12084 26908 12112 27007
rect 13004 26988 13032 27016
rect 13096 27016 15384 27044
rect 12158 26936 12164 26988
rect 12216 26985 12222 26988
rect 12216 26976 12224 26985
rect 12216 26948 12261 26976
rect 12216 26939 12224 26948
rect 12216 26936 12222 26939
rect 12894 26936 12900 26988
rect 12952 26936 12958 26988
rect 12986 26936 12992 26988
rect 13044 26936 13050 26988
rect 11664 26880 12112 26908
rect 11664 26868 11670 26880
rect 12618 26868 12624 26920
rect 12676 26908 12682 26920
rect 13096 26908 13124 27016
rect 15378 27004 15384 27016
rect 15436 27044 15442 27056
rect 15657 27047 15715 27053
rect 15436 27016 15608 27044
rect 15436 27004 15442 27016
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14056 26948 14142 26976
rect 14056 26936 14062 26948
rect 12676 26880 13124 26908
rect 13173 26911 13231 26917
rect 12676 26868 12682 26880
rect 13173 26877 13185 26911
rect 13219 26908 13231 26911
rect 13630 26908 13636 26920
rect 13219 26880 13636 26908
rect 13219 26877 13231 26880
rect 13173 26871 13231 26877
rect 13630 26868 13636 26880
rect 13688 26908 13694 26920
rect 14114 26908 14142 26948
rect 14550 26936 14556 26988
rect 14608 26936 14614 26988
rect 15194 26976 15200 26988
rect 14660 26948 15200 26976
rect 14274 26908 14280 26920
rect 13688 26880 14044 26908
rect 14114 26880 14280 26908
rect 13688 26868 13694 26880
rect 14016 26849 14044 26880
rect 14274 26868 14280 26880
rect 14332 26908 14338 26920
rect 14660 26908 14688 26948
rect 15194 26936 15200 26948
rect 15252 26936 15258 26988
rect 15473 26979 15531 26985
rect 15473 26945 15485 26979
rect 15519 26945 15531 26979
rect 15473 26939 15531 26945
rect 14332 26880 14688 26908
rect 14332 26868 14338 26880
rect 14734 26868 14740 26920
rect 14792 26908 14798 26920
rect 14921 26911 14979 26917
rect 14921 26908 14933 26911
rect 14792 26880 14933 26908
rect 14792 26868 14798 26880
rect 14921 26877 14933 26880
rect 14967 26908 14979 26911
rect 15010 26908 15016 26920
rect 14967 26880 15016 26908
rect 14967 26877 14979 26880
rect 14921 26871 14979 26877
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 14001 26843 14059 26849
rect 14001 26809 14013 26843
rect 14047 26809 14059 26843
rect 15488 26840 15516 26939
rect 15580 26908 15608 27016
rect 15657 27013 15669 27047
rect 15703 27044 15715 27047
rect 16485 27047 16543 27053
rect 16485 27044 16497 27047
rect 15703 27016 16497 27044
rect 15703 27013 15715 27016
rect 15657 27007 15715 27013
rect 16485 27013 16497 27016
rect 16531 27013 16543 27047
rect 16485 27007 16543 27013
rect 15749 26979 15807 26985
rect 15749 26945 15761 26979
rect 15795 26976 15807 26979
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 15795 26948 16681 26976
rect 15795 26945 15807 26948
rect 15749 26939 15807 26945
rect 16669 26945 16681 26948
rect 16715 26976 16727 26979
rect 17144 26976 17172 27072
rect 17218 27004 17224 27056
rect 17276 27044 17282 27056
rect 19420 27047 19478 27053
rect 17276 27016 19196 27044
rect 17276 27004 17282 27016
rect 16715 26948 17172 26976
rect 16715 26945 16727 26948
rect 16669 26939 16727 26945
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 18414 26936 18420 26988
rect 18472 26936 18478 26988
rect 19168 26985 19196 27016
rect 19420 27013 19432 27047
rect 19466 27044 19478 27047
rect 20732 27044 20760 27072
rect 19466 27016 20760 27044
rect 22020 27016 22692 27044
rect 19466 27013 19478 27016
rect 19420 27007 19478 27013
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26945 19211 26979
rect 20346 26976 20352 26988
rect 19153 26939 19211 26945
rect 19260 26948 20352 26976
rect 15841 26911 15899 26917
rect 15841 26908 15853 26911
rect 15580 26880 15853 26908
rect 15841 26877 15853 26880
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 16945 26911 17003 26917
rect 16945 26908 16957 26911
rect 16816 26880 16957 26908
rect 16816 26868 16822 26880
rect 16945 26877 16957 26880
rect 16991 26877 17003 26911
rect 16945 26871 17003 26877
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 18598 26908 18604 26920
rect 17276 26880 18604 26908
rect 17276 26868 17282 26880
rect 18598 26868 18604 26880
rect 18656 26868 18662 26920
rect 19260 26908 19288 26948
rect 20346 26936 20352 26948
rect 20404 26936 20410 26988
rect 20898 26936 20904 26988
rect 20956 26976 20962 26988
rect 22020 26985 22048 27016
rect 22664 26988 22692 27016
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 20956 26948 22017 26976
rect 20956 26936 20962 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22094 26936 22100 26988
rect 22152 26936 22158 26988
rect 22278 26936 22284 26988
rect 22336 26936 22342 26988
rect 22646 26936 22652 26988
rect 22704 26936 22710 26988
rect 22741 26979 22799 26985
rect 22741 26945 22753 26979
rect 22787 26976 22799 26979
rect 22940 26976 22968 27072
rect 25133 27047 25191 27053
rect 22787 26948 22968 26976
rect 23308 27016 23612 27044
rect 22787 26945 22799 26948
rect 22741 26939 22799 26945
rect 23308 26920 23336 27016
rect 23385 26979 23443 26985
rect 23385 26945 23397 26979
rect 23431 26945 23443 26979
rect 23385 26939 23443 26945
rect 18708 26880 19288 26908
rect 16853 26843 16911 26849
rect 16853 26840 16865 26843
rect 15488 26812 16865 26840
rect 14001 26803 14059 26809
rect 16853 26809 16865 26812
rect 16899 26809 16911 26843
rect 16853 26803 16911 26809
rect 17678 26800 17684 26852
rect 17736 26840 17742 26852
rect 18708 26840 18736 26880
rect 20530 26868 20536 26920
rect 20588 26908 20594 26920
rect 20717 26911 20775 26917
rect 20717 26908 20729 26911
rect 20588 26880 20729 26908
rect 20588 26868 20594 26880
rect 20717 26877 20729 26880
rect 20763 26908 20775 26911
rect 20806 26908 20812 26920
rect 20763 26880 20812 26908
rect 20763 26877 20775 26880
rect 20717 26871 20775 26877
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 21174 26868 21180 26920
rect 21232 26908 21238 26920
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 21232 26880 22201 26908
rect 21232 26868 21238 26880
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 22189 26871 22247 26877
rect 23290 26868 23296 26920
rect 23348 26868 23354 26920
rect 21821 26843 21879 26849
rect 21821 26840 21833 26843
rect 17736 26812 18736 26840
rect 20079 26812 21833 26840
rect 17736 26800 17742 26812
rect 12989 26775 13047 26781
rect 12989 26772 13001 26775
rect 11440 26744 13001 26772
rect 12989 26741 13001 26744
rect 13035 26772 13047 26775
rect 13814 26772 13820 26784
rect 13035 26744 13820 26772
rect 13035 26741 13047 26744
rect 12989 26735 13047 26741
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 15102 26732 15108 26784
rect 15160 26772 15166 26784
rect 16761 26775 16819 26781
rect 16761 26772 16773 26775
rect 15160 26744 16773 26772
rect 15160 26732 15166 26744
rect 16761 26741 16773 26744
rect 16807 26741 16819 26775
rect 16761 26735 16819 26741
rect 17310 26732 17316 26784
rect 17368 26772 17374 26784
rect 17862 26772 17868 26784
rect 17368 26744 17868 26772
rect 17368 26732 17374 26744
rect 17862 26732 17868 26744
rect 17920 26732 17926 26784
rect 17954 26732 17960 26784
rect 18012 26732 18018 26784
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 19426 26772 19432 26784
rect 18840 26744 19432 26772
rect 18840 26732 18846 26744
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 19886 26732 19892 26784
rect 19944 26772 19950 26784
rect 20079 26772 20107 26812
rect 21821 26809 21833 26812
rect 21867 26809 21879 26843
rect 23400 26840 23428 26939
rect 23474 26936 23480 26988
rect 23532 26936 23538 26988
rect 23584 26917 23612 27016
rect 25133 27013 25145 27047
rect 25179 27044 25191 27047
rect 25222 27044 25228 27056
rect 25179 27016 25228 27044
rect 25179 27013 25191 27016
rect 25133 27007 25191 27013
rect 25222 27004 25228 27016
rect 25280 27044 25286 27056
rect 26237 27047 26295 27053
rect 26237 27044 26249 27047
rect 25280 27016 26249 27044
rect 25280 27004 25286 27016
rect 26237 27013 26249 27016
rect 26283 27013 26295 27047
rect 26237 27007 26295 27013
rect 26326 27004 26332 27056
rect 26384 27044 26390 27056
rect 26421 27047 26479 27053
rect 26421 27044 26433 27047
rect 26384 27016 26433 27044
rect 26384 27004 26390 27016
rect 26421 27013 26433 27016
rect 26467 27044 26479 27047
rect 26988 27044 27016 27084
rect 27154 27072 27160 27084
rect 27212 27072 27218 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 27982 27112 27988 27124
rect 27672 27084 27988 27112
rect 27672 27072 27678 27084
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 28074 27072 28080 27124
rect 28132 27112 28138 27124
rect 29454 27112 29460 27124
rect 28132 27084 29460 27112
rect 28132 27072 28138 27084
rect 29454 27072 29460 27084
rect 29512 27072 29518 27124
rect 30006 27072 30012 27124
rect 30064 27112 30070 27124
rect 30926 27112 30932 27124
rect 30064 27084 30932 27112
rect 30064 27072 30070 27084
rect 30926 27072 30932 27084
rect 30984 27072 30990 27124
rect 31110 27072 31116 27124
rect 31168 27112 31174 27124
rect 31941 27115 31999 27121
rect 31941 27112 31953 27115
rect 31168 27084 31953 27112
rect 31168 27072 31174 27084
rect 31941 27081 31953 27084
rect 31987 27081 31999 27115
rect 33505 27115 33563 27121
rect 33505 27112 33517 27115
rect 31941 27075 31999 27081
rect 32324 27084 33517 27112
rect 26467 27016 27016 27044
rect 27080 27016 28948 27044
rect 26467 27013 26479 27016
rect 26421 27007 26479 27013
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26976 24271 26979
rect 24946 26976 24952 26988
rect 24259 26948 24952 26976
rect 24259 26945 24271 26948
rect 24213 26939 24271 26945
rect 24946 26936 24952 26948
rect 25004 26936 25010 26988
rect 25038 26936 25044 26988
rect 25096 26936 25102 26988
rect 25682 26936 25688 26988
rect 25740 26936 25746 26988
rect 25866 26936 25872 26988
rect 25924 26936 25930 26988
rect 26142 26936 26148 26988
rect 26200 26976 26206 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 26200 26948 26985 26976
rect 26200 26936 26206 26948
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 26973 26939 27031 26945
rect 23569 26911 23627 26917
rect 23569 26877 23581 26911
rect 23615 26877 23627 26911
rect 23569 26871 23627 26877
rect 24394 26868 24400 26920
rect 24452 26868 24458 26920
rect 24486 26868 24492 26920
rect 24544 26908 24550 26920
rect 25225 26911 25283 26917
rect 24544 26880 25084 26908
rect 24544 26868 24550 26880
rect 24673 26843 24731 26849
rect 24673 26840 24685 26843
rect 23400 26812 24685 26840
rect 21821 26803 21879 26809
rect 24673 26809 24685 26812
rect 24719 26809 24731 26843
rect 25056 26840 25084 26880
rect 25225 26877 25237 26911
rect 25271 26877 25283 26911
rect 25225 26871 25283 26877
rect 25240 26840 25268 26871
rect 25314 26868 25320 26920
rect 25372 26908 25378 26920
rect 27080 26908 27108 27016
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26976 27215 26979
rect 27246 26976 27252 26988
rect 27203 26948 27252 26976
rect 27203 26945 27215 26948
rect 27157 26939 27215 26945
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27433 26979 27491 26985
rect 27433 26945 27445 26979
rect 27479 26976 27491 26979
rect 27614 26976 27620 26988
rect 27479 26948 27620 26976
rect 27479 26945 27491 26948
rect 27433 26939 27491 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 27709 26979 27767 26985
rect 27709 26945 27721 26979
rect 27755 26945 27767 26979
rect 27709 26939 27767 26945
rect 25372 26880 27108 26908
rect 25372 26868 25378 26880
rect 27338 26868 27344 26920
rect 27396 26908 27402 26920
rect 27724 26908 27752 26939
rect 27890 26936 27896 26988
rect 27948 26936 27954 26988
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 28350 26976 28356 26988
rect 28040 26948 28356 26976
rect 28040 26936 28046 26948
rect 28350 26936 28356 26948
rect 28408 26976 28414 26988
rect 28810 26985 28816 26988
rect 28629 26979 28687 26985
rect 28629 26976 28641 26979
rect 28408 26948 28641 26976
rect 28408 26936 28414 26948
rect 28629 26945 28641 26948
rect 28675 26945 28687 26979
rect 28807 26976 28816 26985
rect 28629 26939 28687 26945
rect 28736 26948 28816 26976
rect 28736 26908 28764 26948
rect 28807 26939 28816 26948
rect 28810 26936 28816 26939
rect 28868 26936 28874 26988
rect 27396 26880 27752 26908
rect 28281 26880 28764 26908
rect 28920 26908 28948 27016
rect 29840 27016 30788 27044
rect 29840 26985 29868 27016
rect 30760 26988 30788 27016
rect 31846 27004 31852 27056
rect 31904 27044 31910 27056
rect 32324 27044 32352 27084
rect 33505 27081 33517 27084
rect 33551 27081 33563 27115
rect 33505 27075 33563 27081
rect 33778 27072 33784 27124
rect 33836 27072 33842 27124
rect 34054 27072 34060 27124
rect 34112 27112 34118 27124
rect 34241 27115 34299 27121
rect 34241 27112 34253 27115
rect 34112 27084 34253 27112
rect 34112 27072 34118 27084
rect 34241 27081 34253 27084
rect 34287 27081 34299 27115
rect 34241 27075 34299 27081
rect 31904 27016 32352 27044
rect 32392 27047 32450 27053
rect 31904 27004 31910 27016
rect 32392 27013 32404 27047
rect 32438 27044 32450 27047
rect 33796 27044 33824 27072
rect 32438 27016 33824 27044
rect 32438 27013 32450 27016
rect 32392 27007 32450 27013
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 29825 26939 29883 26945
rect 30305 26969 30363 26975
rect 30305 26935 30317 26969
rect 30351 26966 30363 26969
rect 30351 26938 30420 26966
rect 30351 26935 30363 26938
rect 30305 26929 30363 26935
rect 29917 26911 29975 26917
rect 29917 26908 29929 26911
rect 28920 26880 29929 26908
rect 27396 26868 27402 26880
rect 26510 26840 26516 26852
rect 25056 26812 25268 26840
rect 25613 26812 26516 26840
rect 24673 26803 24731 26809
rect 19944 26744 20107 26772
rect 19944 26732 19950 26744
rect 20530 26732 20536 26784
rect 20588 26732 20594 26784
rect 20714 26732 20720 26784
rect 20772 26772 20778 26784
rect 21361 26775 21419 26781
rect 21361 26772 21373 26775
rect 20772 26744 21373 26772
rect 20772 26732 20778 26744
rect 21361 26741 21373 26744
rect 21407 26741 21419 26775
rect 21361 26735 21419 26741
rect 22186 26732 22192 26784
rect 22244 26772 22250 26784
rect 22833 26775 22891 26781
rect 22833 26772 22845 26775
rect 22244 26744 22845 26772
rect 22244 26732 22250 26744
rect 22833 26741 22845 26744
rect 22879 26741 22891 26775
rect 22833 26735 22891 26741
rect 23845 26775 23903 26781
rect 23845 26741 23857 26775
rect 23891 26772 23903 26775
rect 25613 26772 25641 26812
rect 26510 26800 26516 26812
rect 26568 26800 26574 26852
rect 27617 26843 27675 26849
rect 26620 26812 27568 26840
rect 23891 26744 25641 26772
rect 23891 26741 23903 26744
rect 23845 26735 23903 26741
rect 25682 26732 25688 26784
rect 25740 26732 25746 26784
rect 26620 26781 26648 26812
rect 26605 26775 26663 26781
rect 26605 26741 26617 26775
rect 26651 26741 26663 26775
rect 26605 26735 26663 26741
rect 26786 26732 26792 26784
rect 26844 26732 26850 26784
rect 26973 26775 27031 26781
rect 26973 26741 26985 26775
rect 27019 26772 27031 26775
rect 27430 26772 27436 26784
rect 27019 26744 27436 26772
rect 27019 26741 27031 26744
rect 26973 26735 27031 26741
rect 27430 26732 27436 26744
rect 27488 26732 27494 26784
rect 27540 26772 27568 26812
rect 27617 26809 27629 26843
rect 27663 26840 27675 26843
rect 28281 26840 28309 26880
rect 29917 26877 29929 26880
rect 29963 26877 29975 26911
rect 29917 26871 29975 26877
rect 30101 26911 30159 26917
rect 30101 26877 30113 26911
rect 30147 26908 30159 26911
rect 30190 26908 30196 26920
rect 30147 26880 30196 26908
rect 30147 26877 30159 26880
rect 30101 26871 30159 26877
rect 27663 26812 28309 26840
rect 27663 26809 27675 26812
rect 27617 26803 27675 26809
rect 28350 26800 28356 26852
rect 28408 26840 28414 26852
rect 28408 26812 28948 26840
rect 28408 26800 28414 26812
rect 28920 26784 28948 26812
rect 29730 26800 29736 26852
rect 29788 26840 29794 26852
rect 30116 26840 30144 26871
rect 30190 26868 30196 26880
rect 30248 26868 30254 26920
rect 30392 26908 30420 26938
rect 30742 26936 30748 26988
rect 30800 26936 30806 26988
rect 30834 26936 30840 26988
rect 30892 26936 30898 26988
rect 30926 26936 30932 26988
rect 30984 26936 30990 26988
rect 31018 26936 31024 26988
rect 31076 26936 31082 26988
rect 31202 26936 31208 26988
rect 31260 26936 31266 26988
rect 31294 26936 31300 26988
rect 31352 26936 31358 26988
rect 31938 26936 31944 26988
rect 31996 26936 32002 26988
rect 32122 26936 32128 26988
rect 32180 26936 32186 26988
rect 32214 26936 32220 26988
rect 32272 26976 32278 26988
rect 33781 26979 33839 26985
rect 33781 26976 33793 26979
rect 32272 26948 33793 26976
rect 32272 26936 32278 26948
rect 33781 26945 33793 26948
rect 33827 26945 33839 26979
rect 33781 26939 33839 26945
rect 31956 26908 31984 26936
rect 30392 26880 31984 26908
rect 33597 26911 33655 26917
rect 33597 26877 33609 26911
rect 33643 26908 33655 26911
rect 33870 26908 33876 26920
rect 33643 26880 33876 26908
rect 33643 26877 33655 26880
rect 33597 26871 33655 26877
rect 33870 26868 33876 26880
rect 33928 26908 33934 26920
rect 34072 26908 34100 27072
rect 33928 26880 34100 26908
rect 33928 26868 33934 26880
rect 29788 26812 30144 26840
rect 30469 26843 30527 26849
rect 29788 26800 29794 26812
rect 30469 26809 30481 26843
rect 30515 26840 30527 26843
rect 31846 26840 31852 26852
rect 30515 26812 31852 26840
rect 30515 26809 30527 26812
rect 30469 26803 30527 26809
rect 31846 26800 31852 26812
rect 31904 26800 31910 26852
rect 33965 26843 34023 26849
rect 33965 26840 33977 26843
rect 33060 26812 33977 26840
rect 27706 26772 27712 26784
rect 27540 26744 27712 26772
rect 27706 26732 27712 26744
rect 27764 26732 27770 26784
rect 28074 26732 28080 26784
rect 28132 26732 28138 26784
rect 28626 26732 28632 26784
rect 28684 26732 28690 26784
rect 28902 26732 28908 26784
rect 28960 26732 28966 26784
rect 29365 26775 29423 26781
rect 29365 26741 29377 26775
rect 29411 26772 29423 26775
rect 29454 26772 29460 26784
rect 29411 26744 29460 26772
rect 29411 26741 29423 26744
rect 29365 26735 29423 26741
rect 29454 26732 29460 26744
rect 29512 26772 29518 26784
rect 29822 26772 29828 26784
rect 29512 26744 29828 26772
rect 29512 26732 29518 26744
rect 29822 26732 29828 26744
rect 29880 26772 29886 26784
rect 30374 26772 30380 26784
rect 29880 26744 30380 26772
rect 29880 26732 29886 26744
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 30558 26732 30564 26784
rect 30616 26732 30622 26784
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 31478 26772 31484 26784
rect 30708 26744 31484 26772
rect 30708 26732 30714 26744
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 32030 26732 32036 26784
rect 32088 26772 32094 26784
rect 33060 26772 33088 26812
rect 33965 26809 33977 26812
rect 34011 26809 34023 26843
rect 33965 26803 34023 26809
rect 32088 26744 33088 26772
rect 32088 26732 32094 26744
rect 1104 26682 43884 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 43884 26682
rect 1104 26608 43884 26630
rect 4157 26571 4215 26577
rect 4157 26537 4169 26571
rect 4203 26568 4215 26571
rect 4798 26568 4804 26580
rect 4203 26540 4804 26568
rect 4203 26537 4215 26540
rect 4157 26531 4215 26537
rect 4798 26528 4804 26540
rect 4856 26568 4862 26580
rect 4856 26540 5212 26568
rect 4856 26528 4862 26540
rect 5184 26512 5212 26540
rect 5626 26528 5632 26580
rect 5684 26568 5690 26580
rect 6549 26571 6607 26577
rect 6549 26568 6561 26571
rect 5684 26540 6561 26568
rect 5684 26528 5690 26540
rect 6549 26537 6561 26540
rect 6595 26537 6607 26571
rect 6549 26531 6607 26537
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 7929 26571 7987 26577
rect 7929 26568 7941 26571
rect 7800 26540 7941 26568
rect 7800 26528 7806 26540
rect 7929 26537 7941 26540
rect 7975 26537 7987 26571
rect 7929 26531 7987 26537
rect 8202 26528 8208 26580
rect 8260 26568 8266 26580
rect 8941 26571 8999 26577
rect 8941 26568 8953 26571
rect 8260 26540 8953 26568
rect 8260 26528 8266 26540
rect 8941 26537 8953 26540
rect 8987 26537 8999 26571
rect 11238 26568 11244 26580
rect 8941 26531 8999 26537
rect 9048 26540 11244 26568
rect 1578 26460 1584 26512
rect 1636 26500 1642 26512
rect 4430 26500 4436 26512
rect 1636 26472 4436 26500
rect 1636 26460 1642 26472
rect 4430 26460 4436 26472
rect 4488 26460 4494 26512
rect 4525 26503 4583 26509
rect 4525 26469 4537 26503
rect 4571 26500 4583 26503
rect 4982 26500 4988 26512
rect 4571 26472 4988 26500
rect 4571 26469 4583 26472
rect 4525 26463 4583 26469
rect 4982 26460 4988 26472
rect 5040 26460 5046 26512
rect 5166 26460 5172 26512
rect 5224 26460 5230 26512
rect 5537 26503 5595 26509
rect 5537 26469 5549 26503
rect 5583 26469 5595 26503
rect 5537 26463 5595 26469
rect 4338 26392 4344 26444
rect 4396 26432 4402 26444
rect 4396 26404 5396 26432
rect 4396 26392 4402 26404
rect 1578 26324 1584 26376
rect 1636 26324 1642 26376
rect 3878 26324 3884 26376
rect 3936 26364 3942 26376
rect 4985 26367 5043 26373
rect 4985 26364 4997 26367
rect 3936 26336 4997 26364
rect 3936 26324 3942 26336
rect 4985 26333 4997 26336
rect 5031 26364 5043 26367
rect 5074 26364 5080 26376
rect 5031 26336 5080 26364
rect 5031 26333 5043 26336
rect 4985 26327 5043 26333
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 5166 26324 5172 26376
rect 5224 26324 5230 26376
rect 5368 26373 5396 26404
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26333 5411 26367
rect 5552 26364 5580 26463
rect 5902 26460 5908 26512
rect 5960 26500 5966 26512
rect 6454 26500 6460 26512
rect 5960 26472 6460 26500
rect 5960 26460 5966 26472
rect 6068 26373 6096 26472
rect 6454 26460 6460 26472
rect 6512 26460 6518 26512
rect 7558 26500 7564 26512
rect 6564 26472 7564 26500
rect 6564 26432 6592 26472
rect 7558 26460 7564 26472
rect 7616 26500 7622 26512
rect 9048 26500 9076 26540
rect 11238 26528 11244 26540
rect 11296 26528 11302 26580
rect 12986 26528 12992 26580
rect 13044 26568 13050 26580
rect 14829 26571 14887 26577
rect 14829 26568 14841 26571
rect 13044 26540 14841 26568
rect 13044 26528 13050 26540
rect 14829 26537 14841 26540
rect 14875 26568 14887 26571
rect 16114 26568 16120 26580
rect 14875 26540 16120 26568
rect 14875 26537 14887 26540
rect 14829 26531 14887 26537
rect 16114 26528 16120 26540
rect 16172 26568 16178 26580
rect 16209 26571 16267 26577
rect 16209 26568 16221 26571
rect 16172 26540 16221 26568
rect 16172 26528 16178 26540
rect 16209 26537 16221 26540
rect 16255 26537 16267 26571
rect 16209 26531 16267 26537
rect 17221 26571 17279 26577
rect 17221 26537 17233 26571
rect 17267 26568 17279 26571
rect 17678 26568 17684 26580
rect 17267 26540 17684 26568
rect 17267 26537 17279 26540
rect 17221 26531 17279 26537
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 17770 26528 17776 26580
rect 17828 26528 17834 26580
rect 17954 26528 17960 26580
rect 18012 26528 18018 26580
rect 18490 26571 18548 26577
rect 18490 26537 18502 26571
rect 18536 26568 18548 26571
rect 19613 26571 19671 26577
rect 18536 26540 19196 26568
rect 18536 26537 18548 26540
rect 18490 26531 18548 26537
rect 7616 26472 9076 26500
rect 9401 26503 9459 26509
rect 7616 26460 7622 26472
rect 9401 26469 9413 26503
rect 9447 26500 9459 26503
rect 15013 26503 15071 26509
rect 9447 26472 14780 26500
rect 9447 26469 9459 26472
rect 9401 26463 9459 26469
rect 6196 26404 6592 26432
rect 7213 26404 7834 26432
rect 6196 26373 6224 26404
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5552 26336 5917 26364
rect 5353 26327 5411 26333
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6053 26367 6111 26373
rect 6053 26333 6065 26367
rect 6099 26333 6111 26367
rect 6053 26327 6111 26333
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 2593 26299 2651 26305
rect 2593 26265 2605 26299
rect 2639 26296 2651 26299
rect 2774 26296 2780 26308
rect 2639 26268 2780 26296
rect 2639 26265 2651 26268
rect 2593 26259 2651 26265
rect 2774 26256 2780 26268
rect 2832 26256 2838 26308
rect 3237 26299 3295 26305
rect 3237 26265 3249 26299
rect 3283 26296 3295 26299
rect 3786 26296 3792 26308
rect 3283 26268 3792 26296
rect 3283 26265 3295 26268
rect 3237 26259 3295 26265
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 3970 26256 3976 26308
rect 4028 26296 4034 26308
rect 5261 26299 5319 26305
rect 5261 26296 5273 26299
rect 4028 26268 5273 26296
rect 4028 26256 4034 26268
rect 5261 26265 5273 26268
rect 5307 26265 5319 26299
rect 5368 26296 5396 26327
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 6411 26367 6469 26373
rect 6411 26333 6423 26367
rect 6457 26364 6469 26367
rect 6822 26364 6828 26376
rect 6457 26336 6828 26364
rect 6457 26333 6469 26336
rect 6411 26327 6469 26333
rect 6822 26324 6828 26336
rect 6880 26364 6886 26376
rect 7213 26364 7241 26404
rect 6880 26336 7241 26364
rect 6880 26324 6886 26336
rect 7282 26324 7288 26376
rect 7340 26324 7346 26376
rect 7374 26324 7380 26376
rect 7432 26364 7438 26376
rect 7806 26373 7834 26404
rect 8294 26392 8300 26444
rect 8352 26392 8358 26444
rect 8386 26392 8392 26444
rect 8444 26432 8450 26444
rect 8444 26404 9674 26432
rect 8444 26392 8450 26404
rect 7791 26367 7849 26373
rect 7432 26336 7477 26364
rect 7432 26324 7438 26336
rect 7791 26333 7803 26367
rect 7837 26364 7849 26367
rect 8202 26364 8208 26376
rect 7837 26336 8208 26364
rect 7837 26333 7849 26336
rect 7791 26327 7849 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8312 26336 9137 26364
rect 5626 26296 5632 26308
rect 5368 26268 5632 26296
rect 5261 26259 5319 26265
rect 5626 26256 5632 26268
rect 5684 26296 5690 26308
rect 5684 26268 6960 26296
rect 5684 26256 5690 26268
rect 6012 26240 6040 26268
rect 3605 26231 3663 26237
rect 3605 26197 3617 26231
rect 3651 26228 3663 26231
rect 3694 26228 3700 26240
rect 3651 26200 3700 26228
rect 3651 26197 3663 26200
rect 3605 26191 3663 26197
rect 3694 26188 3700 26200
rect 3752 26188 3758 26240
rect 4893 26231 4951 26237
rect 4893 26197 4905 26231
rect 4939 26228 4951 26231
rect 5166 26228 5172 26240
rect 4939 26200 5172 26228
rect 4939 26197 4951 26200
rect 4893 26191 4951 26197
rect 5166 26188 5172 26200
rect 5224 26188 5230 26240
rect 5534 26188 5540 26240
rect 5592 26228 5598 26240
rect 5810 26228 5816 26240
rect 5592 26200 5816 26228
rect 5592 26188 5598 26200
rect 5810 26188 5816 26200
rect 5868 26188 5874 26240
rect 5994 26188 6000 26240
rect 6052 26188 6058 26240
rect 6932 26237 6960 26268
rect 7558 26256 7564 26308
rect 7616 26256 7622 26308
rect 7653 26299 7711 26305
rect 7653 26265 7665 26299
rect 7699 26296 7711 26299
rect 8110 26296 8116 26308
rect 7699 26268 8116 26296
rect 7699 26265 7711 26268
rect 7653 26259 7711 26265
rect 8110 26256 8116 26268
rect 8168 26296 8174 26308
rect 8312 26296 8340 26336
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 9398 26324 9404 26376
rect 9456 26324 9462 26376
rect 8168 26268 8340 26296
rect 8665 26299 8723 26305
rect 8168 26256 8174 26268
rect 8665 26265 8677 26299
rect 8711 26296 8723 26299
rect 8846 26296 8852 26308
rect 8711 26268 8852 26296
rect 8711 26265 8723 26268
rect 8665 26259 8723 26265
rect 8846 26256 8852 26268
rect 8904 26256 8910 26308
rect 8941 26299 8999 26305
rect 8941 26265 8953 26299
rect 8987 26296 8999 26299
rect 9030 26296 9036 26308
rect 8987 26268 9036 26296
rect 8987 26265 8999 26268
rect 8941 26259 8999 26265
rect 9030 26256 9036 26268
rect 9088 26296 9094 26308
rect 9416 26296 9444 26324
rect 9088 26268 9444 26296
rect 9646 26296 9674 26404
rect 10594 26392 10600 26444
rect 10652 26432 10658 26444
rect 10870 26432 10876 26444
rect 10652 26404 10876 26432
rect 10652 26392 10658 26404
rect 10870 26392 10876 26404
rect 10928 26432 10934 26444
rect 11146 26432 11152 26444
rect 10928 26404 11152 26432
rect 10928 26392 10934 26404
rect 11146 26392 11152 26404
rect 11204 26392 11210 26444
rect 11238 26392 11244 26444
rect 11296 26432 11302 26444
rect 11514 26432 11520 26444
rect 11296 26404 11520 26432
rect 11296 26392 11302 26404
rect 11514 26392 11520 26404
rect 11572 26392 11578 26444
rect 13998 26432 14004 26444
rect 13464 26404 14004 26432
rect 10962 26324 10968 26376
rect 11020 26364 11026 26376
rect 11609 26367 11667 26373
rect 11609 26364 11621 26367
rect 11020 26336 11621 26364
rect 11020 26324 11026 26336
rect 11609 26333 11621 26336
rect 11655 26364 11667 26367
rect 11790 26364 11796 26376
rect 11655 26336 11796 26364
rect 11655 26333 11667 26336
rect 11609 26327 11667 26333
rect 11790 26324 11796 26336
rect 11848 26364 11854 26376
rect 12526 26364 12532 26376
rect 11848 26336 12532 26364
rect 11848 26324 11854 26336
rect 12526 26324 12532 26336
rect 12584 26324 12590 26376
rect 13464 26373 13492 26404
rect 13998 26392 14004 26404
rect 14056 26392 14062 26444
rect 14366 26392 14372 26444
rect 14424 26432 14430 26444
rect 14645 26435 14703 26441
rect 14645 26432 14657 26435
rect 14424 26404 14657 26432
rect 14424 26392 14430 26404
rect 14645 26401 14657 26404
rect 14691 26401 14703 26435
rect 14752 26432 14780 26472
rect 15013 26469 15025 26503
rect 15059 26500 15071 26503
rect 15381 26503 15439 26509
rect 15381 26500 15393 26503
rect 15059 26472 15393 26500
rect 15059 26469 15071 26472
rect 15013 26463 15071 26469
rect 15381 26469 15393 26472
rect 15427 26469 15439 26503
rect 15381 26463 15439 26469
rect 15746 26460 15752 26512
rect 15804 26500 15810 26512
rect 16942 26500 16948 26512
rect 15804 26472 16948 26500
rect 15804 26460 15810 26472
rect 15473 26435 15531 26441
rect 15473 26432 15485 26435
rect 14752 26404 15485 26432
rect 14645 26395 14703 26401
rect 15473 26401 15485 26404
rect 15519 26401 15531 26435
rect 15473 26395 15531 26401
rect 15565 26435 15623 26441
rect 15565 26401 15577 26435
rect 15611 26432 15623 26435
rect 15654 26432 15660 26444
rect 15611 26404 15660 26432
rect 15611 26401 15623 26404
rect 15565 26395 15623 26401
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 13603 26367 13661 26373
rect 13603 26333 13615 26367
rect 13649 26364 13661 26367
rect 13722 26364 13728 26376
rect 13649 26336 13728 26364
rect 13649 26333 13661 26336
rect 13603 26327 13661 26333
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 13814 26324 13820 26376
rect 13872 26324 13878 26376
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 13924 26336 14841 26364
rect 12342 26296 12348 26308
rect 9646 26268 12348 26296
rect 9088 26256 9094 26268
rect 12342 26256 12348 26268
rect 12400 26256 12406 26308
rect 12434 26256 12440 26308
rect 12492 26296 12498 26308
rect 13357 26299 13415 26305
rect 13357 26296 13369 26299
rect 12492 26268 13369 26296
rect 12492 26256 12498 26268
rect 13357 26265 13369 26268
rect 13403 26296 13415 26299
rect 13924 26296 13952 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 13403 26268 13952 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 14550 26256 14556 26308
rect 14608 26256 14614 26308
rect 14844 26296 14872 26327
rect 15286 26324 15292 26376
rect 15344 26324 15350 26376
rect 15378 26324 15384 26376
rect 15436 26364 15442 26376
rect 15580 26364 15608 26395
rect 15654 26392 15660 26404
rect 15712 26392 15718 26444
rect 15856 26441 15884 26472
rect 16942 26460 16948 26472
rect 17000 26460 17006 26512
rect 17788 26500 17816 26528
rect 17604 26472 17816 26500
rect 15841 26435 15899 26441
rect 15841 26401 15853 26435
rect 15887 26401 15899 26435
rect 15841 26395 15899 26401
rect 16132 26404 17549 26432
rect 15436 26336 15608 26364
rect 15749 26367 15807 26373
rect 15436 26324 15442 26336
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 15930 26364 15936 26376
rect 15795 26336 15936 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16132 26296 16160 26404
rect 16390 26324 16396 26376
rect 16448 26324 16454 26376
rect 16482 26324 16488 26376
rect 16540 26364 16546 26376
rect 16666 26364 16672 26376
rect 16540 26336 16672 26364
rect 16540 26324 16546 26336
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 16758 26324 16764 26376
rect 16816 26364 16822 26376
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 16816 26336 17417 26364
rect 16816 26324 16822 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 16408 26296 16436 26324
rect 14844 26268 16160 26296
rect 16224 26268 16436 26296
rect 6917 26231 6975 26237
rect 6917 26197 6929 26231
rect 6963 26228 6975 26231
rect 7098 26228 7104 26240
rect 6963 26200 7104 26228
rect 6963 26197 6975 26200
rect 6917 26191 6975 26197
rect 7098 26188 7104 26200
rect 7156 26228 7162 26240
rect 7742 26228 7748 26240
rect 7156 26200 7748 26228
rect 7156 26188 7162 26200
rect 7742 26188 7748 26200
rect 7800 26228 7806 26240
rect 10318 26228 10324 26240
rect 7800 26200 10324 26228
rect 7800 26188 7806 26200
rect 10318 26188 10324 26200
rect 10376 26188 10382 26240
rect 10502 26188 10508 26240
rect 10560 26228 10566 26240
rect 11054 26228 11060 26240
rect 10560 26200 11060 26228
rect 10560 26188 10566 26200
rect 11054 26188 11060 26200
rect 11112 26228 11118 26240
rect 12452 26228 12480 26256
rect 11112 26200 12480 26228
rect 14369 26231 14427 26237
rect 11112 26188 11118 26200
rect 14369 26197 14381 26231
rect 14415 26228 14427 26231
rect 14458 26228 14464 26240
rect 14415 26200 14464 26228
rect 14415 26197 14427 26200
rect 14369 26191 14427 26197
rect 14458 26188 14464 26200
rect 14516 26188 14522 26240
rect 15102 26188 15108 26240
rect 15160 26188 15166 26240
rect 15838 26188 15844 26240
rect 15896 26228 15902 26240
rect 16224 26237 16252 26268
rect 16942 26256 16948 26308
rect 17000 26256 17006 26308
rect 17129 26299 17187 26305
rect 17129 26265 17141 26299
rect 17175 26296 17187 26299
rect 17310 26296 17316 26308
rect 17175 26268 17316 26296
rect 17175 26265 17187 26268
rect 17129 26259 17187 26265
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 17521 26296 17549 26404
rect 17604 26373 17632 26472
rect 17972 26432 18000 26528
rect 18601 26503 18659 26509
rect 18601 26469 18613 26503
rect 18647 26500 18659 26503
rect 18782 26500 18788 26512
rect 18647 26472 18788 26500
rect 18647 26469 18659 26472
rect 18601 26463 18659 26469
rect 18782 26460 18788 26472
rect 18840 26460 18846 26512
rect 19168 26444 19196 26540
rect 19613 26537 19625 26571
rect 19659 26568 19671 26571
rect 20070 26568 20076 26580
rect 19659 26540 20076 26568
rect 19659 26537 19671 26540
rect 19613 26531 19671 26537
rect 20070 26528 20076 26540
rect 20128 26528 20134 26580
rect 20622 26528 20628 26580
rect 20680 26568 20686 26580
rect 21361 26571 21419 26577
rect 20680 26540 20852 26568
rect 20680 26528 20686 26540
rect 20824 26512 20852 26540
rect 21361 26537 21373 26571
rect 21407 26568 21419 26571
rect 22278 26568 22284 26580
rect 21407 26540 22284 26568
rect 21407 26537 21419 26540
rect 21361 26531 21419 26537
rect 22278 26528 22284 26540
rect 22336 26528 22342 26580
rect 23474 26528 23480 26580
rect 23532 26528 23538 26580
rect 23750 26528 23756 26580
rect 23808 26528 23814 26580
rect 24213 26571 24271 26577
rect 24213 26537 24225 26571
rect 24259 26568 24271 26571
rect 24578 26568 24584 26580
rect 24259 26540 24584 26568
rect 24259 26537 24271 26540
rect 24213 26531 24271 26537
rect 24578 26528 24584 26540
rect 24636 26528 24642 26580
rect 25038 26528 25044 26580
rect 25096 26568 25102 26580
rect 25133 26571 25191 26577
rect 25133 26568 25145 26571
rect 25096 26540 25145 26568
rect 25096 26528 25102 26540
rect 25133 26537 25145 26540
rect 25179 26537 25191 26571
rect 25133 26531 25191 26537
rect 25685 26571 25743 26577
rect 25685 26537 25697 26571
rect 25731 26568 25743 26571
rect 25866 26568 25872 26580
rect 25731 26540 25872 26568
rect 25731 26537 25743 26540
rect 25685 26531 25743 26537
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 26050 26528 26056 26580
rect 26108 26528 26114 26580
rect 26234 26528 26240 26580
rect 26292 26528 26298 26580
rect 26878 26528 26884 26580
rect 26936 26528 26942 26580
rect 27614 26528 27620 26580
rect 27672 26568 27678 26580
rect 28077 26571 28135 26577
rect 28077 26568 28089 26571
rect 27672 26540 28089 26568
rect 27672 26528 27678 26540
rect 28077 26537 28089 26540
rect 28123 26537 28135 26571
rect 28077 26531 28135 26537
rect 28442 26528 28448 26580
rect 28500 26528 28506 26580
rect 28813 26571 28871 26577
rect 28813 26568 28825 26571
rect 28644 26540 28825 26568
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 20864 26472 22692 26500
rect 20864 26460 20870 26472
rect 17696 26404 18000 26432
rect 18156 26404 18368 26432
rect 17696 26373 17724 26404
rect 17589 26367 17647 26373
rect 17589 26333 17601 26367
rect 17635 26333 17647 26367
rect 17589 26327 17647 26333
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 17770 26324 17776 26376
rect 17828 26324 17834 26376
rect 18156 26364 18184 26404
rect 17880 26336 18184 26364
rect 17880 26296 17908 26336
rect 18230 26324 18236 26376
rect 18288 26324 18294 26376
rect 18340 26364 18368 26404
rect 18414 26392 18420 26444
rect 18472 26432 18478 26444
rect 18693 26435 18751 26441
rect 18693 26432 18705 26435
rect 18472 26404 18705 26432
rect 18472 26392 18478 26404
rect 18693 26401 18705 26404
rect 18739 26401 18751 26435
rect 18693 26395 18751 26401
rect 18874 26392 18880 26444
rect 18932 26392 18938 26444
rect 19150 26392 19156 26444
rect 19208 26392 19214 26444
rect 20993 26435 21051 26441
rect 20993 26432 21005 26435
rect 19694 26404 21005 26432
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 18340 26336 19441 26364
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 18248 26296 18276 26324
rect 17521 26268 17908 26296
rect 17972 26268 18276 26296
rect 18325 26299 18383 26305
rect 16209 26231 16267 26237
rect 16209 26228 16221 26231
rect 15896 26200 16221 26228
rect 15896 26188 15902 26200
rect 16209 26197 16221 26200
rect 16255 26197 16267 26231
rect 16209 26191 16267 26197
rect 16390 26188 16396 26240
rect 16448 26188 16454 26240
rect 16666 26188 16672 26240
rect 16724 26188 16730 26240
rect 16960 26228 16988 26256
rect 17218 26228 17224 26240
rect 16960 26200 17224 26228
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 17972 26237 18000 26268
rect 18325 26265 18337 26299
rect 18371 26296 18383 26299
rect 19444 26296 19472 26327
rect 19694 26296 19722 26404
rect 20993 26401 21005 26404
rect 21039 26401 21051 26435
rect 20993 26395 21051 26401
rect 21174 26392 21180 26444
rect 21232 26392 21238 26444
rect 21358 26392 21364 26444
rect 21416 26432 21422 26444
rect 21637 26435 21695 26441
rect 21637 26432 21649 26435
rect 21416 26404 21649 26432
rect 21416 26392 21422 26404
rect 21637 26401 21649 26404
rect 21683 26401 21695 26435
rect 21637 26395 21695 26401
rect 21726 26392 21732 26444
rect 21784 26392 21790 26444
rect 22664 26376 22692 26472
rect 23768 26432 23796 26528
rect 26068 26500 26096 26528
rect 24596 26472 26096 26500
rect 26896 26500 26924 26528
rect 28460 26500 28488 26528
rect 26896 26472 27476 26500
rect 24596 26441 24624 26472
rect 24581 26435 24639 26441
rect 23768 26404 23888 26432
rect 19869 26367 19927 26373
rect 19869 26333 19881 26367
rect 19915 26333 19927 26367
rect 19869 26327 19927 26333
rect 18371 26268 19334 26296
rect 19444 26268 19722 26296
rect 19895 26296 19923 26327
rect 19959 26324 19965 26376
rect 20017 26324 20023 26376
rect 20070 26324 20076 26376
rect 20128 26324 20134 26376
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20346 26364 20352 26376
rect 20303 26336 20352 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 20622 26324 20628 26376
rect 20680 26364 20686 26376
rect 21542 26364 21548 26376
rect 20680 26336 21548 26364
rect 20680 26324 20686 26336
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 20714 26296 20720 26308
rect 19895 26268 20720 26296
rect 18371 26265 18383 26268
rect 18325 26259 18383 26265
rect 17957 26231 18015 26237
rect 17957 26197 17969 26231
rect 18003 26197 18015 26231
rect 19306 26228 19334 26268
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 20990 26256 20996 26308
rect 21048 26296 21054 26308
rect 21836 26296 21864 26327
rect 22002 26324 22008 26376
rect 22060 26324 22066 26376
rect 22646 26324 22652 26376
rect 22704 26364 22710 26376
rect 23290 26364 23296 26376
rect 22704 26336 23296 26364
rect 22704 26324 22710 26336
rect 23290 26324 23296 26336
rect 23348 26364 23354 26376
rect 23750 26373 23756 26376
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 23348 26336 23581 26364
rect 23348 26324 23354 26336
rect 23569 26333 23581 26336
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23717 26367 23756 26373
rect 23717 26333 23729 26367
rect 23717 26327 23756 26333
rect 23750 26324 23756 26327
rect 23808 26324 23814 26376
rect 23860 26364 23888 26404
rect 24581 26401 24593 26435
rect 24627 26401 24639 26435
rect 24581 26395 24639 26401
rect 24034 26367 24092 26373
rect 24034 26364 24046 26367
rect 23860 26336 24046 26364
rect 24034 26333 24046 26336
rect 24080 26333 24092 26367
rect 24596 26364 24624 26395
rect 25406 26392 25412 26444
rect 25464 26392 25470 26444
rect 25498 26392 25504 26444
rect 25556 26432 25562 26444
rect 25556 26404 25913 26432
rect 25556 26392 25562 26404
rect 24034 26327 24092 26333
rect 24136 26336 24624 26364
rect 24765 26367 24823 26373
rect 21048 26268 22416 26296
rect 21048 26256 21054 26268
rect 20438 26228 20444 26240
rect 19306 26200 20444 26228
rect 17957 26191 18015 26197
rect 20438 26188 20444 26200
rect 20496 26188 20502 26240
rect 20530 26188 20536 26240
rect 20588 26188 20594 26240
rect 20901 26231 20959 26237
rect 20901 26197 20913 26231
rect 20947 26228 20959 26231
rect 21082 26228 21088 26240
rect 20947 26200 21088 26228
rect 20947 26197 20959 26200
rect 20901 26191 20959 26197
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 22388 26237 22416 26268
rect 23474 26256 23480 26308
rect 23532 26296 23538 26308
rect 23845 26299 23903 26305
rect 23845 26296 23857 26299
rect 23532 26268 23857 26296
rect 23532 26256 23538 26268
rect 23845 26265 23857 26268
rect 23891 26265 23903 26299
rect 23845 26259 23903 26265
rect 23934 26256 23940 26308
rect 23992 26256 23998 26308
rect 22373 26231 22431 26237
rect 22373 26197 22385 26231
rect 22419 26228 22431 26231
rect 24136 26228 24164 26336
rect 24765 26333 24777 26367
rect 24811 26364 24823 26367
rect 25314 26364 25320 26376
rect 24811 26336 25320 26364
rect 24811 26333 24823 26336
rect 24765 26327 24823 26333
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 25424 26364 25452 26392
rect 25593 26367 25651 26373
rect 25593 26364 25605 26367
rect 25424 26336 25605 26364
rect 25593 26333 25605 26336
rect 25639 26333 25651 26367
rect 25593 26327 25651 26333
rect 25774 26324 25780 26376
rect 25832 26324 25838 26376
rect 24302 26256 24308 26308
rect 24360 26296 24366 26308
rect 24673 26299 24731 26305
rect 24673 26296 24685 26299
rect 24360 26268 24685 26296
rect 24360 26256 24366 26268
rect 24673 26265 24685 26268
rect 24719 26296 24731 26299
rect 25409 26299 25467 26305
rect 25409 26296 25421 26299
rect 24719 26268 25421 26296
rect 24719 26265 24731 26268
rect 24673 26259 24731 26265
rect 25409 26265 25421 26268
rect 25455 26265 25467 26299
rect 25885 26296 25913 26404
rect 25958 26392 25964 26444
rect 26016 26432 26022 26444
rect 26605 26435 26663 26441
rect 26881 26440 26939 26441
rect 26605 26432 26617 26435
rect 26016 26404 26617 26432
rect 26016 26392 26022 26404
rect 26605 26401 26617 26404
rect 26651 26401 26663 26435
rect 26605 26395 26663 26401
rect 26817 26435 26939 26440
rect 26817 26412 26893 26435
rect 26142 26324 26148 26376
rect 26200 26324 26206 26376
rect 26237 26367 26295 26373
rect 26237 26333 26249 26367
rect 26283 26333 26295 26367
rect 26237 26327 26295 26333
rect 26252 26296 26280 26327
rect 26418 26324 26424 26376
rect 26476 26364 26482 26376
rect 26817 26364 26845 26412
rect 26881 26401 26893 26412
rect 26927 26401 26939 26435
rect 26881 26395 26939 26401
rect 27090 26435 27148 26441
rect 27341 26440 27399 26441
rect 27090 26401 27102 26435
rect 27136 26432 27148 26435
rect 27264 26435 27399 26440
rect 27264 26432 27353 26435
rect 27136 26412 27353 26432
rect 27136 26404 27292 26412
rect 27136 26401 27148 26404
rect 27090 26395 27148 26401
rect 27341 26401 27353 26412
rect 27387 26401 27399 26435
rect 27341 26395 27399 26401
rect 26476 26336 26845 26364
rect 26988 26361 27109 26364
rect 27246 26361 27252 26376
rect 26988 26336 27252 26361
rect 26476 26324 26482 26336
rect 26988 26296 27016 26336
rect 27081 26333 27252 26336
rect 27246 26324 27252 26333
rect 27304 26324 27310 26376
rect 25885 26268 27016 26296
rect 27448 26296 27476 26472
rect 27540 26472 28488 26500
rect 27540 26373 27568 26472
rect 27614 26392 27620 26444
rect 27672 26392 27678 26444
rect 28169 26435 28227 26441
rect 28169 26432 28181 26435
rect 27724 26404 28181 26432
rect 27724 26373 27752 26404
rect 28169 26401 28181 26404
rect 28215 26401 28227 26435
rect 28169 26395 28227 26401
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 27709 26367 27767 26373
rect 27801 26370 27859 26373
rect 27709 26333 27721 26367
rect 27755 26333 27767 26367
rect 27709 26327 27767 26333
rect 27724 26296 27752 26327
rect 27798 26318 27804 26370
rect 27856 26358 27862 26370
rect 27985 26367 28043 26373
rect 27856 26330 27895 26358
rect 27985 26333 27997 26367
rect 28031 26333 28043 26367
rect 27856 26318 27862 26330
rect 27985 26327 28043 26333
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26364 28411 26367
rect 28460 26364 28488 26472
rect 28644 26432 28672 26540
rect 28813 26537 28825 26540
rect 28859 26537 28871 26571
rect 28813 26531 28871 26537
rect 28902 26528 28908 26580
rect 28960 26568 28966 26580
rect 29181 26571 29239 26577
rect 29181 26568 29193 26571
rect 28960 26540 29193 26568
rect 28960 26528 28966 26540
rect 29181 26537 29193 26540
rect 29227 26537 29239 26571
rect 29181 26531 29239 26537
rect 29840 26540 30052 26568
rect 28718 26460 28724 26512
rect 28776 26500 28782 26512
rect 29840 26500 29868 26540
rect 28776 26472 29868 26500
rect 30024 26500 30052 26540
rect 30742 26528 30748 26580
rect 30800 26568 30806 26580
rect 31110 26568 31116 26580
rect 30800 26540 31116 26568
rect 30800 26528 30806 26540
rect 31110 26528 31116 26540
rect 31168 26528 31174 26580
rect 31294 26528 31300 26580
rect 31352 26568 31358 26580
rect 33137 26571 33195 26577
rect 33137 26568 33149 26571
rect 31352 26540 33149 26568
rect 31352 26528 31358 26540
rect 33137 26537 33149 26540
rect 33183 26537 33195 26571
rect 33137 26531 33195 26537
rect 33870 26528 33876 26580
rect 33928 26528 33934 26580
rect 30929 26503 30987 26509
rect 30929 26500 30941 26503
rect 30024 26472 30941 26500
rect 28776 26460 28782 26472
rect 30929 26469 30941 26472
rect 30975 26469 30987 26503
rect 30929 26463 30987 26469
rect 32766 26460 32772 26512
rect 32824 26500 32830 26512
rect 33413 26503 33471 26509
rect 33413 26500 33425 26503
rect 32824 26472 33425 26500
rect 32824 26460 32830 26472
rect 33413 26469 33425 26472
rect 33459 26469 33471 26503
rect 33413 26463 33471 26469
rect 28902 26432 28908 26444
rect 28644 26404 28908 26432
rect 28902 26392 28908 26404
rect 28960 26392 28966 26444
rect 29365 26435 29423 26441
rect 29365 26401 29377 26435
rect 29411 26432 29423 26435
rect 29546 26432 29552 26444
rect 29411 26404 29552 26432
rect 29411 26401 29423 26404
rect 29365 26395 29423 26401
rect 29546 26392 29552 26404
rect 29604 26432 29610 26444
rect 29604 26404 29960 26432
rect 29604 26392 29610 26404
rect 29932 26376 29960 26404
rect 30374 26392 30380 26444
rect 30432 26432 30438 26444
rect 30432 26404 31432 26432
rect 30432 26392 30438 26404
rect 29089 26367 29147 26373
rect 29089 26364 29101 26367
rect 28399 26336 29101 26364
rect 28399 26333 28411 26336
rect 28353 26327 28411 26333
rect 29089 26333 29101 26336
rect 29135 26333 29147 26367
rect 29089 26327 29147 26333
rect 29564 26336 29776 26364
rect 27448 26268 27752 26296
rect 25409 26259 25467 26265
rect 28000 26240 28028 26327
rect 28077 26299 28135 26305
rect 28077 26265 28089 26299
rect 28123 26296 28135 26299
rect 28442 26296 28448 26308
rect 28123 26268 28448 26296
rect 28123 26265 28135 26268
rect 28077 26259 28135 26265
rect 28442 26256 28448 26268
rect 28500 26256 28506 26308
rect 28629 26299 28687 26305
rect 28629 26265 28641 26299
rect 28675 26296 28687 26299
rect 28829 26299 28887 26305
rect 28675 26268 28764 26296
rect 28675 26265 28687 26268
rect 28629 26259 28687 26265
rect 28736 26240 28764 26268
rect 28829 26265 28841 26299
rect 28875 26296 28887 26299
rect 29365 26299 29423 26305
rect 28875 26268 29132 26296
rect 28875 26265 28887 26268
rect 28829 26259 28887 26265
rect 29104 26240 29132 26268
rect 29365 26265 29377 26299
rect 29411 26296 29423 26299
rect 29564 26296 29592 26336
rect 29411 26268 29592 26296
rect 29411 26265 29423 26268
rect 29365 26259 29423 26265
rect 22419 26200 24164 26228
rect 22419 26197 22431 26200
rect 22373 26191 22431 26197
rect 26418 26188 26424 26240
rect 26476 26228 26482 26240
rect 26513 26231 26571 26237
rect 26513 26228 26525 26231
rect 26476 26200 26525 26228
rect 26476 26188 26482 26200
rect 26513 26197 26525 26200
rect 26559 26197 26571 26231
rect 26513 26191 26571 26197
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 26973 26231 27031 26237
rect 26973 26228 26985 26231
rect 26844 26200 26985 26228
rect 26844 26188 26850 26200
rect 26973 26197 26985 26200
rect 27019 26197 27031 26231
rect 26973 26191 27031 26197
rect 27246 26188 27252 26240
rect 27304 26188 27310 26240
rect 27982 26188 27988 26240
rect 28040 26188 28046 26240
rect 28534 26188 28540 26240
rect 28592 26188 28598 26240
rect 28718 26188 28724 26240
rect 28776 26188 28782 26240
rect 28994 26188 29000 26240
rect 29052 26188 29058 26240
rect 29086 26188 29092 26240
rect 29144 26188 29150 26240
rect 29546 26188 29552 26240
rect 29604 26188 29610 26240
rect 29748 26228 29776 26336
rect 29822 26324 29828 26376
rect 29880 26324 29886 26376
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 30009 26367 30067 26373
rect 30009 26333 30021 26367
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 30024 26228 30052 26327
rect 30190 26324 30196 26376
rect 30248 26364 30254 26376
rect 30248 26336 30604 26364
rect 30248 26324 30254 26336
rect 30282 26256 30288 26308
rect 30340 26256 30346 26308
rect 30576 26296 30604 26336
rect 30650 26324 30656 26376
rect 30708 26324 30714 26376
rect 30760 26373 30788 26404
rect 30745 26367 30803 26373
rect 30745 26333 30757 26367
rect 30791 26333 30803 26367
rect 30745 26327 30803 26333
rect 30926 26324 30932 26376
rect 30984 26364 30990 26376
rect 31113 26367 31171 26373
rect 31113 26364 31125 26367
rect 30984 26336 31125 26364
rect 30984 26324 30990 26336
rect 31113 26333 31125 26336
rect 31159 26333 31171 26367
rect 31113 26327 31171 26333
rect 31202 26324 31208 26376
rect 31260 26324 31266 26376
rect 31220 26296 31248 26324
rect 30576 26268 31248 26296
rect 31404 26237 31432 26404
rect 31757 26367 31815 26373
rect 31757 26333 31769 26367
rect 31803 26364 31815 26367
rect 31803 26336 32168 26364
rect 31803 26333 31815 26336
rect 31757 26327 31815 26333
rect 32140 26308 32168 26336
rect 32030 26305 32036 26308
rect 32024 26296 32036 26305
rect 31991 26268 32036 26296
rect 32024 26259 32036 26268
rect 32030 26256 32036 26259
rect 32088 26256 32094 26308
rect 32122 26256 32128 26308
rect 32180 26256 32186 26308
rect 29748 26200 30052 26228
rect 31389 26231 31447 26237
rect 31389 26197 31401 26231
rect 31435 26228 31447 26231
rect 32784 26228 32812 26460
rect 31435 26200 32812 26228
rect 31435 26197 31447 26200
rect 31389 26191 31447 26197
rect 1104 26138 43884 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 43884 26138
rect 1104 26064 43884 26086
rect 3878 26024 3884 26036
rect 3620 25996 3884 26024
rect 1664 25891 1722 25897
rect 1664 25857 1676 25891
rect 1710 25888 1722 25891
rect 3234 25888 3240 25900
rect 1710 25860 3240 25888
rect 1710 25857 1722 25860
rect 1664 25851 1722 25857
rect 3234 25848 3240 25860
rect 3292 25848 3298 25900
rect 3620 25888 3648 25996
rect 3878 25984 3884 25996
rect 3936 25984 3942 26036
rect 4890 25984 4896 26036
rect 4948 26024 4954 26036
rect 4985 26027 5043 26033
rect 4985 26024 4997 26027
rect 4948 25996 4997 26024
rect 4948 25984 4954 25996
rect 4985 25993 4997 25996
rect 5031 25993 5043 26027
rect 4985 25987 5043 25993
rect 5074 25984 5080 26036
rect 5132 26024 5138 26036
rect 5629 26027 5687 26033
rect 5132 25996 5393 26024
rect 5132 25984 5138 25996
rect 3694 25916 3700 25968
rect 3752 25956 3758 25968
rect 3973 25959 4031 25965
rect 3973 25956 3985 25959
rect 3752 25928 3985 25956
rect 3752 25916 3758 25928
rect 3973 25925 3985 25928
rect 4019 25956 4031 25959
rect 4617 25959 4675 25965
rect 4019 25928 4476 25956
rect 4019 25925 4031 25928
rect 3973 25919 4031 25925
rect 3789 25891 3847 25897
rect 3789 25888 3801 25891
rect 3620 25860 3801 25888
rect 3789 25857 3801 25860
rect 3835 25857 3847 25891
rect 3789 25851 3847 25857
rect 3878 25848 3884 25900
rect 3936 25888 3942 25900
rect 4061 25891 4119 25897
rect 4061 25888 4073 25891
rect 3936 25860 4073 25888
rect 3936 25848 3942 25860
rect 4061 25857 4073 25860
rect 4107 25857 4119 25891
rect 4061 25851 4119 25857
rect 4157 25891 4215 25897
rect 4157 25857 4169 25891
rect 4203 25888 4215 25891
rect 4338 25888 4344 25900
rect 4203 25860 4344 25888
rect 4203 25857 4215 25860
rect 4157 25851 4215 25857
rect 1394 25780 1400 25832
rect 1452 25780 1458 25832
rect 2777 25755 2835 25761
rect 2777 25721 2789 25755
rect 2823 25721 2835 25755
rect 2777 25715 2835 25721
rect 3329 25755 3387 25761
rect 3329 25721 3341 25755
rect 3375 25752 3387 25755
rect 4172 25752 4200 25851
rect 4338 25848 4344 25860
rect 4396 25848 4402 25900
rect 4448 25897 4476 25928
rect 4617 25925 4629 25959
rect 4663 25956 4675 25959
rect 5166 25956 5172 25968
rect 4663 25928 5172 25956
rect 4663 25925 4675 25928
rect 4617 25919 4675 25925
rect 5166 25916 5172 25928
rect 5224 25916 5230 25968
rect 5365 25956 5393 25996
rect 5629 25993 5641 26027
rect 5675 26024 5687 26027
rect 5810 26024 5816 26036
rect 5675 25996 5816 26024
rect 5675 25993 5687 25996
rect 5629 25987 5687 25993
rect 5810 25984 5816 25996
rect 5868 25984 5874 26036
rect 6730 25984 6736 26036
rect 6788 26024 6794 26036
rect 6788 25996 8984 26024
rect 6788 25984 6794 25996
rect 7926 25956 7932 25968
rect 5365 25928 7932 25956
rect 4433 25891 4491 25897
rect 4433 25857 4445 25891
rect 4479 25857 4491 25891
rect 4433 25851 4491 25857
rect 4448 25820 4476 25851
rect 4706 25848 4712 25900
rect 4764 25848 4770 25900
rect 4801 25891 4859 25897
rect 4801 25857 4813 25891
rect 4847 25888 4859 25891
rect 4982 25888 4988 25900
rect 4847 25860 4988 25888
rect 4847 25857 4859 25860
rect 4801 25851 4859 25857
rect 4982 25848 4988 25860
rect 5040 25848 5046 25900
rect 5074 25848 5080 25900
rect 5132 25848 5138 25900
rect 5258 25848 5264 25900
rect 5316 25848 5322 25900
rect 5353 25891 5411 25897
rect 5353 25857 5365 25891
rect 5399 25857 5411 25891
rect 5353 25851 5411 25857
rect 5491 25891 5549 25897
rect 5491 25857 5503 25891
rect 5537 25888 5549 25891
rect 5626 25888 5632 25900
rect 5537 25860 5632 25888
rect 5537 25857 5549 25860
rect 5491 25851 5549 25857
rect 3375 25724 4200 25752
rect 4264 25792 4476 25820
rect 3375 25721 3387 25724
rect 3329 25715 3387 25721
rect 2792 25684 2820 25715
rect 3970 25684 3976 25696
rect 2792 25656 3976 25684
rect 3970 25644 3976 25656
rect 4028 25644 4034 25696
rect 4264 25684 4292 25792
rect 4614 25780 4620 25832
rect 4672 25820 4678 25832
rect 5365 25820 5393 25851
rect 5626 25848 5632 25860
rect 5684 25848 5690 25900
rect 5718 25848 5724 25900
rect 5776 25888 5782 25900
rect 6546 25888 6552 25900
rect 5776 25860 6552 25888
rect 5776 25848 5782 25860
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 6748 25897 6776 25928
rect 7926 25916 7932 25928
rect 7984 25916 7990 25968
rect 8021 25959 8079 25965
rect 8021 25925 8033 25959
rect 8067 25956 8079 25959
rect 8389 25959 8447 25965
rect 8067 25928 8340 25956
rect 8067 25925 8079 25928
rect 8021 25919 8079 25925
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 6917 25891 6975 25897
rect 6917 25857 6929 25891
rect 6963 25857 6975 25891
rect 6917 25851 6975 25857
rect 4672 25792 5393 25820
rect 4672 25780 4678 25792
rect 6362 25780 6368 25832
rect 6420 25780 6426 25832
rect 6932 25820 6960 25851
rect 7006 25848 7012 25900
rect 7064 25848 7070 25900
rect 7098 25848 7104 25900
rect 7156 25848 7162 25900
rect 8036 25888 8064 25919
rect 8312 25900 8340 25928
rect 8389 25925 8401 25959
rect 8435 25956 8447 25959
rect 8478 25956 8484 25968
rect 8435 25928 8484 25956
rect 8435 25925 8447 25928
rect 8389 25919 8447 25925
rect 8478 25916 8484 25928
rect 8536 25916 8542 25968
rect 8956 25956 8984 25996
rect 9030 25984 9036 26036
rect 9088 25984 9094 26036
rect 9490 25984 9496 26036
rect 9548 26024 9554 26036
rect 10042 26024 10048 26036
rect 9548 25996 10048 26024
rect 9548 25984 9554 25996
rect 10042 25984 10048 25996
rect 10100 25984 10106 26036
rect 10318 25984 10324 26036
rect 10376 26024 10382 26036
rect 11333 26027 11391 26033
rect 10376 25996 11192 26024
rect 10376 25984 10382 25996
rect 10686 25956 10692 25968
rect 8956 25928 10692 25956
rect 10686 25916 10692 25928
rect 10744 25916 10750 25968
rect 10962 25916 10968 25968
rect 11020 25916 11026 25968
rect 11054 25916 11060 25968
rect 11112 25916 11118 25968
rect 7208 25860 8064 25888
rect 7208 25820 7236 25860
rect 8294 25848 8300 25900
rect 8352 25848 8358 25900
rect 8849 25891 8907 25897
rect 8849 25857 8861 25891
rect 8895 25888 8907 25891
rect 9030 25888 9036 25900
rect 8895 25860 9036 25888
rect 8895 25857 8907 25860
rect 8849 25851 8907 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25888 9183 25891
rect 9171 25860 9674 25888
rect 9171 25857 9183 25860
rect 9125 25851 9183 25857
rect 6932 25792 7236 25820
rect 8018 25780 8024 25832
rect 8076 25780 8082 25832
rect 8202 25780 8208 25832
rect 8260 25820 8266 25832
rect 9140 25820 9168 25851
rect 8260 25792 9168 25820
rect 9646 25820 9674 25860
rect 10502 25848 10508 25900
rect 10560 25888 10566 25900
rect 10597 25891 10655 25897
rect 10597 25888 10609 25891
rect 10560 25860 10609 25888
rect 10560 25848 10566 25860
rect 10597 25857 10609 25860
rect 10643 25857 10655 25891
rect 10597 25851 10655 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 10870 25888 10876 25900
rect 10827 25860 10876 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 11164 25897 11192 25996
rect 11333 25993 11345 26027
rect 11379 26024 11391 26027
rect 11606 26024 11612 26036
rect 11379 25996 11612 26024
rect 11379 25993 11391 25996
rect 11333 25987 11391 25993
rect 11606 25984 11612 25996
rect 11664 25984 11670 26036
rect 11701 26027 11759 26033
rect 11701 25993 11713 26027
rect 11747 26024 11759 26027
rect 12434 26024 12440 26036
rect 11747 25996 12440 26024
rect 11747 25993 11759 25996
rect 11701 25987 11759 25993
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 13446 25984 13452 26036
rect 13504 25984 13510 26036
rect 13814 25984 13820 26036
rect 13872 26024 13878 26036
rect 14366 26024 14372 26036
rect 13872 25996 14372 26024
rect 13872 25984 13878 25996
rect 14366 25984 14372 25996
rect 14424 25984 14430 26036
rect 15286 25984 15292 26036
rect 15344 26024 15350 26036
rect 15381 26027 15439 26033
rect 15381 26024 15393 26027
rect 15344 25996 15393 26024
rect 15344 25984 15350 25996
rect 15381 25993 15393 25996
rect 15427 25993 15439 26027
rect 15381 25987 15439 25993
rect 15654 25984 15660 26036
rect 15712 26024 15718 26036
rect 16482 26024 16488 26036
rect 15712 25996 16488 26024
rect 15712 25984 15718 25996
rect 16482 25984 16488 25996
rect 16540 25984 16546 26036
rect 16666 25984 16672 26036
rect 16724 25984 16730 26036
rect 19978 25984 19984 26036
rect 20036 25984 20042 26036
rect 20070 25984 20076 26036
rect 20128 26024 20134 26036
rect 20165 26027 20223 26033
rect 20165 26024 20177 26027
rect 20128 25996 20177 26024
rect 20128 25984 20134 25996
rect 20165 25993 20177 25996
rect 20211 25993 20223 26027
rect 20165 25987 20223 25993
rect 20257 26027 20315 26033
rect 20257 25993 20269 26027
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 11514 25916 11520 25968
rect 11572 25916 11578 25968
rect 12161 25959 12219 25965
rect 12161 25956 12173 25959
rect 11716 25928 12173 25956
rect 11149 25891 11207 25897
rect 11149 25857 11161 25891
rect 11195 25888 11207 25891
rect 11716 25888 11744 25928
rect 12161 25925 12173 25928
rect 12207 25956 12219 25959
rect 15933 25959 15991 25965
rect 12207 25928 12848 25956
rect 12207 25925 12219 25928
rect 12161 25919 12219 25925
rect 11195 25860 11744 25888
rect 11793 25891 11851 25897
rect 11195 25857 11207 25860
rect 11149 25851 11207 25857
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 11839 25860 12296 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 11808 25820 11836 25851
rect 9646 25792 11836 25820
rect 8260 25780 8266 25792
rect 12158 25780 12164 25832
rect 12216 25820 12222 25832
rect 12268 25820 12296 25860
rect 12820 25832 12848 25928
rect 15933 25925 15945 25959
rect 15979 25956 15991 25959
rect 16390 25956 16396 25968
rect 15979 25928 16396 25956
rect 15979 25925 15991 25928
rect 15933 25919 15991 25925
rect 16390 25916 16396 25928
rect 16448 25916 16454 25968
rect 16684 25956 16712 25984
rect 16500 25928 16712 25956
rect 17681 25959 17739 25965
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 13909 25891 13967 25897
rect 13909 25857 13921 25891
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 12216 25792 12296 25820
rect 12216 25780 12222 25792
rect 4341 25755 4399 25761
rect 4341 25721 4353 25755
rect 4387 25752 4399 25755
rect 6380 25752 6408 25780
rect 8036 25752 8064 25780
rect 8478 25752 8484 25764
rect 4387 25724 6408 25752
rect 6569 25724 7880 25752
rect 8036 25724 8484 25752
rect 4387 25721 4399 25724
rect 4341 25715 4399 25721
rect 5074 25684 5080 25696
rect 4264 25656 5080 25684
rect 5074 25644 5080 25656
rect 5132 25644 5138 25696
rect 5626 25644 5632 25696
rect 5684 25684 5690 25696
rect 5997 25687 6055 25693
rect 5997 25684 6009 25687
rect 5684 25656 6009 25684
rect 5684 25644 5690 25656
rect 5997 25653 6009 25656
rect 6043 25684 6055 25687
rect 6569 25684 6597 25724
rect 6043 25656 6597 25684
rect 6043 25653 6055 25656
rect 5997 25647 6055 25653
rect 6638 25644 6644 25696
rect 6696 25644 6702 25696
rect 7282 25644 7288 25696
rect 7340 25644 7346 25696
rect 7561 25687 7619 25693
rect 7561 25653 7573 25687
rect 7607 25684 7619 25687
rect 7742 25684 7748 25696
rect 7607 25656 7748 25684
rect 7607 25653 7619 25656
rect 7561 25647 7619 25653
rect 7742 25644 7748 25656
rect 7800 25644 7806 25696
rect 7852 25684 7880 25724
rect 8478 25712 8484 25724
rect 8536 25712 8542 25764
rect 8754 25712 8760 25764
rect 8812 25752 8818 25764
rect 8849 25755 8907 25761
rect 8849 25752 8861 25755
rect 8812 25724 8861 25752
rect 8812 25712 8818 25724
rect 8849 25721 8861 25724
rect 8895 25721 8907 25755
rect 8849 25715 8907 25721
rect 11330 25712 11336 25764
rect 11388 25752 11394 25764
rect 11517 25755 11575 25761
rect 11517 25752 11529 25755
rect 11388 25724 11529 25752
rect 11388 25712 11394 25724
rect 11517 25721 11529 25724
rect 11563 25721 11575 25755
rect 11517 25715 11575 25721
rect 8570 25684 8576 25696
rect 7852 25656 8576 25684
rect 8570 25644 8576 25656
rect 8628 25684 8634 25696
rect 8665 25687 8723 25693
rect 8665 25684 8677 25687
rect 8628 25656 8677 25684
rect 8628 25644 8634 25656
rect 8665 25653 8677 25656
rect 8711 25684 8723 25687
rect 9306 25684 9312 25696
rect 8711 25656 9312 25684
rect 8711 25653 8723 25656
rect 8665 25647 8723 25653
rect 9306 25644 9312 25656
rect 9364 25684 9370 25696
rect 9861 25687 9919 25693
rect 9861 25684 9873 25687
rect 9364 25656 9873 25684
rect 9364 25644 9370 25656
rect 9861 25653 9873 25656
rect 9907 25684 9919 25687
rect 11054 25684 11060 25696
rect 9907 25656 11060 25684
rect 9907 25653 9919 25656
rect 9861 25647 9919 25653
rect 11054 25644 11060 25656
rect 11112 25684 11118 25696
rect 11974 25684 11980 25696
rect 11112 25656 11980 25684
rect 11112 25644 11118 25656
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12268 25684 12296 25792
rect 12802 25780 12808 25832
rect 12860 25780 12866 25832
rect 13924 25820 13952 25851
rect 14182 25848 14188 25900
rect 14240 25888 14246 25900
rect 14553 25891 14611 25897
rect 14553 25888 14565 25891
rect 14240 25860 14565 25888
rect 14240 25848 14246 25860
rect 14553 25857 14565 25860
rect 14599 25888 14611 25891
rect 15470 25888 15476 25900
rect 14599 25860 15476 25888
rect 14599 25857 14611 25860
rect 14553 25851 14611 25857
rect 15470 25848 15476 25860
rect 15528 25848 15534 25900
rect 15565 25891 15623 25897
rect 15565 25857 15577 25891
rect 15611 25888 15623 25891
rect 15654 25888 15660 25900
rect 15611 25860 15660 25888
rect 15611 25857 15623 25860
rect 15565 25851 15623 25857
rect 15654 25848 15660 25860
rect 15712 25848 15718 25900
rect 15838 25848 15844 25900
rect 15896 25848 15902 25900
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16209 25891 16267 25897
rect 16209 25857 16221 25891
rect 16255 25888 16267 25891
rect 16500 25888 16528 25928
rect 17681 25925 17693 25959
rect 17727 25956 17739 25959
rect 17954 25956 17960 25968
rect 17727 25928 17960 25956
rect 17727 25925 17739 25928
rect 17681 25919 17739 25925
rect 17954 25916 17960 25928
rect 18012 25916 18018 25968
rect 19996 25956 20024 25984
rect 20272 25956 20300 25987
rect 20530 25984 20536 26036
rect 20588 26024 20594 26036
rect 20625 26027 20683 26033
rect 20625 26024 20637 26027
rect 20588 25996 20637 26024
rect 20588 25984 20594 25996
rect 20625 25993 20637 25996
rect 20671 25993 20683 26027
rect 20625 25987 20683 25993
rect 20916 25996 21128 26024
rect 20916 25956 20944 25996
rect 19628 25928 20024 25956
rect 20088 25928 20300 25956
rect 20640 25928 20944 25956
rect 21100 25956 21128 25996
rect 21634 25984 21640 26036
rect 21692 25984 21698 26036
rect 23382 25984 23388 26036
rect 23440 26024 23446 26036
rect 26697 26027 26755 26033
rect 26697 26024 26709 26027
rect 23440 25996 26709 26024
rect 23440 25984 23446 25996
rect 26697 25993 26709 25996
rect 26743 26024 26755 26027
rect 27890 26024 27896 26036
rect 26743 25996 27896 26024
rect 26743 25993 26755 25996
rect 26697 25987 26755 25993
rect 21100 25928 21211 25956
rect 16255 25860 16528 25888
rect 16255 25857 16267 25860
rect 16209 25851 16267 25857
rect 16132 25820 16160 25851
rect 16408 25832 16436 25860
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 16632 25860 16681 25888
rect 16632 25848 16638 25860
rect 16669 25857 16681 25860
rect 16715 25888 16727 25891
rect 17497 25891 17555 25897
rect 17497 25888 17509 25891
rect 16715 25860 17509 25888
rect 16715 25857 16727 25860
rect 16669 25851 16727 25857
rect 17497 25857 17509 25860
rect 17543 25857 17555 25891
rect 17497 25851 17555 25857
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25888 17923 25891
rect 18598 25888 18604 25900
rect 17911 25860 18604 25888
rect 17911 25857 17923 25860
rect 17865 25851 17923 25857
rect 18598 25848 18604 25860
rect 18656 25848 18662 25900
rect 19058 25848 19064 25900
rect 19116 25848 19122 25900
rect 19628 25897 19656 25928
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25888 20039 25891
rect 20088 25888 20116 25928
rect 20640 25888 20668 25928
rect 20027 25860 20116 25888
rect 20180 25860 20668 25888
rect 20027 25857 20039 25860
rect 19981 25851 20039 25857
rect 13924 25792 15700 25820
rect 12526 25712 12532 25764
rect 12584 25752 12590 25764
rect 13262 25752 13268 25764
rect 12584 25724 13268 25752
rect 12584 25712 12590 25724
rect 13262 25712 13268 25724
rect 13320 25712 13326 25764
rect 13924 25684 13952 25792
rect 15672 25764 15700 25792
rect 15764 25792 16160 25820
rect 15764 25764 15792 25792
rect 16390 25780 16396 25832
rect 16448 25780 16454 25832
rect 16482 25780 16488 25832
rect 16540 25820 16546 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 16540 25792 18061 25820
rect 16540 25780 16546 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 19076 25820 19104 25848
rect 20180 25820 20208 25860
rect 20714 25848 20720 25900
rect 20772 25888 20778 25900
rect 20772 25860 20944 25888
rect 20772 25848 20778 25860
rect 19076 25792 20208 25820
rect 18049 25783 18107 25789
rect 20806 25780 20812 25832
rect 20864 25780 20870 25832
rect 20916 25820 20944 25860
rect 20990 25848 20996 25900
rect 21048 25888 21054 25900
rect 21085 25891 21143 25897
rect 21085 25888 21097 25891
rect 21048 25860 21097 25888
rect 21048 25848 21054 25860
rect 21085 25857 21097 25860
rect 21131 25857 21143 25891
rect 21183 25888 21211 25928
rect 24394 25916 24400 25968
rect 24452 25916 24458 25968
rect 25685 25959 25743 25965
rect 25685 25956 25697 25959
rect 24596 25928 25697 25956
rect 22097 25891 22155 25897
rect 22097 25888 22109 25891
rect 21183 25860 22109 25888
rect 21085 25851 21143 25857
rect 22097 25857 22109 25860
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 21634 25820 21640 25832
rect 20916 25792 21640 25820
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22112 25820 22140 25851
rect 22462 25848 22468 25900
rect 22520 25848 22526 25900
rect 22922 25848 22928 25900
rect 22980 25848 22986 25900
rect 23198 25848 23204 25900
rect 23256 25888 23262 25900
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 23256 25860 23305 25888
rect 23256 25848 23262 25860
rect 23293 25857 23305 25860
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 23658 25848 23664 25900
rect 23716 25848 23722 25900
rect 24210 25848 24216 25900
rect 24268 25848 24274 25900
rect 24596 25886 24624 25928
rect 25685 25925 25697 25928
rect 25731 25956 25743 25959
rect 25774 25956 25780 25968
rect 25731 25928 25780 25956
rect 25731 25925 25743 25928
rect 25685 25919 25743 25925
rect 25774 25916 25780 25928
rect 25832 25916 25838 25968
rect 25958 25916 25964 25968
rect 26016 25956 26022 25968
rect 26988 25965 27016 25996
rect 27890 25984 27896 25996
rect 27948 25984 27954 26036
rect 27982 25984 27988 26036
rect 28040 26024 28046 26036
rect 28810 26024 28816 26036
rect 28040 25996 28816 26024
rect 28040 25984 28046 25996
rect 28810 25984 28816 25996
rect 28868 25984 28874 26036
rect 29546 25984 29552 26036
rect 29604 26024 29610 26036
rect 29604 25996 29684 26024
rect 29604 25984 29610 25996
rect 26053 25959 26111 25965
rect 26053 25956 26065 25959
rect 26016 25928 26065 25956
rect 26016 25916 26022 25928
rect 26053 25925 26065 25928
rect 26099 25925 26111 25959
rect 26053 25919 26111 25925
rect 26973 25959 27031 25965
rect 26973 25925 26985 25959
rect 27019 25925 27031 25959
rect 26973 25919 27031 25925
rect 27338 25916 27344 25968
rect 27396 25916 27402 25968
rect 27706 25916 27712 25968
rect 27764 25956 27770 25968
rect 29454 25956 29460 25968
rect 27764 25928 29460 25956
rect 27764 25916 27770 25928
rect 29454 25916 29460 25928
rect 29512 25956 29518 25968
rect 29656 25956 29684 25996
rect 32582 25984 32588 26036
rect 32640 26024 32646 26036
rect 33505 26027 33563 26033
rect 33505 26024 33517 26027
rect 32640 25996 33517 26024
rect 32640 25984 32646 25996
rect 33505 25993 33517 25996
rect 33551 25993 33563 26027
rect 33505 25987 33563 25993
rect 29794 25959 29852 25965
rect 29794 25956 29806 25959
rect 29512 25928 29592 25956
rect 29656 25928 29806 25956
rect 29512 25916 29518 25928
rect 24505 25858 24624 25886
rect 23474 25820 23480 25832
rect 22112 25792 23480 25820
rect 23474 25780 23480 25792
rect 23532 25780 23538 25832
rect 23937 25823 23995 25829
rect 23937 25789 23949 25823
rect 23983 25820 23995 25823
rect 24118 25820 24124 25832
rect 23983 25792 24124 25820
rect 23983 25789 23995 25792
rect 23937 25783 23995 25789
rect 24118 25780 24124 25792
rect 24176 25780 24182 25832
rect 24302 25780 24308 25832
rect 24360 25820 24366 25832
rect 24505 25820 24533 25858
rect 25590 25848 25596 25900
rect 25648 25888 25654 25900
rect 25869 25891 25927 25897
rect 25869 25888 25881 25891
rect 25648 25860 25881 25888
rect 25648 25848 25654 25860
rect 25869 25857 25881 25860
rect 25915 25888 25927 25891
rect 26145 25891 26203 25897
rect 25915 25860 26096 25888
rect 25915 25857 25927 25860
rect 25869 25851 25927 25857
rect 26068 25832 26096 25860
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 24360 25792 24533 25820
rect 24581 25823 24639 25829
rect 24360 25780 24366 25792
rect 24581 25789 24593 25823
rect 24627 25820 24639 25823
rect 24854 25820 24860 25832
rect 24627 25792 24860 25820
rect 24627 25789 24639 25792
rect 24581 25783 24639 25789
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 25222 25780 25228 25832
rect 25280 25780 25286 25832
rect 26050 25780 26056 25832
rect 26108 25780 26114 25832
rect 14844 25724 15614 25752
rect 12268 25656 13952 25684
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 14844 25693 14872 25724
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 14516 25656 14841 25684
rect 14516 25644 14522 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 14829 25647 14887 25653
rect 15286 25644 15292 25696
rect 15344 25644 15350 25696
rect 15586 25684 15614 25724
rect 15654 25712 15660 25764
rect 15712 25712 15718 25764
rect 15746 25712 15752 25764
rect 15804 25712 15810 25764
rect 15930 25712 15936 25764
rect 15988 25712 15994 25764
rect 16666 25752 16672 25764
rect 16040 25724 16672 25752
rect 16040 25684 16068 25724
rect 16666 25712 16672 25724
rect 16724 25752 16730 25764
rect 17129 25755 17187 25761
rect 17129 25752 17141 25755
rect 16724 25724 17141 25752
rect 16724 25712 16730 25724
rect 17129 25721 17141 25724
rect 17175 25752 17187 25755
rect 18230 25752 18236 25764
rect 17175 25724 18236 25752
rect 17175 25721 17187 25724
rect 17129 25715 17187 25721
rect 18230 25712 18236 25724
rect 18288 25712 18294 25764
rect 19242 25712 19248 25764
rect 19300 25752 19306 25764
rect 19300 25724 21496 25752
rect 19300 25712 19306 25724
rect 21468 25696 21496 25724
rect 22370 25712 22376 25764
rect 22428 25752 22434 25764
rect 26160 25752 26188 25851
rect 26234 25848 26240 25900
rect 26292 25848 26298 25900
rect 27356 25820 27384 25916
rect 28166 25848 28172 25900
rect 28224 25888 28230 25900
rect 29564 25897 29592 25928
rect 29794 25925 29806 25928
rect 29840 25925 29852 25959
rect 29794 25919 29852 25925
rect 31846 25916 31852 25968
rect 31904 25956 31910 25968
rect 32370 25959 32428 25965
rect 32370 25956 32382 25959
rect 31904 25928 32382 25956
rect 31904 25916 31910 25928
rect 32370 25925 32382 25928
rect 32416 25925 32428 25959
rect 32370 25919 32428 25925
rect 28353 25891 28411 25897
rect 28353 25888 28365 25891
rect 28224 25860 28365 25888
rect 28224 25848 28230 25860
rect 28353 25857 28365 25860
rect 28399 25857 28411 25891
rect 28353 25851 28411 25857
rect 28537 25891 28595 25897
rect 28537 25857 28549 25891
rect 28583 25857 28595 25891
rect 28537 25851 28595 25857
rect 28629 25891 28687 25897
rect 28629 25857 28641 25891
rect 28675 25888 28687 25891
rect 29549 25891 29607 25897
rect 28675 25860 29500 25888
rect 28675 25857 28687 25860
rect 28629 25851 28687 25857
rect 28442 25820 28448 25832
rect 27356 25792 28448 25820
rect 28442 25780 28448 25792
rect 28500 25820 28506 25832
rect 28552 25820 28580 25851
rect 28500 25792 28580 25820
rect 28500 25780 28506 25792
rect 28902 25780 28908 25832
rect 28960 25780 28966 25832
rect 29472 25820 29500 25860
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 30098 25888 30104 25900
rect 29549 25851 29607 25857
rect 29656 25860 30104 25888
rect 29656 25820 29684 25860
rect 30098 25848 30104 25860
rect 30156 25848 30162 25900
rect 32122 25848 32128 25900
rect 32180 25848 32186 25900
rect 29472 25792 29684 25820
rect 31110 25780 31116 25832
rect 31168 25780 31174 25832
rect 31389 25823 31447 25829
rect 31389 25789 31401 25823
rect 31435 25789 31447 25823
rect 31389 25783 31447 25789
rect 27706 25752 27712 25764
rect 22428 25724 26188 25752
rect 26349 25724 27712 25752
rect 22428 25712 22434 25724
rect 15586 25656 16068 25684
rect 16206 25644 16212 25696
rect 16264 25684 16270 25696
rect 16761 25687 16819 25693
rect 16761 25684 16773 25687
rect 16264 25656 16773 25684
rect 16264 25644 16270 25656
rect 16761 25653 16773 25656
rect 16807 25653 16819 25687
rect 16761 25647 16819 25653
rect 17494 25644 17500 25696
rect 17552 25684 17558 25696
rect 18325 25687 18383 25693
rect 18325 25684 18337 25687
rect 17552 25656 18337 25684
rect 17552 25644 17558 25656
rect 18325 25653 18337 25656
rect 18371 25653 18383 25687
rect 18325 25647 18383 25653
rect 18506 25644 18512 25696
rect 18564 25684 18570 25696
rect 18693 25687 18751 25693
rect 18693 25684 18705 25687
rect 18564 25656 18705 25684
rect 18564 25644 18570 25656
rect 18693 25653 18705 25656
rect 18739 25653 18751 25687
rect 18693 25647 18751 25653
rect 19150 25644 19156 25696
rect 19208 25644 19214 25696
rect 19521 25687 19579 25693
rect 19521 25653 19533 25687
rect 19567 25684 19579 25687
rect 19886 25684 19892 25696
rect 19567 25656 19892 25684
rect 19567 25653 19579 25656
rect 19521 25647 19579 25653
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 19981 25687 20039 25693
rect 19981 25653 19993 25687
rect 20027 25684 20039 25687
rect 20622 25684 20628 25696
rect 20027 25656 20628 25684
rect 20027 25653 20039 25656
rect 19981 25647 20039 25653
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 21082 25644 21088 25696
rect 21140 25684 21146 25696
rect 21177 25687 21235 25693
rect 21177 25684 21189 25687
rect 21140 25656 21189 25684
rect 21140 25644 21146 25656
rect 21177 25653 21189 25656
rect 21223 25653 21235 25687
rect 21177 25647 21235 25653
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 23382 25644 23388 25696
rect 23440 25684 23446 25696
rect 24857 25687 24915 25693
rect 24857 25684 24869 25687
rect 23440 25656 24869 25684
rect 23440 25644 23446 25656
rect 24857 25653 24869 25656
rect 24903 25684 24915 25687
rect 26349 25684 26377 25724
rect 27706 25712 27712 25724
rect 27764 25712 27770 25764
rect 28258 25712 28264 25764
rect 28316 25752 28322 25764
rect 28316 25724 28488 25752
rect 28316 25712 28322 25724
rect 24903 25656 26377 25684
rect 26421 25687 26479 25693
rect 24903 25653 24915 25656
rect 24857 25647 24915 25653
rect 26421 25653 26433 25687
rect 26467 25684 26479 25687
rect 26786 25684 26792 25696
rect 26467 25656 26792 25684
rect 26467 25653 26479 25656
rect 26421 25647 26479 25653
rect 26786 25644 26792 25656
rect 26844 25644 26850 25696
rect 27614 25644 27620 25696
rect 27672 25684 27678 25696
rect 28353 25687 28411 25693
rect 28353 25684 28365 25687
rect 27672 25656 28365 25684
rect 27672 25644 27678 25656
rect 28353 25653 28365 25656
rect 28399 25653 28411 25687
rect 28460 25684 28488 25724
rect 28718 25712 28724 25764
rect 28776 25752 28782 25764
rect 29086 25752 29092 25764
rect 28776 25724 29092 25752
rect 28776 25712 28782 25724
rect 29086 25712 29092 25724
rect 29144 25712 29150 25764
rect 29178 25712 29184 25764
rect 29236 25752 29242 25764
rect 29546 25752 29552 25764
rect 29236 25724 29552 25752
rect 29236 25712 29242 25724
rect 29546 25712 29552 25724
rect 29604 25712 29610 25764
rect 30926 25712 30932 25764
rect 30984 25712 30990 25764
rect 30834 25684 30840 25696
rect 28460 25656 30840 25684
rect 28353 25647 28411 25653
rect 30834 25644 30840 25656
rect 30892 25684 30898 25696
rect 31404 25684 31432 25783
rect 30892 25656 31432 25684
rect 30892 25644 30898 25656
rect 1104 25594 43884 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 43884 25594
rect 1104 25520 43884 25542
rect 2777 25483 2835 25489
rect 2777 25449 2789 25483
rect 2823 25449 2835 25483
rect 2777 25443 2835 25449
rect 2792 25412 2820 25443
rect 3234 25440 3240 25492
rect 3292 25440 3298 25492
rect 3605 25483 3663 25489
rect 3605 25449 3617 25483
rect 3651 25480 3663 25483
rect 3694 25480 3700 25492
rect 3651 25452 3700 25480
rect 3651 25449 3663 25452
rect 3605 25443 3663 25449
rect 3694 25440 3700 25452
rect 3752 25440 3758 25492
rect 5258 25440 5264 25492
rect 5316 25440 5322 25492
rect 5442 25440 5448 25492
rect 5500 25480 5506 25492
rect 5629 25483 5687 25489
rect 5629 25480 5641 25483
rect 5500 25452 5641 25480
rect 5500 25440 5506 25452
rect 5629 25449 5641 25452
rect 5675 25449 5687 25483
rect 5629 25443 5687 25449
rect 6178 25440 6184 25492
rect 6236 25480 6242 25492
rect 6236 25452 7604 25480
rect 6236 25440 6242 25452
rect 3326 25412 3332 25424
rect 2792 25384 3332 25412
rect 3326 25372 3332 25384
rect 3384 25412 3390 25424
rect 3878 25412 3884 25424
rect 3384 25384 3884 25412
rect 3384 25372 3390 25384
rect 3878 25372 3884 25384
rect 3936 25372 3942 25424
rect 2682 25304 2688 25356
rect 2740 25344 2746 25356
rect 4706 25344 4712 25356
rect 2740 25316 4712 25344
rect 2740 25304 2746 25316
rect 4706 25304 4712 25316
rect 4764 25304 4770 25356
rect 5276 25344 5304 25440
rect 5752 25384 7053 25412
rect 5752 25344 5780 25384
rect 6822 25344 6828 25356
rect 5092 25316 5304 25344
rect 5368 25316 5780 25344
rect 6242 25316 6828 25344
rect 1394 25236 1400 25288
rect 1452 25276 1458 25288
rect 2038 25276 2044 25288
rect 1452 25248 2044 25276
rect 1452 25236 1458 25248
rect 2038 25236 2044 25248
rect 2096 25236 2102 25288
rect 2869 25279 2927 25285
rect 2869 25245 2881 25279
rect 2915 25245 2927 25279
rect 2869 25239 2927 25245
rect 1664 25211 1722 25217
rect 1664 25177 1676 25211
rect 1710 25208 1722 25211
rect 1762 25208 1768 25220
rect 1710 25180 1768 25208
rect 1710 25177 1722 25180
rect 1664 25171 1722 25177
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 1486 25100 1492 25152
rect 1544 25140 1550 25152
rect 2884 25140 2912 25239
rect 3050 25236 3056 25288
rect 3108 25236 3114 25288
rect 3881 25279 3939 25285
rect 3881 25245 3893 25279
rect 3927 25276 3939 25279
rect 3970 25276 3976 25288
rect 3927 25248 3976 25276
rect 3927 25245 3939 25248
rect 3881 25239 3939 25245
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 5092 25285 5120 25316
rect 5077 25279 5135 25285
rect 5077 25276 5089 25279
rect 4080 25248 5089 25276
rect 4080 25208 4108 25248
rect 5077 25245 5089 25248
rect 5123 25245 5135 25279
rect 5077 25239 5135 25245
rect 5166 25236 5172 25288
rect 5224 25276 5230 25288
rect 5368 25285 5396 25316
rect 5261 25279 5319 25285
rect 5261 25276 5273 25279
rect 5224 25248 5273 25276
rect 5224 25236 5230 25248
rect 5261 25245 5273 25248
rect 5307 25245 5319 25279
rect 5261 25239 5319 25245
rect 5353 25279 5411 25285
rect 5353 25245 5365 25279
rect 5399 25245 5411 25279
rect 5353 25239 5411 25245
rect 5445 25279 5503 25285
rect 5445 25245 5457 25279
rect 5491 25276 5503 25279
rect 5626 25276 5632 25288
rect 5491 25248 5632 25276
rect 5491 25245 5503 25248
rect 5445 25239 5503 25245
rect 3436 25180 4108 25208
rect 3436 25152 3464 25180
rect 4982 25168 4988 25220
rect 5040 25208 5046 25220
rect 5460 25208 5488 25239
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 5718 25236 5724 25288
rect 5776 25236 5782 25288
rect 5810 25236 5816 25288
rect 5868 25276 5874 25288
rect 5868 25248 5913 25276
rect 5868 25236 5874 25248
rect 5994 25236 6000 25288
rect 6052 25236 6058 25288
rect 6242 25285 6270 25316
rect 6822 25304 6828 25316
rect 6880 25304 6886 25356
rect 7025 25344 7053 25384
rect 7190 25372 7196 25424
rect 7248 25372 7254 25424
rect 7374 25372 7380 25424
rect 7432 25372 7438 25424
rect 7392 25344 7420 25372
rect 7025 25316 7420 25344
rect 6227 25279 6285 25285
rect 6227 25245 6239 25279
rect 6273 25245 6285 25279
rect 6227 25239 6285 25245
rect 6454 25236 6460 25288
rect 6512 25236 6518 25288
rect 6546 25236 6552 25288
rect 6604 25276 6610 25288
rect 6604 25248 6649 25276
rect 6604 25236 6610 25248
rect 6730 25236 6736 25288
rect 6788 25236 6794 25288
rect 6840 25276 6868 25304
rect 6922 25279 6980 25285
rect 6922 25276 6934 25279
rect 6840 25248 6934 25276
rect 6922 25245 6934 25248
rect 6968 25245 6980 25279
rect 6922 25239 6980 25245
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7576 25285 7604 25452
rect 8478 25440 8484 25492
rect 8536 25480 8542 25492
rect 8665 25483 8723 25489
rect 8665 25480 8677 25483
rect 8536 25452 8677 25480
rect 8536 25440 8542 25452
rect 8665 25449 8677 25452
rect 8711 25449 8723 25483
rect 8665 25443 8723 25449
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9493 25483 9551 25489
rect 9493 25480 9505 25483
rect 8812 25452 9505 25480
rect 8812 25440 8818 25452
rect 9493 25449 9505 25452
rect 9539 25449 9551 25483
rect 9493 25443 9551 25449
rect 10413 25483 10471 25489
rect 10413 25449 10425 25483
rect 10459 25480 10471 25483
rect 11514 25480 11520 25492
rect 10459 25452 11520 25480
rect 10459 25449 10471 25452
rect 10413 25443 10471 25449
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 11974 25440 11980 25492
rect 12032 25440 12038 25492
rect 14274 25440 14280 25492
rect 14332 25480 14338 25492
rect 14645 25483 14703 25489
rect 14645 25480 14657 25483
rect 14332 25452 14657 25480
rect 14332 25440 14338 25452
rect 14645 25449 14657 25452
rect 14691 25449 14703 25483
rect 14645 25443 14703 25449
rect 14734 25440 14740 25492
rect 14792 25480 14798 25492
rect 15473 25483 15531 25489
rect 15473 25480 15485 25483
rect 14792 25452 15485 25480
rect 14792 25440 14798 25452
rect 15473 25449 15485 25452
rect 15519 25449 15531 25483
rect 15473 25443 15531 25449
rect 15933 25483 15991 25489
rect 15933 25449 15945 25483
rect 15979 25480 15991 25483
rect 16206 25480 16212 25492
rect 15979 25452 16212 25480
rect 15979 25449 15991 25452
rect 15933 25443 15991 25449
rect 7929 25415 7987 25421
rect 7929 25381 7941 25415
rect 7975 25412 7987 25415
rect 8294 25412 8300 25424
rect 7975 25384 8300 25412
rect 7975 25381 7987 25384
rect 7929 25375 7987 25381
rect 8128 25285 8156 25384
rect 8294 25372 8300 25384
rect 8352 25372 8358 25424
rect 10226 25372 10232 25424
rect 10284 25412 10290 25424
rect 11057 25415 11115 25421
rect 11057 25412 11069 25415
rect 10284 25384 11069 25412
rect 10284 25372 10290 25384
rect 11057 25381 11069 25384
rect 11103 25381 11115 25415
rect 11057 25375 11115 25381
rect 11164 25384 13216 25412
rect 11164 25344 11192 25384
rect 8312 25316 11192 25344
rect 11348 25316 11928 25344
rect 7377 25279 7435 25285
rect 7377 25276 7389 25279
rect 7156 25248 7389 25276
rect 7156 25236 7162 25248
rect 7377 25245 7389 25248
rect 7423 25245 7435 25279
rect 7377 25239 7435 25245
rect 7561 25279 7619 25285
rect 7561 25245 7573 25279
rect 7607 25245 7619 25279
rect 7561 25239 7619 25245
rect 7653 25279 7711 25285
rect 7653 25245 7665 25279
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 5040 25180 5488 25208
rect 6089 25211 6147 25217
rect 5040 25168 5046 25180
rect 5276 25152 5304 25180
rect 6089 25177 6101 25211
rect 6135 25208 6147 25211
rect 6825 25211 6883 25217
rect 6135 25180 6500 25208
rect 6135 25177 6147 25180
rect 6089 25171 6147 25177
rect 6472 25152 6500 25180
rect 6825 25177 6837 25211
rect 6871 25177 6883 25211
rect 6825 25171 6883 25177
rect 1544 25112 2912 25140
rect 1544 25100 1550 25112
rect 3418 25100 3424 25152
rect 3476 25100 3482 25152
rect 4062 25100 4068 25152
rect 4120 25140 4126 25152
rect 4433 25143 4491 25149
rect 4433 25140 4445 25143
rect 4120 25112 4445 25140
rect 4120 25100 4126 25112
rect 4433 25109 4445 25112
rect 4479 25140 4491 25143
rect 4890 25140 4896 25152
rect 4479 25112 4896 25140
rect 4479 25109 4491 25112
rect 4433 25103 4491 25109
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 5258 25100 5264 25152
rect 5316 25100 5322 25152
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 6365 25143 6423 25149
rect 6365 25140 6377 25143
rect 5592 25112 6377 25140
rect 5592 25100 5598 25112
rect 6365 25109 6377 25112
rect 6411 25109 6423 25143
rect 6365 25103 6423 25109
rect 6454 25100 6460 25152
rect 6512 25100 6518 25152
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 6840 25140 6868 25171
rect 7668 25152 7696 25239
rect 8202 25236 8208 25288
rect 8260 25276 8266 25288
rect 8312 25285 8340 25316
rect 8297 25279 8355 25285
rect 8297 25276 8309 25279
rect 8260 25248 8309 25276
rect 8260 25236 8266 25248
rect 8297 25245 8309 25248
rect 8343 25245 8355 25279
rect 8297 25239 8355 25245
rect 8481 25279 8539 25285
rect 8481 25245 8493 25279
rect 8527 25276 8539 25279
rect 8570 25276 8576 25288
rect 8527 25248 8576 25276
rect 8527 25245 8539 25248
rect 8481 25239 8539 25245
rect 8570 25236 8576 25248
rect 8628 25236 8634 25288
rect 9140 25285 9168 25316
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 7926 25168 7932 25220
rect 7984 25208 7990 25220
rect 7984 25180 8248 25208
rect 7984 25168 7990 25180
rect 8220 25152 8248 25180
rect 8386 25168 8392 25220
rect 8444 25168 8450 25220
rect 8662 25168 8668 25220
rect 8720 25208 8726 25220
rect 8956 25208 8984 25239
rect 9214 25236 9220 25288
rect 9272 25236 9278 25288
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 9490 25236 9496 25288
rect 9548 25236 9554 25288
rect 9858 25236 9864 25288
rect 9916 25236 9922 25288
rect 10229 25279 10287 25285
rect 10229 25245 10241 25279
rect 10275 25276 10287 25279
rect 10318 25276 10324 25288
rect 10275 25248 10324 25276
rect 10275 25245 10287 25248
rect 10229 25239 10287 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10594 25276 10600 25288
rect 10551 25248 10600 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 9508 25208 9536 25236
rect 8720 25180 9536 25208
rect 8720 25168 8726 25180
rect 6788 25112 6868 25140
rect 7101 25143 7159 25149
rect 6788 25100 6794 25112
rect 7101 25109 7113 25143
rect 7147 25140 7159 25143
rect 7466 25140 7472 25152
rect 7147 25112 7472 25140
rect 7147 25109 7159 25112
rect 7101 25103 7159 25109
rect 7466 25100 7472 25112
rect 7524 25100 7530 25152
rect 7650 25100 7656 25152
rect 7708 25100 7714 25152
rect 8202 25100 8208 25152
rect 8260 25140 8266 25152
rect 9876 25140 9904 25236
rect 10045 25211 10103 25217
rect 10045 25177 10057 25211
rect 10091 25177 10103 25211
rect 10045 25171 10103 25177
rect 8260 25112 9904 25140
rect 10060 25140 10088 25171
rect 10134 25168 10140 25220
rect 10192 25168 10198 25220
rect 10410 25140 10416 25152
rect 10060 25112 10416 25140
rect 8260 25100 8266 25112
rect 10410 25100 10416 25112
rect 10468 25140 10474 25152
rect 10520 25140 10548 25239
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10704 25285 10732 25316
rect 10689 25279 10747 25285
rect 10689 25245 10701 25279
rect 10735 25245 10747 25279
rect 10689 25239 10747 25245
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 11054 25276 11060 25288
rect 10919 25248 11060 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 11146 25236 11152 25288
rect 11204 25236 11210 25288
rect 11348 25285 11376 25316
rect 11333 25279 11391 25285
rect 11333 25245 11345 25279
rect 11379 25245 11391 25279
rect 11333 25239 11391 25245
rect 11425 25279 11483 25285
rect 11425 25245 11437 25279
rect 11471 25276 11483 25279
rect 11514 25276 11520 25288
rect 11471 25248 11520 25276
rect 11471 25245 11483 25248
rect 11425 25239 11483 25245
rect 11514 25236 11520 25248
rect 11572 25236 11578 25288
rect 11606 25236 11612 25288
rect 11664 25236 11670 25288
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 10781 25211 10839 25217
rect 10781 25177 10793 25211
rect 10827 25177 10839 25211
rect 10781 25171 10839 25177
rect 10468 25112 10548 25140
rect 10468 25100 10474 25112
rect 10594 25100 10600 25152
rect 10652 25140 10658 25152
rect 10796 25140 10824 25171
rect 10962 25168 10968 25220
rect 11020 25208 11026 25220
rect 11716 25208 11744 25239
rect 11020 25180 11744 25208
rect 11900 25208 11928 25316
rect 11992 25316 12655 25344
rect 11992 25288 12020 25316
rect 11974 25236 11980 25288
rect 12032 25236 12038 25288
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 12627 25276 12655 25316
rect 12894 25304 12900 25356
rect 12952 25304 12958 25356
rect 13188 25344 13216 25384
rect 14366 25372 14372 25424
rect 14424 25372 14430 25424
rect 15378 25412 15384 25424
rect 15120 25384 15384 25412
rect 13188 25316 14320 25344
rect 13188 25285 13216 25316
rect 14292 25288 14320 25316
rect 13173 25279 13231 25285
rect 12627 25248 13124 25276
rect 13096 25208 13124 25248
rect 13173 25245 13185 25279
rect 13219 25245 13231 25279
rect 13173 25239 13231 25245
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25276 13507 25279
rect 13722 25276 13728 25288
rect 13495 25248 13728 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 13722 25236 13728 25248
rect 13780 25236 13786 25288
rect 13817 25279 13875 25285
rect 13817 25245 13829 25279
rect 13863 25245 13875 25279
rect 13817 25239 13875 25245
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25276 14151 25279
rect 14182 25276 14188 25288
rect 14139 25248 14188 25276
rect 14139 25245 14151 25248
rect 14093 25239 14151 25245
rect 13538 25208 13544 25220
rect 11900 25180 12940 25208
rect 13096 25180 13544 25208
rect 11020 25168 11026 25180
rect 10652 25112 10824 25140
rect 10652 25100 10658 25112
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11900 25140 11928 25180
rect 12912 25152 12940 25180
rect 13538 25168 13544 25180
rect 13596 25208 13602 25220
rect 13832 25208 13860 25239
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14384 25285 14412 25372
rect 14660 25316 15056 25344
rect 14660 25288 14688 25316
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14642 25236 14648 25288
rect 14700 25236 14706 25288
rect 15028 25285 15056 25316
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 15013 25279 15071 25285
rect 15013 25245 15025 25279
rect 15059 25245 15071 25279
rect 15013 25239 15071 25245
rect 13998 25208 14004 25220
rect 13596 25180 14004 25208
rect 13596 25168 13602 25180
rect 13998 25168 14004 25180
rect 14056 25208 14062 25220
rect 14476 25208 14504 25236
rect 14056 25180 14504 25208
rect 14056 25168 14062 25180
rect 14734 25168 14740 25220
rect 14792 25208 14798 25220
rect 14844 25208 14872 25239
rect 15120 25208 15148 25384
rect 15378 25372 15384 25384
rect 15436 25372 15442 25424
rect 15488 25344 15516 25443
rect 16206 25440 16212 25452
rect 16264 25440 16270 25492
rect 16298 25440 16304 25492
rect 16356 25440 16362 25492
rect 16574 25440 16580 25492
rect 16632 25440 16638 25492
rect 17126 25440 17132 25492
rect 17184 25480 17190 25492
rect 17494 25480 17500 25492
rect 17184 25452 17500 25480
rect 17184 25440 17190 25452
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 17770 25440 17776 25492
rect 17828 25480 17834 25492
rect 17957 25483 18015 25489
rect 17957 25480 17969 25483
rect 17828 25452 17969 25480
rect 17828 25440 17834 25452
rect 17957 25449 17969 25452
rect 18003 25480 18015 25483
rect 18414 25480 18420 25492
rect 18003 25452 18420 25480
rect 18003 25449 18015 25452
rect 17957 25443 18015 25449
rect 18414 25440 18420 25452
rect 18472 25440 18478 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 19613 25483 19671 25489
rect 19613 25480 19625 25483
rect 19576 25452 19625 25480
rect 19576 25440 19582 25452
rect 19613 25449 19625 25452
rect 19659 25449 19671 25483
rect 19613 25443 19671 25449
rect 16022 25344 16028 25356
rect 15488 25316 16028 25344
rect 16022 25304 16028 25316
rect 16080 25304 16086 25356
rect 16316 25344 16344 25440
rect 16850 25372 16856 25424
rect 16908 25412 16914 25424
rect 17681 25415 17739 25421
rect 17681 25412 17693 25415
rect 16908 25384 17693 25412
rect 16908 25372 16914 25384
rect 17681 25381 17693 25384
rect 17727 25381 17739 25415
rect 17681 25375 17739 25381
rect 16316 25316 16528 25344
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 15749 25279 15807 25285
rect 15749 25276 15761 25279
rect 15344 25248 15761 25276
rect 15344 25236 15350 25248
rect 15749 25245 15761 25248
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 14792 25180 15148 25208
rect 15764 25208 15792 25239
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 15988 25248 16221 25276
rect 15988 25236 15994 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 16298 25236 16304 25288
rect 16356 25236 16362 25288
rect 16500 25285 16528 25316
rect 16666 25304 16672 25356
rect 16724 25304 16730 25356
rect 17494 25344 17500 25356
rect 16776 25316 17500 25344
rect 16776 25285 16804 25316
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 17696 25344 17724 25375
rect 18230 25372 18236 25424
rect 18288 25412 18294 25424
rect 18966 25412 18972 25424
rect 18288 25384 18972 25412
rect 18288 25372 18294 25384
rect 18966 25372 18972 25384
rect 19024 25412 19030 25424
rect 19024 25384 19564 25412
rect 19024 25372 19030 25384
rect 17696 25316 18460 25344
rect 16393 25279 16451 25285
rect 16393 25245 16405 25279
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 16485 25279 16543 25285
rect 16485 25245 16497 25279
rect 16531 25245 16543 25279
rect 16485 25239 16543 25245
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 16316 25208 16344 25236
rect 15764 25180 16344 25208
rect 16408 25208 16436 25239
rect 17402 25236 17408 25288
rect 17460 25276 17466 25288
rect 18432 25285 18460 25316
rect 17865 25279 17923 25285
rect 17865 25276 17877 25279
rect 17460 25248 17877 25276
rect 17460 25236 17466 25248
rect 17865 25245 17877 25248
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18506 25236 18512 25288
rect 18564 25276 18570 25288
rect 19334 25276 19340 25288
rect 18564 25248 19340 25276
rect 18564 25236 18570 25248
rect 19334 25236 19340 25248
rect 19392 25236 19398 25288
rect 19536 25276 19564 25384
rect 19628 25344 19656 25443
rect 20162 25440 20168 25492
rect 20220 25440 20226 25492
rect 20346 25440 20352 25492
rect 20404 25440 20410 25492
rect 20530 25440 20536 25492
rect 20588 25480 20594 25492
rect 20588 25452 21220 25480
rect 20588 25440 20594 25452
rect 19886 25372 19892 25424
rect 19944 25412 19950 25424
rect 20364 25412 20392 25440
rect 19944 25384 20392 25412
rect 20441 25415 20499 25421
rect 19944 25372 19950 25384
rect 20441 25381 20453 25415
rect 20487 25412 20499 25415
rect 21192 25412 21220 25452
rect 21266 25440 21272 25492
rect 21324 25440 21330 25492
rect 21637 25483 21695 25489
rect 21637 25449 21649 25483
rect 21683 25480 21695 25483
rect 22002 25480 22008 25492
rect 21683 25452 22008 25480
rect 21683 25449 21695 25452
rect 21637 25443 21695 25449
rect 22002 25440 22008 25452
rect 22060 25440 22066 25492
rect 22922 25440 22928 25492
rect 22980 25440 22986 25492
rect 24670 25480 24676 25492
rect 23768 25452 24676 25480
rect 21913 25415 21971 25421
rect 21913 25412 21925 25415
rect 20487 25384 20852 25412
rect 21192 25384 21925 25412
rect 20487 25381 20499 25384
rect 20441 25375 20499 25381
rect 19628 25316 20760 25344
rect 19978 25276 19984 25288
rect 19536 25248 19984 25276
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 20073 25279 20131 25285
rect 20073 25245 20085 25279
rect 20119 25276 20131 25279
rect 20162 25276 20168 25288
rect 20119 25248 20168 25276
rect 20119 25245 20131 25248
rect 20073 25239 20131 25245
rect 20162 25236 20168 25248
rect 20220 25236 20226 25288
rect 20349 25279 20407 25285
rect 20349 25245 20361 25279
rect 20395 25245 20407 25279
rect 20349 25239 20407 25245
rect 17034 25208 17040 25220
rect 16408 25180 17040 25208
rect 14792 25168 14798 25180
rect 17034 25168 17040 25180
rect 17092 25168 17098 25220
rect 17129 25211 17187 25217
rect 17129 25177 17141 25211
rect 17175 25208 17187 25211
rect 17175 25180 17356 25208
rect 17175 25177 17187 25180
rect 17129 25171 17187 25177
rect 17328 25152 17356 25180
rect 17586 25168 17592 25220
rect 17644 25208 17650 25220
rect 20364 25208 20392 25239
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 20533 25279 20591 25285
rect 20533 25276 20545 25279
rect 20496 25248 20545 25276
rect 20496 25236 20502 25248
rect 20533 25245 20545 25248
rect 20579 25245 20591 25279
rect 20533 25239 20591 25245
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20732 25276 20760 25316
rect 20824 25288 20852 25384
rect 21913 25381 21925 25384
rect 21959 25381 21971 25415
rect 21913 25375 21971 25381
rect 23014 25372 23020 25424
rect 23072 25412 23078 25424
rect 23293 25415 23351 25421
rect 23293 25412 23305 25415
rect 23072 25384 23305 25412
rect 23072 25372 23078 25384
rect 23293 25381 23305 25384
rect 23339 25412 23351 25415
rect 23768 25412 23796 25452
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 25130 25440 25136 25492
rect 25188 25480 25194 25492
rect 28629 25483 28687 25489
rect 28629 25480 28641 25483
rect 25188 25452 28641 25480
rect 25188 25440 25194 25452
rect 28629 25449 28641 25452
rect 28675 25449 28687 25483
rect 28629 25443 28687 25449
rect 28966 25452 29592 25480
rect 23339 25384 23796 25412
rect 23339 25381 23351 25384
rect 23293 25375 23351 25381
rect 22830 25304 22836 25356
rect 22888 25344 22894 25356
rect 22888 25316 23428 25344
rect 22888 25304 22894 25316
rect 20671 25248 20760 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20806 25236 20812 25288
rect 20864 25236 20870 25288
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 21085 25279 21143 25285
rect 21085 25276 21097 25279
rect 21048 25248 21097 25276
rect 21048 25236 21054 25248
rect 21085 25245 21097 25248
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25276 21603 25279
rect 21634 25276 21640 25288
rect 21591 25248 21640 25276
rect 21591 25245 21603 25248
rect 21545 25239 21603 25245
rect 21634 25236 21640 25248
rect 21692 25236 21698 25288
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 21729 25239 21787 25245
rect 20714 25208 20720 25220
rect 17644 25180 19334 25208
rect 20364 25180 20720 25208
rect 17644 25168 17650 25180
rect 11204 25112 11928 25140
rect 11204 25100 11210 25112
rect 12894 25100 12900 25152
rect 12952 25140 12958 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 12952 25112 14841 25140
rect 12952 25100 12958 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 14829 25103 14887 25109
rect 15378 25100 15384 25152
rect 15436 25140 15442 25152
rect 15565 25143 15623 25149
rect 15565 25140 15577 25143
rect 15436 25112 15577 25140
rect 15436 25100 15442 25112
rect 15565 25109 15577 25112
rect 15611 25109 15623 25143
rect 15565 25103 15623 25109
rect 15838 25100 15844 25152
rect 15896 25140 15902 25152
rect 16758 25140 16764 25152
rect 15896 25112 16764 25140
rect 15896 25100 15902 25112
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 16942 25100 16948 25152
rect 17000 25100 17006 25152
rect 17310 25100 17316 25152
rect 17368 25100 17374 25152
rect 17494 25100 17500 25152
rect 17552 25149 17558 25152
rect 17552 25140 17564 25149
rect 19306 25140 19334 25180
rect 20714 25168 20720 25180
rect 20772 25168 20778 25220
rect 20901 25211 20959 25217
rect 20901 25177 20913 25211
rect 20947 25208 20959 25211
rect 21450 25208 21456 25220
rect 20947 25180 21456 25208
rect 20947 25177 20959 25180
rect 20901 25171 20959 25177
rect 21450 25168 21456 25180
rect 21508 25168 21514 25220
rect 19794 25140 19800 25152
rect 17552 25112 17597 25140
rect 19306 25112 19800 25140
rect 17552 25103 17564 25112
rect 17552 25100 17558 25103
rect 19794 25100 19800 25112
rect 19852 25100 19858 25152
rect 20070 25100 20076 25152
rect 20128 25140 20134 25152
rect 21744 25140 21772 25239
rect 22094 25236 22100 25288
rect 22152 25236 22158 25288
rect 22186 25236 22192 25288
rect 22244 25236 22250 25288
rect 22370 25236 22376 25288
rect 22428 25236 22434 25288
rect 22462 25236 22468 25288
rect 22520 25236 22526 25288
rect 23109 25279 23167 25285
rect 23109 25245 23121 25279
rect 23155 25245 23167 25279
rect 23109 25239 23167 25245
rect 23124 25208 23152 25239
rect 23198 25236 23204 25288
rect 23256 25236 23262 25288
rect 23400 25285 23428 25316
rect 23768 25285 23796 25384
rect 24397 25415 24455 25421
rect 24397 25381 24409 25415
rect 24443 25381 24455 25415
rect 24397 25375 24455 25381
rect 24412 25344 24440 25375
rect 24486 25372 24492 25424
rect 24544 25412 24550 25424
rect 25406 25412 25412 25424
rect 24544 25384 25412 25412
rect 24544 25372 24550 25384
rect 25406 25372 25412 25384
rect 25464 25372 25470 25424
rect 27617 25415 27675 25421
rect 27617 25381 27629 25415
rect 27663 25412 27675 25415
rect 28966 25412 28994 25452
rect 29564 25424 29592 25452
rect 29638 25440 29644 25492
rect 29696 25440 29702 25492
rect 31110 25440 31116 25492
rect 31168 25480 31174 25492
rect 32309 25483 32367 25489
rect 32309 25480 32321 25483
rect 31168 25452 32321 25480
rect 31168 25440 31174 25452
rect 32309 25449 32321 25452
rect 32355 25449 32367 25483
rect 32309 25443 32367 25449
rect 32490 25440 32496 25492
rect 32548 25440 32554 25492
rect 32950 25440 32956 25492
rect 33008 25480 33014 25492
rect 33505 25483 33563 25489
rect 33505 25480 33517 25483
rect 33008 25452 33517 25480
rect 33008 25440 33014 25452
rect 33505 25449 33517 25452
rect 33551 25480 33563 25483
rect 43254 25480 43260 25492
rect 33551 25452 43260 25480
rect 33551 25449 33563 25452
rect 33505 25443 33563 25449
rect 43254 25440 43260 25452
rect 43312 25440 43318 25492
rect 27663 25384 28994 25412
rect 27663 25381 27675 25384
rect 27617 25375 27675 25381
rect 29454 25372 29460 25424
rect 29512 25372 29518 25424
rect 29546 25372 29552 25424
rect 29604 25372 29610 25424
rect 31573 25415 31631 25421
rect 31573 25381 31585 25415
rect 31619 25381 31631 25415
rect 31573 25375 31631 25381
rect 24412 25316 24808 25344
rect 23374 25279 23432 25285
rect 23374 25245 23386 25279
rect 23420 25245 23432 25279
rect 23374 25239 23432 25245
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 23934 25276 23940 25288
rect 23891 25248 23940 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 24026 25236 24032 25288
rect 24084 25236 24090 25288
rect 24121 25279 24179 25285
rect 24121 25245 24133 25279
rect 24167 25276 24179 25279
rect 24167 25248 24532 25276
rect 24167 25245 24179 25248
rect 24121 25239 24179 25245
rect 23124 25180 23336 25208
rect 23308 25152 23336 25180
rect 20128 25112 21772 25140
rect 20128 25100 20134 25112
rect 22094 25100 22100 25152
rect 22152 25140 22158 25152
rect 22830 25140 22836 25152
rect 22152 25112 22836 25140
rect 22152 25100 22158 25112
rect 22830 25100 22836 25112
rect 22888 25100 22894 25152
rect 23290 25100 23296 25152
rect 23348 25100 23354 25152
rect 23566 25100 23572 25152
rect 23624 25100 23630 25152
rect 23952 25140 23980 25236
rect 24394 25168 24400 25220
rect 24452 25168 24458 25220
rect 24504 25208 24532 25248
rect 24578 25236 24584 25288
rect 24636 25276 24642 25288
rect 24780 25285 24808 25316
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 24912 25316 24992 25344
rect 24912 25304 24918 25316
rect 24964 25285 24992 25316
rect 26510 25304 26516 25356
rect 26568 25344 26574 25356
rect 26973 25347 27031 25353
rect 26973 25344 26985 25347
rect 26568 25316 26985 25344
rect 26568 25304 26574 25316
rect 26973 25313 26985 25316
rect 27019 25313 27031 25347
rect 26973 25307 27031 25313
rect 27982 25304 27988 25356
rect 28040 25304 28046 25356
rect 28902 25304 28908 25356
rect 28960 25344 28966 25356
rect 29472 25344 29500 25372
rect 30193 25347 30251 25353
rect 30193 25344 30205 25347
rect 28960 25316 29040 25344
rect 29472 25316 30205 25344
rect 28960 25304 28966 25316
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24636 25248 24685 25276
rect 24636 25236 24642 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25245 24823 25279
rect 24765 25239 24823 25245
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 25065 25279 25123 25285
rect 25065 25245 25077 25279
rect 25111 25276 25123 25279
rect 25111 25248 25360 25276
rect 25111 25245 25123 25248
rect 25065 25239 25123 25245
rect 25332 25220 25360 25248
rect 26694 25236 26700 25288
rect 26752 25236 26758 25288
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 27338 25276 27344 25288
rect 26927 25248 27344 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 27338 25236 27344 25248
rect 27396 25236 27402 25288
rect 29012 25285 29040 25316
rect 30193 25313 30205 25316
rect 30239 25313 30251 25347
rect 31588 25344 31616 25375
rect 31665 25347 31723 25353
rect 31665 25344 31677 25347
rect 31588 25316 31677 25344
rect 30193 25307 30251 25313
rect 31665 25313 31677 25316
rect 31711 25313 31723 25347
rect 31665 25307 31723 25313
rect 32674 25304 32680 25356
rect 32732 25304 32738 25356
rect 28997 25279 29055 25285
rect 28997 25276 29009 25279
rect 27448 25248 29009 25276
rect 24857 25211 24915 25217
rect 24857 25208 24869 25211
rect 24504 25180 24869 25208
rect 24857 25177 24869 25180
rect 24903 25177 24915 25211
rect 24857 25171 24915 25177
rect 25314 25168 25320 25220
rect 25372 25208 25378 25220
rect 27448 25208 27476 25248
rect 28997 25245 29009 25248
rect 29043 25245 29055 25279
rect 29089 25276 29147 25282
rect 29089 25266 29101 25276
rect 29135 25266 29147 25276
rect 29181 25279 29239 25285
rect 28997 25239 29055 25245
rect 25372 25180 27476 25208
rect 28721 25211 28779 25217
rect 29086 25214 29092 25266
rect 29144 25214 29150 25266
rect 29181 25245 29193 25279
rect 29227 25276 29239 25279
rect 29270 25276 29276 25288
rect 29227 25248 29276 25276
rect 29227 25245 29239 25248
rect 29181 25239 29239 25245
rect 29270 25236 29276 25248
rect 29328 25236 29334 25288
rect 29377 25279 29435 25285
rect 29377 25245 29389 25279
rect 29423 25276 29435 25279
rect 29549 25279 29607 25285
rect 29423 25248 29500 25276
rect 29423 25245 29435 25248
rect 29377 25239 29435 25245
rect 25372 25168 25378 25180
rect 28721 25177 28733 25211
rect 28767 25208 28779 25211
rect 29472 25208 29500 25248
rect 29549 25245 29561 25279
rect 29595 25276 29607 25279
rect 29730 25276 29736 25288
rect 29595 25248 29736 25276
rect 29595 25245 29607 25248
rect 29549 25239 29607 25245
rect 29730 25236 29736 25248
rect 29788 25236 29794 25288
rect 30006 25236 30012 25288
rect 30064 25276 30070 25288
rect 31570 25276 31576 25288
rect 30064 25248 31576 25276
rect 30064 25236 30070 25248
rect 31570 25236 31576 25248
rect 31628 25236 31634 25288
rect 32401 25279 32459 25285
rect 32401 25276 32413 25279
rect 31772 25248 32413 25276
rect 30190 25208 30196 25220
rect 28767 25180 29040 25208
rect 29472 25180 30196 25208
rect 28767 25177 28779 25180
rect 28721 25171 28779 25177
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 23952 25112 24593 25140
rect 24581 25109 24593 25112
rect 24627 25140 24639 25143
rect 25133 25143 25191 25149
rect 25133 25140 25145 25143
rect 24627 25112 25145 25140
rect 24627 25109 24639 25112
rect 24581 25103 24639 25109
rect 25133 25109 25145 25112
rect 25179 25109 25191 25143
rect 25133 25103 25191 25109
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25140 26847 25143
rect 27246 25140 27252 25152
rect 26835 25112 27252 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 27246 25100 27252 25112
rect 27304 25100 27310 25152
rect 29012 25140 29040 25180
rect 30190 25168 30196 25180
rect 30248 25168 30254 25220
rect 30460 25211 30518 25217
rect 30460 25177 30472 25211
rect 30506 25208 30518 25211
rect 30558 25208 30564 25220
rect 30506 25180 30564 25208
rect 30506 25177 30518 25180
rect 30460 25171 30518 25177
rect 30558 25168 30564 25180
rect 30616 25168 30622 25220
rect 31772 25152 31800 25248
rect 32401 25245 32413 25248
rect 32447 25276 32459 25279
rect 32953 25279 33011 25285
rect 32953 25276 32965 25279
rect 32447 25248 32965 25276
rect 32447 25245 32459 25248
rect 32401 25239 32459 25245
rect 32953 25245 32965 25248
rect 32999 25245 33011 25279
rect 32953 25239 33011 25245
rect 29086 25140 29092 25152
rect 29012 25112 29092 25140
rect 29086 25100 29092 25112
rect 29144 25100 29150 25152
rect 31754 25100 31760 25152
rect 31812 25100 31818 25152
rect 32214 25100 32220 25152
rect 32272 25140 32278 25152
rect 32677 25143 32735 25149
rect 32677 25140 32689 25143
rect 32272 25112 32689 25140
rect 32272 25100 32278 25112
rect 32677 25109 32689 25112
rect 32723 25109 32735 25143
rect 32677 25103 32735 25109
rect 1104 25050 43884 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 43884 25050
rect 1104 24976 43884 24998
rect 1762 24896 1768 24948
rect 1820 24896 1826 24948
rect 5166 24896 5172 24948
rect 5224 24896 5230 24948
rect 5350 24896 5356 24948
rect 5408 24896 5414 24948
rect 5442 24896 5448 24948
rect 5500 24936 5506 24948
rect 6730 24936 6736 24948
rect 5500 24908 6736 24936
rect 5500 24896 5506 24908
rect 6730 24896 6736 24908
rect 6788 24896 6794 24948
rect 8389 24939 8447 24945
rect 8389 24905 8401 24939
rect 8435 24936 8447 24939
rect 8662 24936 8668 24948
rect 8435 24908 8668 24936
rect 8435 24905 8447 24908
rect 8389 24899 8447 24905
rect 8662 24896 8668 24908
rect 8720 24896 8726 24948
rect 9030 24896 9036 24948
rect 9088 24896 9094 24948
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 10689 24939 10747 24945
rect 9916 24908 10456 24936
rect 9916 24896 9922 24908
rect 2038 24828 2044 24880
rect 2096 24868 2102 24880
rect 5074 24868 5080 24880
rect 2096 24840 2636 24868
rect 2096 24828 2102 24840
rect 2608 24809 2636 24840
rect 2700 24840 5080 24868
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 2501 24803 2559 24809
rect 2501 24800 2513 24803
rect 1627 24772 2513 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 2501 24769 2513 24772
rect 2547 24769 2559 24803
rect 2501 24763 2559 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24769 2651 24803
rect 2593 24763 2651 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1486 24732 1492 24744
rect 1443 24704 1492 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1486 24692 1492 24704
rect 1544 24692 1550 24744
rect 1949 24735 2007 24741
rect 1949 24701 1961 24735
rect 1995 24732 2007 24735
rect 2700 24732 2728 24840
rect 5074 24828 5080 24840
rect 5132 24828 5138 24880
rect 5184 24868 5212 24896
rect 5184 24840 5393 24868
rect 2860 24803 2918 24809
rect 2860 24769 2872 24803
rect 2906 24800 2918 24803
rect 3602 24800 3608 24812
rect 2906 24772 3608 24800
rect 2906 24769 2918 24772
rect 2860 24763 2918 24769
rect 3602 24760 3608 24772
rect 3660 24760 3666 24812
rect 3694 24760 3700 24812
rect 3752 24800 3758 24812
rect 4614 24800 4620 24812
rect 3752 24772 4620 24800
rect 3752 24760 3758 24772
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 4798 24760 4804 24812
rect 4856 24760 4862 24812
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24769 5043 24803
rect 4985 24763 5043 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5258 24800 5264 24812
rect 5215 24772 5264 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 4065 24735 4123 24741
rect 4065 24732 4077 24735
rect 1995 24704 2544 24732
rect 1995 24701 2007 24704
rect 1949 24695 2007 24701
rect 2516 24596 2544 24704
rect 2608 24704 2728 24732
rect 3988 24704 4077 24732
rect 2608 24676 2636 24704
rect 2590 24624 2596 24676
rect 2648 24624 2654 24676
rect 3988 24673 4016 24704
rect 4065 24701 4077 24704
rect 4111 24732 4123 24735
rect 4522 24732 4528 24744
rect 4111 24704 4528 24732
rect 4111 24701 4123 24704
rect 4065 24695 4123 24701
rect 4522 24692 4528 24704
rect 4580 24692 4586 24744
rect 3973 24667 4031 24673
rect 3973 24633 3985 24667
rect 4019 24633 4031 24667
rect 4816 24664 4844 24760
rect 5000 24732 5028 24763
rect 5258 24760 5264 24772
rect 5316 24760 5322 24812
rect 5365 24732 5393 24840
rect 5902 24828 5908 24880
rect 5960 24828 5966 24880
rect 6914 24868 6920 24880
rect 6058 24840 6920 24868
rect 5534 24760 5540 24812
rect 5592 24760 5598 24812
rect 6058 24809 6086 24840
rect 6914 24828 6920 24840
rect 6972 24868 6978 24880
rect 7285 24871 7343 24877
rect 7285 24868 7297 24871
rect 6972 24840 7297 24868
rect 6972 24828 6978 24840
rect 7285 24837 7297 24840
rect 7331 24868 7343 24871
rect 7650 24868 7656 24880
rect 7331 24840 7656 24868
rect 7331 24837 7343 24840
rect 7285 24831 7343 24837
rect 7650 24828 7656 24840
rect 7708 24868 7714 24880
rect 7708 24840 8064 24868
rect 7708 24828 7714 24840
rect 5685 24803 5743 24809
rect 5685 24769 5697 24803
rect 5731 24769 5743 24803
rect 5685 24763 5743 24769
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6043 24803 6101 24809
rect 5859 24772 5948 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 5000 24704 5393 24732
rect 5700 24732 5728 24763
rect 5920 24744 5948 24772
rect 6043 24769 6055 24803
rect 6089 24769 6101 24803
rect 6043 24763 6101 24769
rect 6270 24760 6276 24812
rect 6328 24760 6334 24812
rect 6365 24803 6423 24809
rect 6365 24769 6377 24803
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 5700 24704 5764 24732
rect 5534 24664 5540 24676
rect 4816 24636 5540 24664
rect 3973 24627 4031 24633
rect 5534 24624 5540 24636
rect 5592 24624 5598 24676
rect 5736 24664 5764 24704
rect 5902 24692 5908 24744
rect 5960 24692 5966 24744
rect 6288 24664 6316 24760
rect 5736 24636 6316 24664
rect 6380 24664 6408 24763
rect 6546 24760 6552 24812
rect 6604 24760 6610 24812
rect 6638 24760 6644 24812
rect 6696 24760 6702 24812
rect 6730 24760 6736 24812
rect 6788 24760 6794 24812
rect 7006 24760 7012 24812
rect 7064 24760 7070 24812
rect 7190 24809 7196 24812
rect 7157 24803 7196 24809
rect 7157 24769 7169 24803
rect 7157 24763 7196 24769
rect 7190 24760 7196 24763
rect 7248 24760 7254 24812
rect 7377 24803 7435 24809
rect 7377 24769 7389 24803
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 7515 24803 7573 24809
rect 7515 24769 7527 24803
rect 7561 24800 7573 24803
rect 7926 24800 7932 24812
rect 7561 24772 7932 24800
rect 7561 24769 7573 24772
rect 7515 24763 7573 24769
rect 7392 24732 7420 24763
rect 7926 24760 7932 24772
rect 7984 24760 7990 24812
rect 7742 24732 7748 24744
rect 7392 24704 7748 24732
rect 7742 24692 7748 24704
rect 7800 24692 7806 24744
rect 8036 24732 8064 24840
rect 8202 24760 8208 24812
rect 8260 24800 8266 24812
rect 8680 24809 8708 24896
rect 9401 24871 9459 24877
rect 9401 24837 9413 24871
rect 9447 24868 9459 24871
rect 9674 24868 9680 24880
rect 9447 24840 9680 24868
rect 9447 24837 9459 24840
rect 9401 24831 9459 24837
rect 9674 24828 9680 24840
rect 9732 24868 9738 24880
rect 10321 24871 10379 24877
rect 10321 24868 10333 24871
rect 9732 24840 10333 24868
rect 9732 24828 9738 24840
rect 10321 24837 10333 24840
rect 10367 24837 10379 24871
rect 10428 24868 10456 24908
rect 10689 24905 10701 24939
rect 10735 24936 10747 24939
rect 10962 24936 10968 24948
rect 10735 24908 10968 24936
rect 10735 24905 10747 24908
rect 10689 24899 10747 24905
rect 10962 24896 10968 24908
rect 11020 24896 11026 24948
rect 11238 24896 11244 24948
rect 11296 24896 11302 24948
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 12066 24936 12072 24948
rect 11756 24908 12072 24936
rect 11756 24896 11762 24908
rect 12066 24896 12072 24908
rect 12124 24936 12130 24948
rect 12618 24936 12624 24948
rect 12124 24908 12624 24936
rect 12124 24896 12130 24908
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 13449 24939 13507 24945
rect 13449 24905 13461 24939
rect 13495 24936 13507 24939
rect 13630 24936 13636 24948
rect 13495 24908 13636 24936
rect 13495 24905 13507 24908
rect 13449 24899 13507 24905
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 14274 24896 14280 24948
rect 14332 24936 14338 24948
rect 15930 24936 15936 24948
rect 14332 24908 15936 24936
rect 14332 24896 14338 24908
rect 15930 24896 15936 24908
rect 15988 24896 15994 24948
rect 16206 24936 16212 24948
rect 16040 24908 16212 24936
rect 11256 24868 11284 24896
rect 13081 24871 13139 24877
rect 10428 24840 11008 24868
rect 10321 24831 10379 24837
rect 10980 24812 11008 24840
rect 11072 24840 11284 24868
rect 11532 24840 12204 24868
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8260 24772 8493 24800
rect 8260 24760 8266 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24769 8723 24803
rect 8665 24763 8723 24769
rect 8754 24760 8760 24812
rect 8812 24760 8818 24812
rect 8849 24803 8907 24809
rect 8849 24769 8861 24803
rect 8895 24800 8907 24803
rect 9030 24800 9036 24812
rect 8895 24772 9036 24800
rect 8895 24769 8907 24772
rect 8849 24763 8907 24769
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 9122 24760 9128 24812
rect 9180 24760 9186 24812
rect 9306 24809 9312 24812
rect 9263 24803 9312 24809
rect 9263 24769 9275 24803
rect 9309 24769 9312 24803
rect 9263 24763 9312 24769
rect 9306 24760 9312 24763
rect 9364 24760 9370 24812
rect 9490 24760 9496 24812
rect 9548 24760 9554 24812
rect 9590 24803 9648 24809
rect 9590 24769 9602 24803
rect 9636 24800 9648 24803
rect 9858 24800 9864 24812
rect 9636 24772 9864 24800
rect 9636 24769 9648 24772
rect 9590 24763 9648 24769
rect 9605 24732 9633 24763
rect 9858 24760 9864 24772
rect 9916 24760 9922 24812
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10137 24763 10195 24769
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10870 24800 10876 24812
rect 10551 24772 10876 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 8036 24704 9633 24732
rect 8021 24667 8079 24673
rect 8021 24664 8033 24667
rect 6380 24636 8033 24664
rect 8021 24633 8033 24636
rect 8067 24664 8079 24667
rect 10152 24664 10180 24763
rect 10428 24732 10456 24763
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 10962 24760 10968 24812
rect 11020 24760 11026 24812
rect 11072 24809 11100 24840
rect 11057 24803 11115 24809
rect 11057 24769 11069 24803
rect 11103 24769 11115 24803
rect 11057 24763 11115 24769
rect 11241 24803 11299 24809
rect 11241 24769 11253 24803
rect 11287 24769 11299 24803
rect 11241 24763 11299 24769
rect 11146 24732 11152 24744
rect 10428 24704 11152 24732
rect 11146 24692 11152 24704
rect 11204 24692 11210 24744
rect 11256 24732 11284 24763
rect 11330 24760 11336 24812
rect 11388 24760 11394 24812
rect 11532 24732 11560 24840
rect 11609 24803 11667 24809
rect 11609 24769 11621 24803
rect 11655 24800 11667 24803
rect 11698 24800 11704 24812
rect 11655 24772 11704 24800
rect 11655 24769 11667 24772
rect 11609 24763 11667 24769
rect 11698 24760 11704 24772
rect 11756 24760 11762 24812
rect 11793 24803 11851 24809
rect 11793 24769 11805 24803
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 11256 24704 11560 24732
rect 11808 24732 11836 24763
rect 11882 24760 11888 24812
rect 11940 24760 11946 24812
rect 11974 24760 11980 24812
rect 12032 24760 12038 24812
rect 11808 24704 11928 24732
rect 10502 24664 10508 24676
rect 8067 24636 9904 24664
rect 10152 24636 10508 24664
rect 8067 24633 8079 24636
rect 8021 24627 8079 24633
rect 9876 24608 9904 24636
rect 10502 24624 10508 24636
rect 10560 24624 10566 24676
rect 11900 24608 11928 24704
rect 12176 24673 12204 24840
rect 13081 24837 13093 24871
rect 13127 24868 13139 24871
rect 14182 24868 14188 24880
rect 13127 24840 14188 24868
rect 13127 24837 13139 24840
rect 13081 24831 13139 24837
rect 14182 24828 14188 24840
rect 14240 24828 14246 24880
rect 15378 24828 15384 24880
rect 15436 24868 15442 24880
rect 16040 24877 16068 24908
rect 16206 24896 16212 24908
rect 16264 24896 16270 24948
rect 16298 24896 16304 24948
rect 16356 24896 16362 24948
rect 19242 24936 19248 24948
rect 16408 24908 19248 24936
rect 16025 24871 16083 24877
rect 15436 24840 15884 24868
rect 15436 24828 15442 24840
rect 12250 24760 12256 24812
rect 12308 24800 12314 24812
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12308 24772 12909 24800
rect 12308 24760 12314 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 12897 24763 12955 24769
rect 12912 24732 12940 24763
rect 13170 24760 13176 24812
rect 13228 24760 13234 24812
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24800 13323 24803
rect 13446 24800 13452 24812
rect 13311 24772 13452 24800
rect 13311 24769 13323 24772
rect 13265 24763 13323 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13538 24760 13544 24812
rect 13596 24760 13602 24812
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 14458 24800 14464 24812
rect 13964 24772 14464 24800
rect 13964 24760 13970 24772
rect 14458 24760 14464 24772
rect 14516 24760 14522 24812
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24800 15347 24803
rect 15335 24772 15424 24800
rect 15335 24769 15347 24772
rect 15289 24763 15347 24769
rect 14001 24735 14059 24741
rect 14001 24732 14013 24735
rect 12912 24704 14013 24732
rect 14001 24701 14013 24704
rect 14047 24701 14059 24735
rect 14001 24695 14059 24701
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 14369 24735 14427 24741
rect 14369 24732 14381 24735
rect 14332 24704 14381 24732
rect 14332 24692 14338 24704
rect 14369 24701 14381 24704
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 12161 24667 12219 24673
rect 12161 24633 12173 24667
rect 12207 24633 12219 24667
rect 12161 24627 12219 24633
rect 14182 24624 14188 24676
rect 14240 24664 14246 24676
rect 14645 24667 14703 24673
rect 14645 24664 14657 24667
rect 14240 24636 14657 24664
rect 14240 24624 14246 24636
rect 14645 24633 14657 24636
rect 14691 24633 14703 24667
rect 14645 24627 14703 24633
rect 15286 24624 15292 24676
rect 15344 24664 15350 24676
rect 15396 24664 15424 24772
rect 15562 24760 15568 24812
rect 15620 24760 15626 24812
rect 15856 24798 15884 24840
rect 16025 24837 16037 24871
rect 16071 24837 16083 24871
rect 16316 24868 16344 24896
rect 16408 24880 16436 24908
rect 19242 24896 19248 24908
rect 19300 24896 19306 24948
rect 19352 24908 20760 24936
rect 16025 24831 16083 24837
rect 16132 24840 16344 24868
rect 16132 24809 16160 24840
rect 16390 24828 16396 24880
rect 16448 24828 16454 24880
rect 19352 24868 19380 24908
rect 20625 24871 20683 24877
rect 20625 24868 20637 24871
rect 16500 24840 17356 24868
rect 15933 24803 15991 24809
rect 15933 24798 15945 24803
rect 15856 24770 15945 24798
rect 15933 24769 15945 24770
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16117 24763 16175 24769
rect 16255 24803 16313 24809
rect 16255 24769 16267 24803
rect 16301 24800 16313 24803
rect 16500 24800 16528 24840
rect 17328 24812 17356 24840
rect 17788 24840 18368 24868
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16301 24772 16528 24800
rect 16592 24772 16681 24800
rect 16301 24769 16313 24772
rect 16255 24763 16313 24769
rect 16592 24744 16620 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16758 24760 16764 24812
rect 16816 24760 16822 24812
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16908 24772 16957 24800
rect 16908 24760 16914 24772
rect 16945 24769 16957 24772
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17678 24760 17684 24812
rect 17736 24760 17742 24812
rect 16393 24735 16451 24741
rect 16393 24701 16405 24735
rect 16439 24701 16451 24735
rect 16393 24695 16451 24701
rect 16408 24664 16436 24695
rect 16574 24692 16580 24744
rect 16632 24692 16638 24744
rect 16776 24732 16804 24760
rect 17129 24735 17187 24741
rect 17129 24732 17141 24735
rect 16776 24704 17141 24732
rect 17129 24701 17141 24704
rect 17175 24732 17187 24735
rect 17586 24732 17592 24744
rect 17175 24704 17592 24732
rect 17175 24701 17187 24704
rect 17129 24695 17187 24701
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 15344 24636 16436 24664
rect 15344 24624 15350 24636
rect 2866 24596 2872 24608
rect 2516 24568 2872 24596
rect 2866 24556 2872 24568
rect 2924 24556 2930 24608
rect 4706 24556 4712 24608
rect 4764 24556 4770 24608
rect 6181 24599 6239 24605
rect 6181 24565 6193 24599
rect 6227 24596 6239 24599
rect 6270 24596 6276 24608
rect 6227 24568 6276 24596
rect 6227 24565 6239 24568
rect 6181 24559 6239 24565
rect 6270 24556 6276 24568
rect 6328 24556 6334 24608
rect 6914 24556 6920 24608
rect 6972 24556 6978 24608
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 7653 24599 7711 24605
rect 7653 24596 7665 24599
rect 7616 24568 7665 24596
rect 7616 24556 7622 24568
rect 7653 24565 7665 24568
rect 7699 24565 7711 24599
rect 7653 24559 7711 24565
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 9306 24596 9312 24608
rect 7984 24568 9312 24596
rect 7984 24556 7990 24568
rect 9306 24556 9312 24568
rect 9364 24556 9370 24608
rect 9766 24556 9772 24608
rect 9824 24556 9830 24608
rect 9858 24556 9864 24608
rect 9916 24556 9922 24608
rect 10686 24556 10692 24608
rect 10744 24596 10750 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10744 24568 10793 24596
rect 10744 24556 10750 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 11882 24556 11888 24608
rect 11940 24556 11946 24608
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 13446 24596 13452 24608
rect 12860 24568 13452 24596
rect 12860 24556 12866 24568
rect 13446 24556 13452 24568
rect 13504 24556 13510 24608
rect 15746 24556 15752 24608
rect 15804 24556 15810 24608
rect 16408 24596 16436 24636
rect 16758 24624 16764 24676
rect 16816 24624 16822 24676
rect 17788 24664 17816 24840
rect 18340 24812 18368 24840
rect 18984 24840 19380 24868
rect 19435 24840 20637 24868
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 17957 24803 18015 24809
rect 17957 24769 17969 24803
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 16868 24636 17816 24664
rect 16868 24596 16896 24636
rect 16408 24568 16896 24596
rect 17494 24556 17500 24608
rect 17552 24556 17558 24608
rect 17880 24596 17908 24763
rect 17972 24664 18000 24763
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 18322 24760 18328 24812
rect 18380 24760 18386 24812
rect 18782 24760 18788 24812
rect 18840 24760 18846 24812
rect 18248 24732 18276 24760
rect 18598 24732 18604 24744
rect 18248 24704 18604 24732
rect 18598 24692 18604 24704
rect 18656 24732 18662 24744
rect 18984 24732 19012 24840
rect 19242 24760 19248 24812
rect 19300 24800 19306 24812
rect 19435 24800 19463 24840
rect 20625 24837 20637 24840
rect 20671 24837 20683 24871
rect 20732 24868 20760 24908
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 21085 24939 21143 24945
rect 21085 24936 21097 24939
rect 20864 24908 21097 24936
rect 20864 24896 20870 24908
rect 21085 24905 21097 24908
rect 21131 24936 21143 24939
rect 21542 24936 21548 24948
rect 21131 24908 21548 24936
rect 21131 24905 21143 24908
rect 21085 24899 21143 24905
rect 21542 24896 21548 24908
rect 21600 24936 21606 24948
rect 22738 24936 22744 24948
rect 21600 24908 22744 24936
rect 21600 24896 21606 24908
rect 22738 24896 22744 24908
rect 22796 24896 22802 24948
rect 24486 24936 24492 24948
rect 23952 24908 24492 24936
rect 20990 24868 20996 24880
rect 20732 24840 20996 24868
rect 20625 24831 20683 24837
rect 20990 24828 20996 24840
rect 21048 24868 21054 24880
rect 21048 24840 21312 24868
rect 21048 24828 21054 24840
rect 19300 24772 19463 24800
rect 19889 24803 19947 24809
rect 19300 24760 19306 24772
rect 19521 24771 19579 24777
rect 18656 24704 19012 24732
rect 18656 24692 18662 24704
rect 19058 24692 19064 24744
rect 19116 24732 19122 24744
rect 19334 24732 19340 24744
rect 19116 24704 19340 24732
rect 19116 24692 19122 24704
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 19521 24737 19533 24771
rect 19567 24737 19579 24771
rect 19889 24769 19901 24803
rect 19935 24800 19947 24803
rect 20070 24800 20076 24812
rect 19935 24772 20076 24800
rect 19935 24769 19947 24772
rect 19889 24763 19947 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 20257 24806 20315 24809
rect 20346 24806 20352 24812
rect 20257 24803 20352 24806
rect 20257 24769 20269 24803
rect 20303 24778 20352 24803
rect 20303 24769 20315 24778
rect 20257 24763 20315 24769
rect 19521 24731 19579 24737
rect 19679 24735 19737 24741
rect 19426 24664 19432 24676
rect 17972 24636 19432 24664
rect 19426 24624 19432 24636
rect 19484 24624 19490 24676
rect 19536 24664 19564 24731
rect 19679 24701 19691 24735
rect 19725 24732 19737 24735
rect 19794 24732 19800 24744
rect 19725 24704 19800 24732
rect 19725 24701 19737 24704
rect 19679 24695 19737 24701
rect 19794 24692 19800 24704
rect 19852 24692 19858 24744
rect 20180 24732 20208 24763
rect 20346 24760 20352 24778
rect 20404 24760 20410 24812
rect 20530 24760 20536 24812
rect 20588 24760 20594 24812
rect 20806 24760 20812 24812
rect 20864 24760 20870 24812
rect 21284 24809 21312 24840
rect 21358 24828 21364 24880
rect 21416 24868 21422 24880
rect 21818 24868 21824 24880
rect 21416 24840 21824 24868
rect 21416 24828 21422 24840
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24769 21327 24803
rect 21269 24763 21327 24769
rect 20548 24732 20576 24760
rect 21100 24732 21128 24763
rect 21450 24760 21456 24812
rect 21508 24760 21514 24812
rect 21652 24809 21680 24840
rect 21818 24828 21824 24840
rect 21876 24868 21882 24880
rect 22370 24868 22376 24880
rect 21876 24840 22376 24868
rect 21876 24828 21882 24840
rect 22370 24828 22376 24840
rect 22428 24828 22434 24880
rect 23106 24868 23112 24880
rect 22480 24840 23112 24868
rect 21637 24803 21695 24809
rect 21637 24769 21649 24803
rect 21683 24769 21695 24803
rect 21637 24763 21695 24769
rect 21910 24760 21916 24812
rect 21968 24800 21974 24812
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 21968 24772 22017 24800
rect 21968 24760 21974 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22189 24803 22247 24809
rect 22189 24769 22201 24803
rect 22235 24800 22247 24803
rect 22480 24800 22508 24840
rect 23106 24828 23112 24840
rect 23164 24828 23170 24880
rect 23952 24877 23980 24908
rect 24486 24896 24492 24908
rect 24544 24896 24550 24948
rect 24578 24896 24584 24948
rect 24636 24936 24642 24948
rect 24636 24908 25636 24936
rect 24636 24896 24642 24908
rect 25608 24880 25636 24908
rect 27522 24896 27528 24948
rect 27580 24896 27586 24948
rect 27709 24939 27767 24945
rect 27709 24905 27721 24939
rect 27755 24905 27767 24939
rect 27709 24899 27767 24905
rect 23201 24871 23259 24877
rect 23201 24837 23213 24871
rect 23247 24837 23259 24871
rect 23937 24871 23995 24877
rect 23937 24868 23949 24871
rect 23201 24831 23259 24837
rect 23308 24840 23949 24868
rect 22235 24772 22508 24800
rect 22235 24769 22247 24772
rect 22189 24763 22247 24769
rect 20180 24704 20392 24732
rect 20548 24704 21128 24732
rect 19536 24636 20208 24664
rect 18138 24596 18144 24608
rect 17880 24568 18144 24596
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 18874 24556 18880 24608
rect 18932 24596 18938 24608
rect 19536 24596 19564 24636
rect 20180 24608 20208 24636
rect 20254 24624 20260 24676
rect 20312 24624 20318 24676
rect 18932 24568 19564 24596
rect 18932 24556 18938 24568
rect 19886 24556 19892 24608
rect 19944 24556 19950 24608
rect 20162 24556 20168 24608
rect 20220 24556 20226 24608
rect 20364 24596 20392 24704
rect 21358 24692 21364 24744
rect 21416 24732 21422 24744
rect 21928 24732 21956 24760
rect 21416 24704 21956 24732
rect 21416 24692 21422 24704
rect 20438 24624 20444 24676
rect 20496 24624 20502 24676
rect 20533 24667 20591 24673
rect 20533 24633 20545 24667
rect 20579 24664 20591 24667
rect 20622 24664 20628 24676
rect 20579 24636 20628 24664
rect 20579 24633 20591 24636
rect 20533 24627 20591 24633
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 20898 24624 20904 24676
rect 20956 24664 20962 24676
rect 22204 24664 22232 24763
rect 22830 24760 22836 24812
rect 22888 24800 22894 24812
rect 23017 24803 23075 24809
rect 23017 24800 23029 24803
rect 22888 24772 23029 24800
rect 22888 24760 22894 24772
rect 23017 24769 23029 24772
rect 23063 24769 23075 24803
rect 23216 24800 23244 24831
rect 23308 24809 23336 24840
rect 23937 24837 23949 24840
rect 23983 24837 23995 24871
rect 23937 24831 23995 24837
rect 24029 24871 24087 24877
rect 24029 24837 24041 24871
rect 24075 24837 24087 24871
rect 24029 24831 24087 24837
rect 23017 24763 23075 24769
rect 23124 24772 23244 24800
rect 23293 24803 23351 24809
rect 23124 24732 23152 24772
rect 23293 24769 23305 24803
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24800 23443 24803
rect 23566 24800 23572 24812
rect 23431 24772 23572 24800
rect 23431 24769 23443 24772
rect 23385 24763 23443 24769
rect 23566 24760 23572 24772
rect 23624 24760 23630 24812
rect 23750 24760 23756 24812
rect 23808 24800 23814 24812
rect 23845 24803 23903 24809
rect 23845 24800 23857 24803
rect 23808 24772 23857 24800
rect 23808 24760 23814 24772
rect 23845 24769 23857 24772
rect 23891 24769 23903 24803
rect 24044 24800 24072 24831
rect 24118 24828 24124 24880
rect 24176 24877 24182 24880
rect 24176 24871 24205 24877
rect 24193 24868 24205 24871
rect 24193 24840 24532 24868
rect 24193 24837 24205 24840
rect 24176 24831 24205 24837
rect 24176 24828 24182 24831
rect 24394 24800 24400 24812
rect 24044 24772 24400 24800
rect 23845 24763 23903 24769
rect 24394 24760 24400 24772
rect 24452 24760 24458 24812
rect 20956 24636 22232 24664
rect 23032 24704 23152 24732
rect 20956 24624 20962 24636
rect 23032 24608 23060 24704
rect 23198 24692 23204 24744
rect 23256 24732 23262 24744
rect 24305 24735 24363 24741
rect 24305 24732 24317 24735
rect 23256 24704 24317 24732
rect 23256 24692 23262 24704
rect 24305 24701 24317 24704
rect 24351 24701 24363 24735
rect 24305 24695 24363 24701
rect 24412 24664 24440 24760
rect 24504 24732 24532 24840
rect 24670 24828 24676 24880
rect 24728 24828 24734 24880
rect 24765 24871 24823 24877
rect 24765 24837 24777 24871
rect 24811 24868 24823 24871
rect 25038 24868 25044 24880
rect 24811 24840 25044 24868
rect 24811 24837 24823 24840
rect 24765 24831 24823 24837
rect 25038 24828 25044 24840
rect 25096 24868 25102 24880
rect 25314 24868 25320 24880
rect 25096 24840 25320 24868
rect 25096 24828 25102 24840
rect 25314 24828 25320 24840
rect 25372 24828 25378 24880
rect 25590 24828 25596 24880
rect 25648 24828 25654 24880
rect 27154 24828 27160 24880
rect 27212 24868 27218 24880
rect 27540 24868 27568 24896
rect 27724 24868 27752 24899
rect 28258 24896 28264 24948
rect 28316 24936 28322 24948
rect 28810 24936 28816 24948
rect 28316 24908 28816 24936
rect 28316 24896 28322 24908
rect 28810 24896 28816 24908
rect 28868 24896 28874 24948
rect 30098 24896 30104 24948
rect 30156 24936 30162 24948
rect 30469 24939 30527 24945
rect 30469 24936 30481 24939
rect 30156 24908 30481 24936
rect 30156 24896 30162 24908
rect 30469 24905 30481 24908
rect 30515 24905 30527 24939
rect 30469 24899 30527 24905
rect 32674 24896 32680 24948
rect 32732 24936 32738 24948
rect 32769 24939 32827 24945
rect 32769 24936 32781 24939
rect 32732 24908 32781 24936
rect 32732 24896 32738 24908
rect 32769 24905 32781 24908
rect 32815 24905 32827 24939
rect 33870 24936 33876 24948
rect 32769 24899 32827 24905
rect 33520 24908 33876 24936
rect 28718 24868 28724 24880
rect 27212 24840 27660 24868
rect 27724 24840 28724 24868
rect 27212 24828 27218 24840
rect 24578 24760 24584 24812
rect 24636 24760 24642 24812
rect 24883 24803 24941 24809
rect 24883 24800 24895 24803
rect 24826 24772 24895 24800
rect 24826 24732 24854 24772
rect 24883 24769 24895 24772
rect 24929 24800 24941 24803
rect 25498 24800 25504 24812
rect 24929 24772 25504 24800
rect 24929 24769 24941 24772
rect 24883 24763 24941 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 26326 24760 26332 24812
rect 26384 24800 26390 24812
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26384 24772 26985 24800
rect 26384 24760 26390 24772
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27065 24803 27123 24809
rect 27065 24769 27077 24803
rect 27111 24800 27123 24803
rect 27338 24800 27344 24812
rect 27111 24772 27344 24800
rect 27111 24769 27123 24772
rect 27065 24763 27123 24769
rect 27338 24760 27344 24772
rect 27396 24760 27402 24812
rect 27433 24803 27491 24809
rect 27433 24769 27445 24803
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 24504 24704 24854 24732
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24701 25099 24735
rect 25041 24695 25099 24701
rect 24486 24664 24492 24676
rect 24412 24636 24492 24664
rect 24486 24624 24492 24636
rect 24544 24624 24550 24676
rect 24578 24624 24584 24676
rect 24636 24664 24642 24676
rect 24854 24664 24860 24676
rect 24636 24636 24860 24664
rect 24636 24624 24642 24636
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 25056 24664 25084 24695
rect 25130 24692 25136 24744
rect 25188 24732 25194 24744
rect 27249 24735 27307 24741
rect 27249 24732 27261 24735
rect 25188 24704 27261 24732
rect 25188 24692 25194 24704
rect 27249 24701 27261 24704
rect 27295 24701 27307 24735
rect 27448 24732 27476 24763
rect 27522 24760 27528 24812
rect 27580 24760 27586 24812
rect 27632 24800 27660 24840
rect 28718 24828 28724 24840
rect 28776 24828 28782 24880
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 27632 24772 27997 24800
rect 27985 24769 27997 24772
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 28166 24760 28172 24812
rect 28224 24760 28230 24812
rect 28258 24760 28264 24812
rect 28316 24760 28322 24812
rect 28828 24809 28856 24896
rect 33137 24871 33195 24877
rect 33137 24837 33149 24871
rect 33183 24868 33195 24871
rect 33520 24868 33548 24908
rect 33870 24896 33876 24908
rect 33928 24936 33934 24948
rect 34057 24939 34115 24945
rect 34057 24936 34069 24939
rect 33928 24908 34069 24936
rect 33928 24896 33934 24908
rect 34057 24905 34069 24908
rect 34103 24905 34115 24939
rect 34057 24899 34115 24905
rect 33183 24840 33548 24868
rect 33183 24837 33195 24840
rect 33137 24831 33195 24837
rect 28353 24803 28411 24809
rect 28353 24769 28365 24803
rect 28399 24800 28411 24803
rect 28813 24803 28871 24809
rect 28399 24772 28764 24800
rect 28399 24769 28411 24772
rect 28353 24763 28411 24769
rect 27893 24735 27951 24741
rect 27893 24732 27905 24735
rect 27448 24704 27905 24732
rect 27249 24695 27307 24701
rect 27893 24701 27905 24704
rect 27939 24701 27951 24735
rect 27893 24695 27951 24701
rect 28077 24735 28135 24741
rect 28077 24701 28089 24735
rect 28123 24732 28135 24735
rect 28276 24732 28304 24760
rect 28123 24704 28304 24732
rect 28123 24701 28135 24704
rect 28077 24695 28135 24701
rect 25056 24636 25360 24664
rect 25332 24608 25360 24636
rect 21082 24596 21088 24608
rect 20364 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24596 21146 24608
rect 22370 24596 22376 24608
rect 21140 24568 22376 24596
rect 21140 24556 21146 24568
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22830 24556 22836 24608
rect 22888 24556 22894 24608
rect 23014 24556 23020 24608
rect 23072 24556 23078 24608
rect 23566 24556 23572 24608
rect 23624 24556 23630 24608
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24596 23719 24599
rect 24302 24596 24308 24608
rect 23707 24568 24308 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 24302 24556 24308 24568
rect 24360 24556 24366 24608
rect 24397 24599 24455 24605
rect 24397 24565 24409 24599
rect 24443 24596 24455 24599
rect 24946 24596 24952 24608
rect 24443 24568 24952 24596
rect 24443 24565 24455 24568
rect 24397 24559 24455 24565
rect 24946 24556 24952 24568
rect 25004 24556 25010 24608
rect 25314 24556 25320 24608
rect 25372 24556 25378 24608
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 26602 24596 26608 24608
rect 25924 24568 26608 24596
rect 25924 24556 25930 24568
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 27157 24599 27215 24605
rect 27157 24565 27169 24599
rect 27203 24596 27215 24599
rect 27798 24596 27804 24608
rect 27203 24568 27804 24596
rect 27203 24565 27215 24568
rect 27157 24559 27215 24565
rect 27798 24556 27804 24568
rect 27856 24556 27862 24608
rect 27908 24596 27936 24695
rect 28442 24692 28448 24744
rect 28500 24692 28506 24744
rect 28736 24732 28764 24772
rect 28813 24769 28825 24803
rect 28859 24769 28871 24803
rect 28813 24763 28871 24769
rect 28902 24760 28908 24812
rect 28960 24760 28966 24812
rect 29356 24803 29414 24809
rect 29356 24769 29368 24803
rect 29402 24800 29414 24803
rect 31205 24803 31263 24809
rect 31205 24800 31217 24803
rect 29402 24772 31217 24800
rect 29402 24769 29414 24772
rect 29356 24763 29414 24769
rect 31205 24769 31217 24772
rect 31251 24769 31263 24803
rect 31205 24763 31263 24769
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24800 31447 24803
rect 32214 24800 32220 24812
rect 31435 24772 32220 24800
rect 31435 24769 31447 24772
rect 31389 24763 31447 24769
rect 32214 24760 32220 24772
rect 32272 24760 32278 24812
rect 32861 24803 32919 24809
rect 32861 24769 32873 24803
rect 32907 24800 32919 24803
rect 32950 24800 32956 24812
rect 32907 24772 32956 24800
rect 32907 24769 32919 24772
rect 32861 24763 32919 24769
rect 32950 24760 32956 24772
rect 33008 24760 33014 24812
rect 33520 24809 33548 24840
rect 33505 24803 33563 24809
rect 33505 24769 33517 24803
rect 33551 24769 33563 24803
rect 33505 24763 33563 24769
rect 33594 24760 33600 24812
rect 33652 24800 33658 24812
rect 34517 24803 34575 24809
rect 34517 24800 34529 24803
rect 33652 24772 34529 24800
rect 33652 24760 33658 24772
rect 34517 24769 34529 24772
rect 34563 24800 34575 24803
rect 36446 24800 36452 24812
rect 34563 24772 36452 24800
rect 34563 24769 34575 24772
rect 34517 24763 34575 24769
rect 36446 24760 36452 24772
rect 36504 24760 36510 24812
rect 28920 24732 28948 24760
rect 28736 24704 28948 24732
rect 29086 24692 29092 24744
rect 29144 24692 29150 24744
rect 30561 24735 30619 24741
rect 30561 24732 30573 24735
rect 30116 24704 30573 24732
rect 28166 24624 28172 24676
rect 28224 24664 28230 24676
rect 28224 24636 28396 24664
rect 28224 24624 28230 24636
rect 28258 24596 28264 24608
rect 27908 24568 28264 24596
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 28368 24605 28396 24636
rect 28626 24624 28632 24676
rect 28684 24664 28690 24676
rect 28905 24667 28963 24673
rect 28905 24664 28917 24667
rect 28684 24636 28917 24664
rect 28684 24624 28690 24636
rect 28905 24633 28917 24636
rect 28951 24633 28963 24667
rect 28905 24627 28963 24633
rect 28994 24624 29000 24676
rect 29052 24624 29058 24676
rect 28353 24599 28411 24605
rect 28353 24565 28365 24599
rect 28399 24565 28411 24599
rect 28353 24559 28411 24565
rect 28718 24556 28724 24608
rect 28776 24556 28782 24608
rect 29012 24596 29040 24624
rect 30116 24596 30144 24704
rect 30561 24701 30573 24704
rect 30607 24701 30619 24735
rect 30561 24695 30619 24701
rect 32125 24735 32183 24741
rect 32125 24701 32137 24735
rect 32171 24732 32183 24735
rect 32398 24732 32404 24744
rect 32171 24704 32404 24732
rect 32171 24701 32183 24704
rect 32125 24695 32183 24701
rect 32398 24692 32404 24704
rect 32456 24692 32462 24744
rect 29012 24568 30144 24596
rect 31938 24556 31944 24608
rect 31996 24556 32002 24608
rect 33778 24556 33784 24608
rect 33836 24556 33842 24608
rect 1104 24506 43884 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 43884 24506
rect 1104 24432 43884 24454
rect 2869 24395 2927 24401
rect 2869 24361 2881 24395
rect 2915 24392 2927 24395
rect 3050 24392 3056 24404
rect 2915 24364 3056 24392
rect 2915 24361 2927 24364
rect 2869 24355 2927 24361
rect 3050 24352 3056 24364
rect 3108 24352 3114 24404
rect 3602 24352 3608 24404
rect 3660 24352 3666 24404
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 3936 24364 4660 24392
rect 3936 24352 3942 24364
rect 3620 24324 3648 24352
rect 4433 24327 4491 24333
rect 4433 24324 4445 24327
rect 3620 24296 4445 24324
rect 4433 24293 4445 24296
rect 4479 24293 4491 24327
rect 4433 24287 4491 24293
rect 4522 24284 4528 24336
rect 4580 24284 4586 24336
rect 4632 24324 4660 24364
rect 4982 24352 4988 24404
rect 5040 24392 5046 24404
rect 6914 24392 6920 24404
rect 5040 24364 5580 24392
rect 5040 24352 5046 24364
rect 5077 24327 5135 24333
rect 5077 24324 5089 24327
rect 4632 24296 5089 24324
rect 5077 24293 5089 24296
rect 5123 24293 5135 24327
rect 5077 24287 5135 24293
rect 1210 24216 1216 24268
rect 1268 24256 1274 24268
rect 1857 24259 1915 24265
rect 1857 24256 1869 24259
rect 1268 24228 1869 24256
rect 1268 24216 1274 24228
rect 1857 24225 1869 24228
rect 1903 24225 1915 24259
rect 1857 24219 1915 24225
rect 2774 24216 2780 24268
rect 2832 24256 2838 24268
rect 3510 24256 3516 24268
rect 2832 24228 3516 24256
rect 2832 24216 2838 24228
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 1578 24148 1584 24200
rect 1636 24148 1642 24200
rect 3329 24191 3387 24197
rect 3329 24188 3341 24191
rect 3068 24160 3341 24188
rect 3068 24132 3096 24160
rect 3329 24157 3341 24160
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24188 3847 24191
rect 3878 24188 3884 24200
rect 3835 24160 3884 24188
rect 3835 24157 3847 24160
rect 3789 24151 3847 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 4062 24148 4068 24200
rect 4120 24148 4126 24200
rect 4540 24197 4568 24284
rect 4706 24216 4712 24268
rect 4764 24216 4770 24268
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24157 4583 24191
rect 4724 24188 4752 24216
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4724 24160 4813 24188
rect 4525 24151 4583 24157
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 4982 24188 4988 24200
rect 4939 24160 4988 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 5074 24148 5080 24200
rect 5132 24188 5138 24200
rect 5169 24191 5227 24197
rect 5169 24188 5181 24191
rect 5132 24160 5181 24188
rect 5132 24148 5138 24160
rect 5169 24157 5181 24160
rect 5215 24157 5227 24191
rect 5169 24151 5227 24157
rect 5258 24148 5264 24200
rect 5316 24188 5322 24200
rect 5552 24197 5580 24364
rect 6426 24364 6920 24392
rect 6426 24256 6454 24364
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 7006 24352 7012 24404
rect 7064 24392 7070 24404
rect 8757 24395 8815 24401
rect 8757 24392 8769 24395
rect 7064 24364 8769 24392
rect 7064 24352 7070 24364
rect 8757 24361 8769 24364
rect 8803 24361 8815 24395
rect 8757 24355 8815 24361
rect 9122 24352 9128 24404
rect 9180 24392 9186 24404
rect 9585 24395 9643 24401
rect 9585 24392 9597 24395
rect 9180 24364 9597 24392
rect 9180 24352 9186 24364
rect 9585 24361 9597 24364
rect 9631 24361 9643 24395
rect 11241 24395 11299 24401
rect 9585 24355 9643 24361
rect 9692 24364 11211 24392
rect 6822 24324 6828 24336
rect 6012 24228 6454 24256
rect 6496 24296 6828 24324
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5316 24160 5457 24188
rect 5316 24148 5322 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 5445 24151 5503 24157
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24188 5595 24191
rect 5583 24160 5856 24188
rect 5583 24157 5595 24160
rect 5537 24151 5595 24157
rect 3050 24080 3056 24132
rect 3108 24080 3114 24132
rect 3237 24123 3295 24129
rect 3237 24089 3249 24123
rect 3283 24120 3295 24123
rect 4080 24120 4108 24148
rect 4709 24123 4767 24129
rect 4709 24120 4721 24123
rect 3283 24092 4108 24120
rect 4540 24092 4721 24120
rect 3283 24089 3295 24092
rect 3237 24083 3295 24089
rect 4062 24012 4068 24064
rect 4120 24052 4126 24064
rect 4540 24052 4568 24092
rect 4709 24089 4721 24092
rect 4755 24089 4767 24123
rect 4709 24083 4767 24089
rect 5350 24080 5356 24132
rect 5408 24080 5414 24132
rect 4120 24024 4568 24052
rect 4120 24012 4126 24024
rect 5626 24012 5632 24064
rect 5684 24052 5690 24064
rect 5721 24055 5779 24061
rect 5721 24052 5733 24055
rect 5684 24024 5733 24052
rect 5684 24012 5690 24024
rect 5721 24021 5733 24024
rect 5767 24021 5779 24055
rect 5828 24052 5856 24160
rect 5902 24148 5908 24200
rect 5960 24148 5966 24200
rect 6012 24197 6040 24228
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 6086 24148 6092 24200
rect 6144 24188 6150 24200
rect 6144 24160 6189 24188
rect 6144 24148 6150 24160
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 6496 24197 6524 24296
rect 6822 24284 6828 24296
rect 6880 24324 6886 24336
rect 7926 24324 7932 24336
rect 6880 24296 7932 24324
rect 6880 24284 6886 24296
rect 7926 24284 7932 24296
rect 7984 24284 7990 24336
rect 8662 24284 8668 24336
rect 8720 24324 8726 24336
rect 9692 24324 9720 24364
rect 8720 24296 9720 24324
rect 9953 24327 10011 24333
rect 8720 24284 8726 24296
rect 7530 24228 8386 24256
rect 6481 24191 6539 24197
rect 6481 24157 6493 24191
rect 6527 24157 6539 24191
rect 6481 24151 6539 24157
rect 6638 24148 6644 24200
rect 6696 24188 6702 24200
rect 7006 24188 7012 24200
rect 6696 24160 7012 24188
rect 6696 24148 6702 24160
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 7530 24197 7558 24228
rect 7157 24191 7215 24197
rect 7157 24157 7169 24191
rect 7203 24157 7215 24191
rect 7157 24151 7215 24157
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7515 24191 7573 24197
rect 7515 24157 7527 24191
rect 7561 24157 7573 24191
rect 7515 24151 7573 24157
rect 5920 24120 5948 24148
rect 6273 24123 6331 24129
rect 6273 24120 6285 24123
rect 5920 24092 6285 24120
rect 6273 24089 6285 24092
rect 6319 24089 6331 24123
rect 6822 24120 6828 24132
rect 6273 24083 6331 24089
rect 6380 24092 6828 24120
rect 6380 24052 6408 24092
rect 6822 24080 6828 24092
rect 6880 24080 6886 24132
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7172 24120 7200 24151
rect 6972 24092 7200 24120
rect 6972 24080 6978 24092
rect 5828 24024 6408 24052
rect 6641 24055 6699 24061
rect 5721 24015 5779 24021
rect 6641 24021 6653 24055
rect 6687 24052 6699 24055
rect 7098 24052 7104 24064
rect 6687 24024 7104 24052
rect 6687 24021 6699 24024
rect 6641 24015 6699 24021
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 7300 24052 7328 24151
rect 7926 24148 7932 24200
rect 7984 24148 7990 24200
rect 8110 24148 8116 24200
rect 8168 24148 8174 24200
rect 8202 24148 8208 24200
rect 8260 24188 8266 24200
rect 8358 24188 8386 24228
rect 8619 24191 8677 24197
rect 8619 24188 8631 24191
rect 8260 24160 8305 24188
rect 8358 24160 8631 24188
rect 8260 24148 8266 24160
rect 8619 24157 8631 24160
rect 8665 24188 8677 24191
rect 8665 24160 8896 24188
rect 8665 24157 8677 24160
rect 8619 24151 8677 24157
rect 7374 24080 7380 24132
rect 7432 24080 7438 24132
rect 8386 24120 8392 24132
rect 7484 24092 8392 24120
rect 7484 24052 7512 24092
rect 8386 24080 8392 24092
rect 8444 24080 8450 24132
rect 8478 24080 8484 24132
rect 8536 24120 8542 24132
rect 8754 24120 8760 24132
rect 8536 24092 8760 24120
rect 8536 24080 8542 24092
rect 8754 24080 8760 24092
rect 8812 24080 8818 24132
rect 7300 24024 7512 24052
rect 7558 24012 7564 24064
rect 7616 24052 7622 24064
rect 7653 24055 7711 24061
rect 7653 24052 7665 24055
rect 7616 24024 7665 24052
rect 7616 24012 7622 24024
rect 7653 24021 7665 24024
rect 7699 24021 7711 24055
rect 8868 24052 8896 24160
rect 8938 24148 8944 24200
rect 8996 24148 9002 24200
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9232 24197 9260 24296
rect 9953 24293 9965 24327
rect 9999 24324 10011 24327
rect 10226 24324 10232 24336
rect 9999 24296 10232 24324
rect 9999 24293 10011 24296
rect 9953 24287 10011 24293
rect 10226 24284 10232 24296
rect 10284 24284 10290 24336
rect 10502 24284 10508 24336
rect 10560 24284 10566 24336
rect 9306 24216 9312 24268
rect 9364 24256 9370 24268
rect 11183 24256 11211 24364
rect 11241 24361 11253 24395
rect 11287 24392 11299 24395
rect 11330 24392 11336 24404
rect 11287 24364 11336 24392
rect 11287 24361 11299 24364
rect 11241 24355 11299 24361
rect 11330 24352 11336 24364
rect 11388 24352 11394 24404
rect 11606 24352 11612 24404
rect 11664 24392 11670 24404
rect 11885 24395 11943 24401
rect 11885 24392 11897 24395
rect 11664 24364 11897 24392
rect 11664 24352 11670 24364
rect 11885 24361 11897 24364
rect 11931 24361 11943 24395
rect 11885 24355 11943 24361
rect 11974 24352 11980 24404
rect 12032 24392 12038 24404
rect 13722 24392 13728 24404
rect 12032 24364 13728 24392
rect 12032 24352 12038 24364
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 14461 24395 14519 24401
rect 14461 24392 14473 24395
rect 14148 24364 14473 24392
rect 14148 24352 14154 24364
rect 14461 24361 14473 24364
rect 14507 24361 14519 24395
rect 14461 24355 14519 24361
rect 15289 24395 15347 24401
rect 15289 24361 15301 24395
rect 15335 24392 15347 24395
rect 15470 24392 15476 24404
rect 15335 24364 15476 24392
rect 15335 24361 15347 24364
rect 15289 24355 15347 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 15749 24395 15807 24401
rect 15749 24361 15761 24395
rect 15795 24392 15807 24395
rect 16574 24392 16580 24404
rect 15795 24364 16580 24392
rect 15795 24361 15807 24364
rect 15749 24355 15807 24361
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 17865 24395 17923 24401
rect 17865 24361 17877 24395
rect 17911 24392 17923 24395
rect 17954 24392 17960 24404
rect 17911 24364 17960 24392
rect 17911 24361 17923 24364
rect 17865 24355 17923 24361
rect 17954 24352 17960 24364
rect 18012 24392 18018 24404
rect 18782 24392 18788 24404
rect 18012 24364 18788 24392
rect 18012 24352 18018 24364
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 19886 24392 19892 24404
rect 18892 24364 19892 24392
rect 11882 24256 11888 24268
rect 9364 24228 11100 24256
rect 11183 24228 11888 24256
rect 9364 24216 9370 24228
rect 9462 24197 9490 24228
rect 11072 24200 11100 24228
rect 9217 24191 9275 24197
rect 9088 24160 9133 24188
rect 9088 24148 9094 24160
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9447 24191 9505 24197
rect 9447 24157 9459 24191
rect 9493 24157 9505 24191
rect 9447 24151 9505 24157
rect 9674 24148 9680 24200
rect 9732 24148 9738 24200
rect 10686 24148 10692 24200
rect 10744 24148 10750 24200
rect 10962 24148 10968 24200
rect 11020 24148 11026 24200
rect 11054 24148 11060 24200
rect 11112 24148 11118 24200
rect 11238 24148 11244 24200
rect 11296 24188 11302 24200
rect 11333 24191 11391 24197
rect 11333 24188 11345 24191
rect 11296 24160 11345 24188
rect 11296 24148 11302 24160
rect 11333 24157 11345 24160
rect 11379 24157 11391 24191
rect 11440 24188 11468 24228
rect 11882 24216 11888 24228
rect 11940 24216 11946 24268
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 11440 24160 11529 24188
rect 11333 24151 11391 24157
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11606 24148 11612 24200
rect 11664 24148 11670 24200
rect 11701 24191 11759 24197
rect 11701 24157 11713 24191
rect 11747 24188 11759 24191
rect 11992 24188 12020 24352
rect 13354 24324 13360 24336
rect 13004 24296 13360 24324
rect 12710 24216 12716 24268
rect 12768 24216 12774 24268
rect 11747 24160 12020 24188
rect 11747 24157 11759 24160
rect 11701 24151 11759 24157
rect 12894 24148 12900 24200
rect 12952 24148 12958 24200
rect 13004 24197 13032 24296
rect 13354 24284 13360 24296
rect 13412 24284 13418 24336
rect 13909 24327 13967 24333
rect 13909 24324 13921 24327
rect 13464 24296 13921 24324
rect 13464 24256 13492 24296
rect 13909 24293 13921 24296
rect 13955 24293 13967 24327
rect 14366 24324 14372 24336
rect 13909 24287 13967 24293
rect 14016 24296 14372 24324
rect 13814 24256 13820 24268
rect 13280 24228 13492 24256
rect 13648 24228 13820 24256
rect 13280 24197 13308 24228
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24157 13047 24191
rect 12989 24151 13047 24157
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24157 13323 24191
rect 13265 24151 13323 24157
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24188 13415 24191
rect 13648 24188 13676 24228
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 13403 24160 13676 24188
rect 13403 24157 13415 24160
rect 13357 24151 13415 24157
rect 9306 24080 9312 24132
rect 9364 24080 9370 24132
rect 9692 24120 9720 24148
rect 10873 24123 10931 24129
rect 10873 24120 10885 24123
rect 9692 24092 10885 24120
rect 10873 24089 10885 24092
rect 10919 24120 10931 24123
rect 10919 24092 11054 24120
rect 10919 24089 10931 24092
rect 10873 24083 10931 24089
rect 9490 24052 9496 24064
rect 8868 24024 9496 24052
rect 7653 24015 7711 24021
rect 9490 24012 9496 24024
rect 9548 24012 9554 24064
rect 11026 24052 11054 24092
rect 12066 24080 12072 24132
rect 12124 24120 12130 24132
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 12124 24092 12265 24120
rect 12124 24080 12130 24092
rect 12253 24089 12265 24092
rect 12299 24089 12311 24123
rect 13188 24120 13216 24151
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 13906 24188 13912 24200
rect 13780 24160 13912 24188
rect 13780 24148 13786 24160
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 13446 24120 13452 24132
rect 13188 24092 13452 24120
rect 12253 24083 12311 24089
rect 13446 24080 13452 24092
rect 13504 24080 13510 24132
rect 13541 24123 13599 24129
rect 13541 24089 13553 24123
rect 13587 24089 13599 24123
rect 13541 24083 13599 24089
rect 13633 24123 13691 24129
rect 13633 24089 13645 24123
rect 13679 24120 13691 24123
rect 14016 24120 14044 24296
rect 14366 24284 14372 24296
rect 14424 24284 14430 24336
rect 14476 24296 15056 24324
rect 14090 24216 14096 24268
rect 14148 24256 14154 24268
rect 14476 24256 14504 24296
rect 14148 24228 14504 24256
rect 15028 24256 15056 24296
rect 15378 24284 15384 24336
rect 15436 24324 15442 24336
rect 15562 24324 15568 24336
rect 15436 24296 15568 24324
rect 15436 24284 15442 24296
rect 15562 24284 15568 24296
rect 15620 24324 15626 24336
rect 16666 24324 16672 24336
rect 15620 24296 16672 24324
rect 15620 24284 15626 24296
rect 16666 24284 16672 24296
rect 16724 24324 16730 24336
rect 17218 24324 17224 24336
rect 16724 24296 17224 24324
rect 16724 24284 16730 24296
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 17310 24284 17316 24336
rect 17368 24324 17374 24336
rect 17368 24296 18184 24324
rect 17368 24284 17374 24296
rect 18046 24256 18052 24268
rect 15028 24228 18052 24256
rect 14148 24216 14154 24228
rect 18046 24216 18052 24228
rect 18104 24216 18110 24268
rect 18156 24256 18184 24296
rect 18506 24284 18512 24336
rect 18564 24324 18570 24336
rect 18892 24324 18920 24364
rect 19886 24352 19892 24364
rect 19944 24392 19950 24404
rect 21361 24395 21419 24401
rect 21361 24392 21373 24395
rect 19944 24364 21373 24392
rect 19944 24352 19950 24364
rect 21361 24361 21373 24364
rect 21407 24361 21419 24395
rect 21361 24355 21419 24361
rect 21545 24395 21603 24401
rect 21545 24361 21557 24395
rect 21591 24392 21603 24395
rect 21634 24392 21640 24404
rect 21591 24364 21640 24392
rect 21591 24361 21603 24364
rect 21545 24355 21603 24361
rect 18564 24296 18920 24324
rect 18564 24284 18570 24296
rect 18966 24284 18972 24336
rect 19024 24324 19030 24336
rect 20070 24324 20076 24336
rect 19024 24296 20076 24324
rect 19024 24284 19030 24296
rect 20070 24284 20076 24296
rect 20128 24284 20134 24336
rect 20162 24284 20168 24336
rect 20220 24324 20226 24336
rect 21376 24324 21404 24355
rect 21634 24352 21640 24364
rect 21692 24352 21698 24404
rect 21726 24352 21732 24404
rect 21784 24352 21790 24404
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24361 22155 24395
rect 23198 24392 23204 24404
rect 22097 24355 22155 24361
rect 22296 24364 23204 24392
rect 21744 24324 21772 24352
rect 20220 24296 20944 24324
rect 21376 24296 21772 24324
rect 20220 24284 20226 24296
rect 20254 24256 20260 24268
rect 18156 24228 20260 24256
rect 20254 24216 20260 24228
rect 20312 24216 20318 24268
rect 20916 24265 20944 24296
rect 20901 24259 20959 24265
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 22112 24256 22140 24355
rect 20947 24228 22140 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 14645 24191 14703 24197
rect 14645 24188 14657 24191
rect 13679 24092 14044 24120
rect 14476 24160 14657 24188
rect 13679 24089 13691 24092
rect 13633 24083 13691 24089
rect 13556 24052 13584 24083
rect 14182 24052 14188 24064
rect 11026 24024 14188 24052
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 14476 24052 14504 24160
rect 14645 24157 14657 24160
rect 14691 24157 14703 24191
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14645 24151 14703 24157
rect 14752 24160 14933 24188
rect 14550 24080 14556 24132
rect 14608 24120 14614 24132
rect 14752 24120 14780 24160
rect 14921 24157 14933 24160
rect 14967 24188 14979 24191
rect 15565 24191 15623 24197
rect 15565 24188 15577 24191
rect 14967 24160 15577 24188
rect 14967 24157 14979 24160
rect 14921 24151 14979 24157
rect 15565 24157 15577 24160
rect 15611 24157 15623 24191
rect 15565 24151 15623 24157
rect 14608 24092 14780 24120
rect 14829 24123 14887 24129
rect 14608 24080 14614 24092
rect 14829 24089 14841 24123
rect 14875 24120 14887 24123
rect 15286 24120 15292 24132
rect 14875 24092 15292 24120
rect 14875 24089 14887 24092
rect 14829 24083 14887 24089
rect 15286 24080 15292 24092
rect 15344 24080 15350 24132
rect 15381 24123 15439 24129
rect 15381 24089 15393 24123
rect 15427 24089 15439 24123
rect 15580 24120 15608 24151
rect 15654 24148 15660 24200
rect 15712 24188 15718 24200
rect 16114 24188 16120 24200
rect 15712 24160 16120 24188
rect 15712 24148 15718 24160
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 16482 24148 16488 24200
rect 16540 24148 16546 24200
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16942 24188 16948 24200
rect 16899 24160 16948 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17218 24148 17224 24200
rect 17276 24148 17282 24200
rect 17405 24191 17463 24197
rect 17405 24157 17417 24191
rect 17451 24188 17463 24191
rect 17954 24188 17960 24200
rect 17451 24160 17960 24188
rect 17451 24157 17463 24160
rect 17405 24151 17463 24157
rect 17954 24148 17960 24160
rect 18012 24148 18018 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24157 18291 24191
rect 18233 24151 18291 24157
rect 17310 24120 17316 24132
rect 15580 24092 17316 24120
rect 15381 24083 15439 24089
rect 15396 24052 15424 24083
rect 17310 24080 17316 24092
rect 17368 24080 17374 24132
rect 18248 24120 18276 24151
rect 18598 24148 18604 24200
rect 18656 24148 18662 24200
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 19058 24148 19064 24200
rect 19116 24148 19122 24200
rect 19426 24148 19432 24200
rect 19484 24148 19490 24200
rect 19702 24188 19708 24200
rect 19628 24160 19708 24188
rect 18892 24120 18920 24148
rect 19628 24120 19656 24160
rect 19702 24148 19708 24160
rect 19760 24148 19766 24200
rect 19794 24148 19800 24200
rect 19852 24188 19858 24200
rect 20533 24191 20591 24197
rect 19852 24160 20484 24188
rect 19852 24148 19858 24160
rect 20456 24132 20484 24160
rect 20533 24157 20545 24191
rect 20579 24188 20591 24191
rect 20806 24188 20812 24200
rect 20579 24160 20812 24188
rect 20579 24157 20591 24160
rect 20533 24151 20591 24157
rect 19978 24120 19984 24132
rect 18248 24092 18920 24120
rect 19306 24092 19656 24120
rect 19720 24092 19984 24120
rect 15562 24052 15568 24064
rect 14476 24024 15568 24052
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 15930 24012 15936 24064
rect 15988 24012 15994 24064
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 17770 24052 17776 24064
rect 16356 24024 17776 24052
rect 16356 24012 16362 24024
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 19306 24052 19334 24092
rect 18380 24024 19334 24052
rect 19613 24055 19671 24061
rect 18380 24012 18386 24024
rect 19613 24021 19625 24055
rect 19659 24052 19671 24055
rect 19720 24052 19748 24092
rect 19978 24080 19984 24092
rect 20036 24080 20042 24132
rect 20438 24080 20444 24132
rect 20496 24080 20502 24132
rect 19659 24024 19748 24052
rect 19659 24021 19671 24024
rect 19613 24015 19671 24021
rect 19794 24012 19800 24064
rect 19852 24052 19858 24064
rect 20070 24052 20076 24064
rect 19852 24024 20076 24052
rect 19852 24012 19858 24024
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 20162 24012 20168 24064
rect 20220 24052 20226 24064
rect 20548 24052 20576 24151
rect 20806 24148 20812 24160
rect 20864 24148 20870 24200
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21082 24188 21088 24200
rect 21039 24160 21088 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21082 24148 21088 24160
rect 21140 24148 21146 24200
rect 21174 24148 21180 24200
rect 21232 24188 21238 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21232 24160 21373 24188
rect 21232 24148 21238 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21542 24148 21548 24200
rect 21600 24188 21606 24200
rect 21729 24191 21787 24197
rect 21729 24188 21741 24191
rect 21600 24160 21741 24188
rect 21600 24148 21606 24160
rect 21729 24157 21741 24160
rect 21775 24157 21787 24191
rect 21729 24151 21787 24157
rect 22094 24148 22100 24200
rect 22152 24148 22158 24200
rect 22296 24120 22324 24364
rect 23198 24352 23204 24364
rect 23256 24392 23262 24404
rect 23385 24395 23443 24401
rect 23385 24392 23397 24395
rect 23256 24364 23397 24392
rect 23256 24352 23262 24364
rect 23385 24361 23397 24364
rect 23431 24361 23443 24395
rect 23385 24355 23443 24361
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 24026 24392 24032 24404
rect 23891 24364 24032 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 24762 24352 24768 24404
rect 24820 24352 24826 24404
rect 25038 24352 25044 24404
rect 25096 24352 25102 24404
rect 25406 24352 25412 24404
rect 25464 24392 25470 24404
rect 26326 24392 26332 24404
rect 25464 24364 26332 24392
rect 25464 24352 25470 24364
rect 26326 24352 26332 24364
rect 26384 24352 26390 24404
rect 27154 24352 27160 24404
rect 27212 24352 27218 24404
rect 27522 24352 27528 24404
rect 27580 24352 27586 24404
rect 27706 24352 27712 24404
rect 27764 24392 27770 24404
rect 28994 24392 29000 24404
rect 27764 24364 29000 24392
rect 27764 24352 27770 24364
rect 28994 24352 29000 24364
rect 29052 24392 29058 24404
rect 29733 24395 29791 24401
rect 29733 24392 29745 24395
rect 29052 24364 29745 24392
rect 29052 24352 29058 24364
rect 29733 24361 29745 24364
rect 29779 24392 29791 24395
rect 30190 24392 30196 24404
rect 29779 24364 30196 24392
rect 29779 24361 29791 24364
rect 29733 24355 29791 24361
rect 30190 24352 30196 24364
rect 30248 24392 30254 24404
rect 30285 24395 30343 24401
rect 30285 24392 30297 24395
rect 30248 24364 30297 24392
rect 30248 24352 30254 24364
rect 30285 24361 30297 24364
rect 30331 24392 30343 24395
rect 31938 24392 31944 24404
rect 30331 24364 30512 24392
rect 30331 24361 30343 24364
rect 30285 24355 30343 24361
rect 23750 24284 23756 24336
rect 23808 24324 23814 24336
rect 24780 24324 24808 24352
rect 23808 24296 24808 24324
rect 23808 24284 23814 24296
rect 23290 24216 23296 24268
rect 23348 24216 23354 24268
rect 23474 24216 23480 24268
rect 23532 24216 23538 24268
rect 25056 24256 25084 24352
rect 26694 24324 26700 24336
rect 25516 24296 26096 24324
rect 25516 24268 25544 24296
rect 24688 24228 25084 24256
rect 22370 24148 22376 24200
rect 22428 24148 22434 24200
rect 23308 24188 23336 24216
rect 23661 24191 23719 24197
rect 23661 24188 23673 24191
rect 23308 24160 23673 24188
rect 23661 24157 23673 24160
rect 23707 24188 23719 24191
rect 24026 24188 24032 24200
rect 23707 24160 24032 24188
rect 23707 24157 23719 24160
rect 23661 24151 23719 24157
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 24688 24197 24716 24228
rect 25498 24216 25504 24268
rect 25556 24216 25562 24268
rect 25866 24256 25872 24268
rect 25700 24228 25872 24256
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24157 24731 24191
rect 24673 24151 24731 24157
rect 24762 24148 24768 24200
rect 24820 24148 24826 24200
rect 24854 24148 24860 24200
rect 24912 24148 24918 24200
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24188 25099 24191
rect 25590 24188 25596 24200
rect 25087 24160 25596 24188
rect 25087 24157 25099 24160
rect 25041 24151 25099 24157
rect 25590 24148 25596 24160
rect 25648 24148 25654 24200
rect 25700 24197 25728 24228
rect 25866 24216 25872 24228
rect 25924 24216 25930 24268
rect 26068 24197 26096 24296
rect 26528 24296 26700 24324
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24157 25743 24191
rect 25961 24191 26019 24197
rect 25961 24188 25973 24191
rect 25685 24151 25743 24157
rect 25792 24160 25973 24188
rect 20916 24092 22324 24120
rect 20916 24064 20944 24092
rect 23382 24080 23388 24132
rect 23440 24080 23446 24132
rect 24302 24080 24308 24132
rect 24360 24120 24366 24132
rect 24360 24092 24533 24120
rect 24360 24080 24366 24092
rect 20220 24024 20576 24052
rect 20220 24012 20226 24024
rect 20898 24012 20904 24064
rect 20956 24012 20962 24064
rect 20990 24012 20996 24064
rect 21048 24052 21054 24064
rect 21450 24052 21456 24064
rect 21048 24024 21456 24052
rect 21048 24012 21054 24024
rect 21450 24012 21456 24024
rect 21508 24052 21514 24064
rect 21913 24055 21971 24061
rect 21913 24052 21925 24055
rect 21508 24024 21925 24052
rect 21508 24012 21514 24024
rect 21913 24021 21925 24024
rect 21959 24021 21971 24055
rect 21913 24015 21971 24021
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 24118 24052 24124 24064
rect 23532 24024 24124 24052
rect 23532 24012 23538 24024
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24394 24012 24400 24064
rect 24452 24012 24458 24064
rect 24505 24052 24533 24092
rect 24578 24080 24584 24132
rect 24636 24120 24642 24132
rect 25792 24120 25820 24160
rect 25961 24157 25973 24160
rect 26007 24157 26019 24191
rect 25961 24151 26019 24157
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 24636 24092 25820 24120
rect 24636 24080 24642 24092
rect 25866 24080 25872 24132
rect 25924 24080 25930 24132
rect 26068 24120 26096 24151
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26528 24197 26556 24296
rect 26694 24284 26700 24296
rect 26752 24324 26758 24336
rect 27172 24324 27200 24352
rect 26752 24296 27200 24324
rect 26752 24284 26758 24296
rect 26878 24256 26884 24268
rect 26620 24228 26884 24256
rect 26620 24197 26648 24228
rect 26878 24216 26884 24228
rect 26936 24216 26942 24268
rect 26329 24191 26387 24197
rect 26329 24188 26341 24191
rect 26200 24160 26341 24188
rect 26200 24148 26206 24160
rect 26329 24157 26341 24160
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 26513 24191 26571 24197
rect 26513 24157 26525 24191
rect 26559 24157 26571 24191
rect 26513 24151 26571 24157
rect 26605 24191 26663 24197
rect 26605 24157 26617 24191
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 27433 24191 27491 24197
rect 27433 24157 27445 24191
rect 27479 24157 27491 24191
rect 27540 24188 27568 24352
rect 27798 24284 27804 24336
rect 27856 24324 27862 24336
rect 28718 24324 28724 24336
rect 27856 24296 28724 24324
rect 27856 24284 27862 24296
rect 28718 24284 28724 24296
rect 28776 24284 28782 24336
rect 30484 24265 30512 24364
rect 30668 24364 31944 24392
rect 30469 24259 30527 24265
rect 30469 24225 30481 24259
rect 30515 24225 30527 24259
rect 30469 24219 30527 24225
rect 27617 24191 27675 24197
rect 27617 24188 27629 24191
rect 27540 24160 27629 24188
rect 27433 24151 27491 24157
rect 27617 24157 27629 24160
rect 27663 24157 27675 24191
rect 27617 24151 27675 24157
rect 26712 24120 26740 24151
rect 26970 24120 26976 24132
rect 26068 24092 26418 24120
rect 25222 24052 25228 24064
rect 24505 24024 25228 24052
rect 25222 24012 25228 24024
rect 25280 24012 25286 24064
rect 25682 24012 25688 24064
rect 25740 24052 25746 24064
rect 26142 24052 26148 24064
rect 25740 24024 26148 24052
rect 25740 24012 25746 24024
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26280 24061 26286 24064
rect 26237 24055 26286 24061
rect 26237 24021 26249 24055
rect 26283 24021 26286 24055
rect 26237 24015 26286 24021
rect 26280 24012 26286 24015
rect 26338 24012 26344 24064
rect 26390 24052 26418 24092
rect 26712 24092 26976 24120
rect 26712 24052 26740 24092
rect 26970 24080 26976 24092
rect 27028 24080 27034 24132
rect 27448 24120 27476 24151
rect 27798 24148 27804 24200
rect 27856 24148 27862 24200
rect 30668 24197 30696 24364
rect 31938 24352 31944 24364
rect 31996 24352 32002 24404
rect 33778 24352 33784 24404
rect 33836 24352 33842 24404
rect 32122 24216 32128 24268
rect 32180 24256 32186 24268
rect 32401 24259 32459 24265
rect 32401 24256 32413 24259
rect 32180 24228 32413 24256
rect 32180 24216 32186 24228
rect 32401 24225 32413 24228
rect 32447 24225 32459 24259
rect 32401 24219 32459 24225
rect 30653 24191 30711 24197
rect 30653 24157 30665 24191
rect 30699 24157 30711 24191
rect 30653 24151 30711 24157
rect 30929 24191 30987 24197
rect 30929 24157 30941 24191
rect 30975 24157 30987 24191
rect 30929 24151 30987 24157
rect 32668 24191 32726 24197
rect 32668 24157 32680 24191
rect 32714 24188 32726 24191
rect 33796 24188 33824 24352
rect 32714 24160 33824 24188
rect 32714 24157 32726 24160
rect 32668 24151 32726 24157
rect 27522 24120 27528 24132
rect 27448 24092 27528 24120
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 27709 24123 27767 24129
rect 27709 24089 27721 24123
rect 27755 24089 27767 24123
rect 27709 24083 27767 24089
rect 26390 24024 26740 24052
rect 26878 24012 26884 24064
rect 26936 24012 26942 24064
rect 27154 24012 27160 24064
rect 27212 24052 27218 24064
rect 27249 24055 27307 24061
rect 27249 24052 27261 24055
rect 27212 24024 27261 24052
rect 27212 24012 27218 24024
rect 27249 24021 27261 24024
rect 27295 24052 27307 24055
rect 27724 24052 27752 24083
rect 27890 24080 27896 24132
rect 27948 24120 27954 24132
rect 28077 24123 28135 24129
rect 28077 24120 28089 24123
rect 27948 24092 28089 24120
rect 27948 24080 27954 24092
rect 28077 24089 28089 24092
rect 28123 24089 28135 24123
rect 28077 24083 28135 24089
rect 28905 24123 28963 24129
rect 28905 24089 28917 24123
rect 28951 24120 28963 24123
rect 29086 24120 29092 24132
rect 28951 24092 29092 24120
rect 28951 24089 28963 24092
rect 28905 24083 28963 24089
rect 29086 24080 29092 24092
rect 29144 24120 29150 24132
rect 29454 24120 29460 24132
rect 29144 24092 29460 24120
rect 29144 24080 29150 24092
rect 29454 24080 29460 24092
rect 29512 24120 29518 24132
rect 30944 24120 30972 24151
rect 31174 24123 31232 24129
rect 31174 24120 31186 24123
rect 29512 24092 30972 24120
rect 31036 24092 31186 24120
rect 29512 24080 29518 24092
rect 27295 24024 27752 24052
rect 27295 24021 27307 24024
rect 27249 24015 27307 24021
rect 27982 24012 27988 24064
rect 28040 24012 28046 24064
rect 30837 24055 30895 24061
rect 30837 24021 30849 24055
rect 30883 24052 30895 24055
rect 31036 24052 31064 24092
rect 31174 24089 31186 24092
rect 31220 24089 31232 24123
rect 31174 24083 31232 24089
rect 30883 24024 31064 24052
rect 30883 24021 30895 24024
rect 30837 24015 30895 24021
rect 32306 24012 32312 24064
rect 32364 24012 32370 24064
rect 33778 24012 33784 24064
rect 33836 24012 33842 24064
rect 1104 23962 43884 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 43884 23962
rect 1104 23888 43884 23910
rect 1949 23851 2007 23857
rect 1949 23817 1961 23851
rect 1995 23848 2007 23851
rect 4062 23848 4068 23860
rect 1995 23820 4068 23848
rect 1995 23817 2007 23820
rect 1949 23811 2007 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 4764 23820 4844 23848
rect 4764 23808 4770 23820
rect 4816 23789 4844 23820
rect 5534 23808 5540 23860
rect 5592 23808 5598 23860
rect 5718 23808 5724 23860
rect 5776 23848 5782 23860
rect 6733 23851 6791 23857
rect 6733 23848 6745 23851
rect 5776 23820 6745 23848
rect 5776 23808 5782 23820
rect 6733 23817 6745 23820
rect 6779 23817 6791 23851
rect 6733 23811 6791 23817
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 7469 23851 7527 23857
rect 7469 23848 7481 23851
rect 6880 23820 7481 23848
rect 6880 23808 6886 23820
rect 7469 23817 7481 23820
rect 7515 23848 7527 23851
rect 7650 23848 7656 23860
rect 7515 23820 7656 23848
rect 7515 23817 7527 23820
rect 7469 23811 7527 23817
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 8662 23808 8668 23860
rect 8720 23808 8726 23860
rect 8938 23808 8944 23860
rect 8996 23848 9002 23860
rect 9125 23851 9183 23857
rect 9125 23848 9137 23851
rect 8996 23820 9137 23848
rect 8996 23808 9002 23820
rect 9125 23817 9137 23820
rect 9171 23817 9183 23851
rect 9125 23811 9183 23817
rect 9766 23808 9772 23860
rect 9824 23808 9830 23860
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 13078 23848 13084 23860
rect 9916 23820 13084 23848
rect 9916 23808 9922 23820
rect 13078 23808 13084 23820
rect 13136 23808 13142 23860
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 13633 23851 13691 23857
rect 13633 23848 13645 23851
rect 13504 23820 13645 23848
rect 13504 23808 13510 23820
rect 13633 23817 13645 23820
rect 13679 23817 13691 23851
rect 13633 23811 13691 23817
rect 13998 23808 14004 23860
rect 14056 23848 14062 23860
rect 14185 23851 14243 23857
rect 14185 23848 14197 23851
rect 14056 23820 14197 23848
rect 14056 23808 14062 23820
rect 14185 23817 14197 23820
rect 14231 23817 14243 23851
rect 14734 23848 14740 23860
rect 14185 23811 14243 23817
rect 14476 23820 14740 23848
rect 4801 23783 4859 23789
rect 3528 23752 4569 23780
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23712 1639 23715
rect 2130 23712 2136 23724
rect 1627 23684 2136 23712
rect 1627 23681 1639 23684
rect 1581 23675 1639 23681
rect 2130 23672 2136 23684
rect 2188 23672 2194 23724
rect 2308 23715 2366 23721
rect 2308 23681 2320 23715
rect 2354 23712 2366 23715
rect 3142 23712 3148 23724
rect 2354 23684 3148 23712
rect 2354 23681 2366 23684
rect 2308 23675 2366 23681
rect 3142 23672 3148 23684
rect 3200 23672 3206 23724
rect 3326 23672 3332 23724
rect 3384 23712 3390 23724
rect 3528 23721 3556 23752
rect 3513 23715 3571 23721
rect 3513 23712 3525 23715
rect 3384 23684 3525 23712
rect 3384 23672 3390 23684
rect 3513 23681 3525 23684
rect 3559 23681 3571 23715
rect 3513 23675 3571 23681
rect 3786 23672 3792 23724
rect 3844 23712 3850 23724
rect 4541 23721 4569 23752
rect 4801 23749 4813 23783
rect 4847 23749 4859 23783
rect 4801 23743 4859 23749
rect 5184 23752 6408 23780
rect 5184 23724 5212 23752
rect 4433 23715 4491 23721
rect 4433 23712 4445 23715
rect 3844 23684 4445 23712
rect 3844 23672 3850 23684
rect 4433 23681 4445 23684
rect 4479 23681 4491 23715
rect 4433 23675 4491 23681
rect 4526 23715 4584 23721
rect 4526 23681 4538 23715
rect 4572 23681 4584 23715
rect 4526 23675 4584 23681
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23681 4767 23715
rect 4709 23675 4767 23681
rect 4939 23715 4997 23721
rect 4939 23681 4951 23715
rect 4985 23712 4997 23715
rect 5074 23712 5080 23724
rect 4985 23684 5080 23712
rect 4985 23681 4997 23684
rect 4939 23675 4997 23681
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23613 1731 23647
rect 1673 23607 1731 23613
rect 1688 23576 1716 23607
rect 1762 23604 1768 23656
rect 1820 23644 1826 23656
rect 2038 23644 2044 23656
rect 1820 23616 2044 23644
rect 1820 23604 1826 23616
rect 2038 23604 2044 23616
rect 2096 23604 2102 23656
rect 4154 23644 4160 23656
rect 3344 23616 4160 23644
rect 1688 23548 1992 23576
rect 1964 23508 1992 23548
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 3344 23576 3372 23616
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 4724 23644 4752 23675
rect 5074 23672 5080 23684
rect 5132 23672 5138 23724
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23712 5687 23715
rect 5810 23712 5816 23724
rect 5675 23684 5816 23712
rect 5675 23681 5687 23684
rect 5629 23675 5687 23681
rect 4798 23644 4804 23656
rect 4724 23616 4804 23644
rect 4798 23604 4804 23616
rect 4856 23604 4862 23656
rect 5644 23644 5672 23675
rect 5810 23672 5816 23684
rect 5868 23672 5874 23724
rect 5994 23672 6000 23724
rect 6052 23672 6058 23724
rect 6380 23721 6408 23752
rect 7006 23740 7012 23792
rect 7064 23780 7070 23792
rect 8680 23780 8708 23808
rect 9490 23780 9496 23792
rect 7064 23752 8708 23780
rect 8956 23752 9496 23780
rect 7064 23740 7070 23752
rect 6365 23715 6423 23721
rect 6365 23681 6377 23715
rect 6411 23681 6423 23715
rect 6365 23675 6423 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 6730 23712 6736 23724
rect 6595 23684 6736 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 6730 23672 6736 23684
rect 6788 23712 6794 23724
rect 8956 23721 8984 23752
rect 9490 23740 9496 23752
rect 9548 23780 9554 23792
rect 11974 23780 11980 23792
rect 9548 23752 11980 23780
rect 9548 23740 9554 23752
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 13372 23752 14228 23780
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 6788 23684 8953 23712
rect 6788 23672 6794 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 10778 23672 10784 23724
rect 10836 23672 10842 23724
rect 11238 23672 11244 23724
rect 11296 23712 11302 23724
rect 11790 23712 11796 23724
rect 11296 23684 11796 23712
rect 11296 23672 11302 23684
rect 11790 23672 11796 23684
rect 11848 23672 11854 23724
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 12986 23712 12992 23724
rect 12676 23684 12992 23712
rect 12676 23672 12682 23684
rect 12986 23672 12992 23684
rect 13044 23712 13050 23724
rect 13081 23715 13139 23721
rect 13081 23712 13093 23715
rect 13044 23684 13093 23712
rect 13044 23672 13050 23684
rect 13081 23681 13093 23684
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 13262 23672 13268 23724
rect 13320 23672 13326 23724
rect 13372 23721 13400 23752
rect 14200 23724 14228 23752
rect 13357 23715 13415 23721
rect 13357 23681 13369 23715
rect 13403 23681 13415 23715
rect 13357 23675 13415 23681
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 5148 23616 5672 23644
rect 6012 23644 6040 23672
rect 7282 23644 7288 23656
rect 6012 23616 7288 23644
rect 3292 23548 3372 23576
rect 3421 23579 3479 23585
rect 3292 23536 3298 23548
rect 3421 23545 3433 23579
rect 3467 23576 3479 23579
rect 5148 23576 5176 23616
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 7466 23604 7472 23656
rect 7524 23644 7530 23656
rect 7834 23644 7840 23656
rect 7524 23616 7840 23644
rect 7524 23604 7530 23616
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8757 23647 8815 23653
rect 8757 23613 8769 23647
rect 8803 23644 8815 23647
rect 9030 23644 9036 23656
rect 8803 23616 9036 23644
rect 8803 23613 8815 23616
rect 8757 23607 8815 23613
rect 9030 23604 9036 23616
rect 9088 23644 9094 23656
rect 9214 23644 9220 23656
rect 9088 23616 9220 23644
rect 9088 23604 9094 23616
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 10502 23604 10508 23656
rect 10560 23644 10566 23656
rect 10965 23647 11023 23653
rect 10965 23644 10977 23647
rect 10560 23616 10977 23644
rect 10560 23604 10566 23616
rect 10965 23613 10977 23616
rect 11011 23613 11023 23647
rect 11900 23644 11928 23672
rect 13280 23644 13308 23672
rect 11900 23616 13308 23644
rect 10965 23607 11023 23613
rect 3467 23548 5176 23576
rect 3467 23545 3479 23548
rect 3421 23539 3479 23545
rect 5258 23536 5264 23588
rect 5316 23576 5322 23588
rect 8665 23579 8723 23585
rect 8665 23576 8677 23579
rect 5316 23548 8677 23576
rect 5316 23536 5322 23548
rect 8665 23545 8677 23548
rect 8711 23576 8723 23579
rect 9122 23576 9128 23588
rect 8711 23548 9128 23576
rect 8711 23545 8723 23548
rect 8665 23539 8723 23545
rect 9122 23536 9128 23548
rect 9180 23576 9186 23588
rect 9180 23548 10640 23576
rect 9180 23536 9186 23548
rect 10612 23520 10640 23548
rect 10870 23536 10876 23588
rect 10928 23576 10934 23588
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 10928 23548 12173 23576
rect 10928 23536 10934 23548
rect 12161 23545 12173 23548
rect 12207 23545 12219 23579
rect 12161 23539 12219 23545
rect 3326 23508 3332 23520
rect 1964 23480 3332 23508
rect 3326 23468 3332 23480
rect 3384 23468 3390 23520
rect 4062 23468 4068 23520
rect 4120 23508 4126 23520
rect 5077 23511 5135 23517
rect 5077 23508 5089 23511
rect 4120 23480 5089 23508
rect 4120 23468 4126 23480
rect 5077 23477 5089 23480
rect 5123 23477 5135 23511
rect 5077 23471 5135 23477
rect 5166 23468 5172 23520
rect 5224 23508 5230 23520
rect 5626 23508 5632 23520
rect 5224 23480 5632 23508
rect 5224 23468 5230 23480
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 5810 23468 5816 23520
rect 5868 23468 5874 23520
rect 6181 23511 6239 23517
rect 6181 23477 6193 23511
rect 6227 23508 6239 23511
rect 6822 23508 6828 23520
rect 6227 23480 6828 23508
rect 6227 23477 6239 23480
rect 6181 23471 6239 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7006 23468 7012 23520
rect 7064 23468 7070 23520
rect 7834 23468 7840 23520
rect 7892 23468 7898 23520
rect 8202 23468 8208 23520
rect 8260 23468 8266 23520
rect 9950 23468 9956 23520
rect 10008 23508 10014 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 10008 23480 10057 23508
rect 10008 23468 10014 23480
rect 10045 23477 10057 23480
rect 10091 23477 10103 23511
rect 10045 23471 10103 23477
rect 10594 23468 10600 23520
rect 10652 23468 10658 23520
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 11606 23508 11612 23520
rect 10744 23480 11612 23508
rect 10744 23468 10750 23480
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 12176 23508 12204 23539
rect 12250 23536 12256 23588
rect 12308 23576 12314 23588
rect 13464 23576 13492 23675
rect 14182 23672 14188 23724
rect 14240 23672 14246 23724
rect 14476 23721 14504 23820
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 15194 23808 15200 23860
rect 15252 23808 15258 23860
rect 19794 23848 19800 23860
rect 16684 23820 16896 23848
rect 14550 23740 14556 23792
rect 14608 23780 14614 23792
rect 14645 23783 14703 23789
rect 14645 23780 14657 23783
rect 14608 23752 14657 23780
rect 14608 23740 14614 23752
rect 14645 23749 14657 23752
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 14826 23740 14832 23792
rect 14884 23740 14890 23792
rect 16040 23752 16528 23780
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23681 14519 23715
rect 14844 23712 14872 23740
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14844 23684 14933 23712
rect 14461 23675 14519 23681
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 14921 23675 14979 23681
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15930 23672 15936 23724
rect 15988 23672 15994 23724
rect 16040 23721 16068 23752
rect 16025 23715 16083 23721
rect 16025 23681 16037 23715
rect 16071 23681 16083 23715
rect 16025 23675 16083 23681
rect 16393 23715 16451 23721
rect 16393 23681 16405 23715
rect 16439 23681 16451 23715
rect 16393 23675 16451 23681
rect 14274 23604 14280 23656
rect 14332 23644 14338 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 14332 23616 14841 23644
rect 14332 23604 14338 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 14829 23607 14887 23613
rect 15010 23604 15016 23656
rect 15068 23644 15074 23656
rect 15194 23644 15200 23656
rect 15068 23616 15200 23644
rect 15068 23604 15074 23616
rect 15194 23604 15200 23616
rect 15252 23644 15258 23656
rect 15381 23647 15439 23653
rect 15381 23644 15393 23647
rect 15252 23616 15393 23644
rect 15252 23604 15258 23616
rect 15381 23613 15393 23616
rect 15427 23613 15439 23647
rect 15381 23607 15439 23613
rect 16040 23576 16068 23675
rect 12308 23548 16068 23576
rect 16408 23576 16436 23675
rect 16500 23644 16528 23752
rect 16684 23721 16712 23820
rect 16868 23780 16896 23820
rect 18432 23820 19800 23848
rect 17494 23780 17500 23792
rect 16868 23752 17500 23780
rect 17494 23740 17500 23752
rect 17552 23780 17558 23792
rect 17589 23783 17647 23789
rect 17589 23780 17601 23783
rect 17552 23752 17601 23780
rect 17552 23740 17558 23752
rect 17589 23749 17601 23752
rect 17635 23749 17647 23783
rect 17589 23743 17647 23749
rect 17954 23740 17960 23792
rect 18012 23780 18018 23792
rect 18432 23780 18460 23820
rect 19794 23808 19800 23820
rect 19852 23808 19858 23860
rect 20622 23848 20628 23860
rect 19895 23820 20628 23848
rect 18012 23752 18460 23780
rect 18012 23740 18018 23752
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16758 23672 16764 23724
rect 16816 23672 16822 23724
rect 16945 23715 17003 23721
rect 16853 23705 16911 23711
rect 16776 23644 16804 23672
rect 16853 23671 16865 23705
rect 16899 23671 16911 23705
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 17175 23684 17632 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 16853 23665 16911 23671
rect 16500 23616 16804 23644
rect 16868 23576 16896 23665
rect 16960 23644 16988 23675
rect 17604 23656 17632 23684
rect 17770 23672 17776 23724
rect 17828 23712 17834 23724
rect 18432 23721 18460 23752
rect 18506 23740 18512 23792
rect 18564 23740 18570 23792
rect 19895 23780 19923 23820
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 20714 23808 20720 23860
rect 20772 23848 20778 23860
rect 21082 23848 21088 23860
rect 20772 23820 21088 23848
rect 20772 23808 20778 23820
rect 21082 23808 21088 23820
rect 21140 23848 21146 23860
rect 21177 23851 21235 23857
rect 21177 23848 21189 23851
rect 21140 23820 21189 23848
rect 21140 23808 21146 23820
rect 21177 23817 21189 23820
rect 21223 23848 21235 23851
rect 21266 23848 21272 23860
rect 21223 23820 21272 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 21453 23851 21511 23857
rect 21453 23848 21465 23851
rect 21416 23820 21465 23848
rect 21416 23808 21422 23820
rect 21453 23817 21465 23820
rect 21499 23817 21511 23851
rect 21634 23848 21640 23860
rect 21453 23811 21511 23817
rect 21560 23820 21640 23848
rect 19260 23752 19756 23780
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 17828 23684 18061 23712
rect 17828 23672 17834 23684
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23681 18475 23715
rect 18524 23711 18552 23740
rect 19260 23724 19288 23752
rect 18966 23721 18972 23724
rect 18943 23715 18972 23721
rect 18417 23675 18475 23681
rect 18509 23705 18567 23711
rect 18509 23671 18521 23705
rect 18555 23671 18567 23705
rect 18943 23681 18955 23715
rect 18943 23675 18972 23681
rect 18966 23672 18972 23675
rect 19024 23672 19030 23724
rect 19242 23672 19248 23724
rect 19300 23672 19306 23724
rect 19334 23672 19340 23724
rect 19392 23672 19398 23724
rect 19728 23721 19756 23752
rect 19812 23752 19923 23780
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 18509 23665 18567 23671
rect 16960 23616 17264 23644
rect 17126 23576 17132 23588
rect 16408 23548 17132 23576
rect 12308 23536 12314 23548
rect 17126 23536 17132 23548
rect 17184 23536 17190 23588
rect 17236 23576 17264 23616
rect 17586 23604 17592 23656
rect 17644 23604 17650 23656
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 18138 23576 18144 23588
rect 17236 23548 18144 23576
rect 18138 23536 18144 23548
rect 18196 23536 18202 23588
rect 18233 23579 18291 23585
rect 18233 23545 18245 23579
rect 18279 23576 18291 23579
rect 18414 23576 18420 23588
rect 18279 23548 18420 23576
rect 18279 23545 18291 23548
rect 18233 23539 18291 23545
rect 18414 23536 18420 23548
rect 18472 23536 18478 23588
rect 12618 23508 12624 23520
rect 12176 23480 12624 23508
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 12989 23511 13047 23517
rect 12989 23477 13001 23511
rect 13035 23508 13047 23511
rect 13998 23508 14004 23520
rect 13035 23480 14004 23508
rect 13035 23477 13047 23480
rect 12989 23471 13047 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15562 23468 15568 23520
rect 15620 23508 15626 23520
rect 16298 23508 16304 23520
rect 15620 23480 16304 23508
rect 15620 23468 15626 23480
rect 16298 23468 16304 23480
rect 16356 23468 16362 23520
rect 16758 23468 16764 23520
rect 16816 23468 16822 23520
rect 17144 23508 17172 23536
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17144 23480 17233 23508
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 17221 23471 17279 23477
rect 18046 23468 18052 23520
rect 18104 23468 18110 23520
rect 18874 23468 18880 23520
rect 18932 23468 18938 23520
rect 19444 23508 19472 23675
rect 19518 23536 19524 23588
rect 19576 23576 19582 23588
rect 19812 23576 19840 23752
rect 20070 23740 20076 23792
rect 20128 23780 20134 23792
rect 20165 23783 20223 23789
rect 20165 23780 20177 23783
rect 20128 23752 20177 23780
rect 20128 23740 20134 23752
rect 20165 23749 20177 23752
rect 20211 23749 20223 23783
rect 21560 23780 21588 23820
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 23661 23851 23719 23857
rect 22060 23820 23428 23848
rect 22060 23808 22066 23820
rect 23400 23792 23428 23820
rect 23661 23817 23673 23851
rect 23707 23817 23719 23851
rect 23661 23811 23719 23817
rect 22094 23780 22100 23792
rect 20165 23743 20223 23749
rect 20548 23752 21588 23780
rect 21652 23752 22100 23780
rect 20548 23724 20576 23752
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 19576 23548 19840 23576
rect 19904 23684 20269 23712
rect 19904 23576 19932 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20257 23675 20315 23681
rect 20438 23672 20444 23724
rect 20496 23672 20502 23724
rect 20530 23672 20536 23724
rect 20588 23672 20594 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 21376 23721 21404 23752
rect 20901 23715 20959 23721
rect 20901 23712 20913 23715
rect 20772 23684 20913 23712
rect 20772 23672 20778 23684
rect 20901 23681 20913 23684
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 21361 23715 21419 23721
rect 21361 23681 21373 23715
rect 21407 23681 21419 23715
rect 21361 23675 21419 23681
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20990 23644 20996 23656
rect 20036 23616 20996 23644
rect 20036 23604 20042 23616
rect 20990 23604 20996 23616
rect 21048 23644 21054 23656
rect 21100 23644 21128 23675
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 21545 23715 21603 23721
rect 21545 23712 21557 23715
rect 21508 23684 21557 23712
rect 21508 23672 21514 23684
rect 21545 23681 21557 23684
rect 21591 23681 21603 23715
rect 21545 23675 21603 23681
rect 21652 23644 21680 23752
rect 22094 23740 22100 23752
rect 22152 23780 22158 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 22152 23752 22293 23780
rect 22152 23740 22158 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 23014 23780 23020 23792
rect 22281 23743 22339 23749
rect 22388 23752 23020 23780
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 21048 23616 21128 23644
rect 21284 23616 21680 23644
rect 22020 23644 22048 23675
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 22388 23721 22416 23752
rect 23014 23740 23020 23752
rect 23072 23780 23078 23792
rect 23290 23780 23296 23792
rect 23072 23752 23296 23780
rect 23072 23740 23078 23752
rect 23290 23740 23296 23752
rect 23348 23740 23354 23792
rect 23382 23740 23388 23792
rect 23440 23740 23446 23792
rect 23676 23780 23704 23811
rect 23750 23808 23756 23860
rect 23808 23848 23814 23860
rect 25314 23848 25320 23860
rect 23808 23820 25320 23848
rect 23808 23808 23814 23820
rect 24044 23789 24072 23820
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 25498 23808 25504 23860
rect 25556 23808 25562 23860
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 25924 23820 27108 23848
rect 25924 23808 25930 23820
rect 24029 23783 24087 23789
rect 23676 23752 23880 23780
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 22554 23672 22560 23724
rect 22612 23712 22618 23724
rect 23109 23715 23167 23721
rect 23109 23712 23121 23715
rect 22612 23684 23121 23712
rect 22612 23672 22618 23684
rect 23109 23681 23121 23684
rect 23155 23681 23167 23715
rect 23109 23675 23167 23681
rect 23474 23672 23480 23724
rect 23532 23672 23538 23724
rect 23566 23672 23572 23724
rect 23624 23718 23630 23724
rect 23753 23718 23811 23721
rect 23624 23715 23811 23718
rect 23624 23690 23765 23715
rect 23624 23672 23630 23690
rect 23732 23684 23765 23690
rect 23753 23681 23765 23684
rect 23799 23681 23811 23715
rect 23852 23712 23880 23752
rect 24029 23749 24041 23783
rect 24075 23749 24087 23783
rect 24029 23743 24087 23749
rect 24949 23783 25007 23789
rect 24949 23749 24961 23783
rect 24995 23780 25007 23783
rect 25038 23780 25044 23792
rect 24995 23752 25044 23780
rect 24995 23749 25007 23752
rect 24949 23743 25007 23749
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 23852 23684 23889 23712
rect 23753 23675 23811 23681
rect 23492 23644 23520 23672
rect 22020 23616 23520 23644
rect 23861 23644 23889 23684
rect 23934 23672 23940 23724
rect 23992 23672 23998 23724
rect 24118 23672 24124 23724
rect 24176 23712 24182 23724
rect 24762 23712 24768 23724
rect 24176 23684 24768 23712
rect 24176 23672 24182 23684
rect 24762 23672 24768 23684
rect 24820 23672 24826 23724
rect 24854 23672 24860 23724
rect 24912 23712 24918 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24912 23684 25145 23712
rect 24912 23672 24918 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 25409 23715 25467 23721
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 23861 23616 25360 23644
rect 21048 23604 21054 23616
rect 20070 23576 20076 23588
rect 19904 23548 20076 23576
rect 19576 23536 19582 23548
rect 20070 23536 20076 23548
rect 20128 23536 20134 23588
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 20533 23579 20591 23585
rect 20533 23576 20545 23579
rect 20312 23548 20545 23576
rect 20312 23536 20318 23548
rect 20533 23545 20545 23548
rect 20579 23576 20591 23579
rect 21284 23576 21312 23616
rect 20579 23548 21312 23576
rect 20579 23545 20591 23548
rect 20533 23539 20591 23545
rect 21358 23536 21364 23588
rect 21416 23536 21422 23588
rect 21634 23536 21640 23588
rect 21692 23576 21698 23588
rect 22278 23576 22284 23588
rect 21692 23548 22284 23576
rect 21692 23536 21698 23548
rect 22278 23536 22284 23548
rect 22336 23576 22342 23588
rect 22462 23576 22468 23588
rect 22336 23548 22468 23576
rect 22336 23536 22342 23548
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 22557 23579 22615 23585
rect 22557 23545 22569 23579
rect 22603 23576 22615 23579
rect 25038 23576 25044 23588
rect 22603 23548 25044 23576
rect 22603 23545 22615 23548
rect 22557 23539 22615 23545
rect 25038 23536 25044 23548
rect 25096 23576 25102 23588
rect 25225 23579 25283 23585
rect 25225 23576 25237 23579
rect 25096 23548 25237 23576
rect 25096 23536 25102 23548
rect 25225 23545 25237 23548
rect 25271 23545 25283 23579
rect 25225 23539 25283 23545
rect 20346 23508 20352 23520
rect 19444 23480 20352 23508
rect 20346 23468 20352 23480
rect 20404 23508 20410 23520
rect 21266 23508 21272 23520
rect 20404 23480 21272 23508
rect 20404 23468 20410 23480
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 21376 23508 21404 23536
rect 25332 23520 25360 23616
rect 25424 23576 25452 23675
rect 25682 23672 25688 23724
rect 25740 23672 25746 23724
rect 25885 23721 25913 23808
rect 27080 23792 27108 23820
rect 27890 23808 27896 23860
rect 27948 23848 27954 23860
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 27948 23820 28457 23848
rect 27948 23808 27954 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 28445 23811 28503 23817
rect 28905 23851 28963 23857
rect 28905 23817 28917 23851
rect 28951 23848 28963 23851
rect 28994 23848 29000 23860
rect 28951 23820 29000 23848
rect 28951 23817 28963 23820
rect 28905 23811 28963 23817
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 30006 23808 30012 23860
rect 30064 23848 30070 23860
rect 30837 23851 30895 23857
rect 30837 23848 30849 23851
rect 30064 23820 30849 23848
rect 30064 23808 30070 23820
rect 30837 23817 30849 23820
rect 30883 23817 30895 23851
rect 33778 23848 33784 23860
rect 30837 23811 30895 23817
rect 32600 23820 33784 23848
rect 25958 23740 25964 23792
rect 26016 23740 26022 23792
rect 27062 23740 27068 23792
rect 27120 23780 27126 23792
rect 27249 23783 27307 23789
rect 27249 23780 27261 23783
rect 27120 23752 27261 23780
rect 27120 23740 27126 23752
rect 27249 23749 27261 23752
rect 27295 23749 27307 23783
rect 27249 23743 27307 23749
rect 27430 23740 27436 23792
rect 27488 23780 27494 23792
rect 27801 23783 27859 23789
rect 27801 23780 27813 23783
rect 27488 23752 27813 23780
rect 27488 23740 27494 23752
rect 27801 23749 27813 23752
rect 27847 23749 27859 23783
rect 27801 23743 27859 23749
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 26970 23672 26976 23724
rect 27028 23672 27034 23724
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23712 27399 23715
rect 27614 23712 27620 23724
rect 27387 23684 27620 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 27172 23644 27200 23675
rect 27614 23672 27620 23684
rect 27672 23672 27678 23724
rect 27890 23672 27896 23724
rect 27948 23672 27954 23724
rect 29012 23721 29040 23808
rect 29546 23780 29552 23792
rect 29196 23752 29552 23780
rect 29196 23721 29224 23752
rect 29546 23740 29552 23752
rect 29604 23740 29610 23792
rect 31662 23740 31668 23792
rect 31720 23740 31726 23792
rect 27985 23715 28043 23721
rect 27985 23681 27997 23715
rect 28031 23681 28043 23715
rect 27985 23675 28043 23681
rect 28997 23715 29055 23721
rect 28997 23681 29009 23715
rect 29043 23681 29055 23715
rect 28997 23675 29055 23681
rect 29181 23715 29239 23721
rect 29181 23681 29193 23715
rect 29227 23681 29239 23715
rect 29181 23675 29239 23681
rect 29365 23715 29423 23721
rect 29365 23681 29377 23715
rect 29411 23712 29423 23715
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29411 23684 29745 23712
rect 29411 23681 29423 23684
rect 29365 23675 29423 23681
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23712 31631 23715
rect 32306 23712 32312 23724
rect 31619 23684 32312 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 26712 23616 27200 23644
rect 25958 23576 25964 23588
rect 25424 23548 25964 23576
rect 25958 23536 25964 23548
rect 26016 23536 26022 23588
rect 26050 23536 26056 23588
rect 26108 23576 26114 23588
rect 26712 23585 26740 23616
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 28000 23644 28028 23675
rect 32306 23672 32312 23684
rect 32364 23672 32370 23724
rect 32600 23721 32628 23820
rect 33778 23808 33784 23820
rect 33836 23808 33842 23860
rect 32585 23715 32643 23721
rect 32585 23681 32597 23715
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 27856 23616 28028 23644
rect 27856 23604 27862 23616
rect 29454 23604 29460 23656
rect 29512 23604 29518 23656
rect 26697 23579 26755 23585
rect 26697 23576 26709 23579
rect 26108 23548 26709 23576
rect 26108 23536 26114 23548
rect 26697 23545 26709 23548
rect 26743 23545 26755 23579
rect 26697 23539 26755 23545
rect 23750 23508 23756 23520
rect 21376 23480 23756 23508
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 24305 23511 24363 23517
rect 24305 23477 24317 23511
rect 24351 23508 24363 23511
rect 25130 23508 25136 23520
rect 24351 23480 25136 23508
rect 24351 23477 24363 23480
rect 24305 23471 24363 23477
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 25314 23468 25320 23520
rect 25372 23468 25378 23520
rect 25774 23468 25780 23520
rect 25832 23508 25838 23520
rect 26237 23511 26295 23517
rect 26237 23508 26249 23511
rect 25832 23480 26249 23508
rect 25832 23468 25838 23480
rect 26237 23477 26249 23480
rect 26283 23477 26295 23511
rect 26237 23471 26295 23477
rect 27522 23468 27528 23520
rect 27580 23468 27586 23520
rect 28166 23468 28172 23520
rect 28224 23468 28230 23520
rect 33134 23468 33140 23520
rect 33192 23468 33198 23520
rect 1104 23418 43884 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 43884 23418
rect 1104 23344 43884 23366
rect 2866 23264 2872 23316
rect 2924 23264 2930 23316
rect 3326 23264 3332 23316
rect 3384 23304 3390 23316
rect 4893 23307 4951 23313
rect 4893 23304 4905 23307
rect 3384 23276 4905 23304
rect 3384 23264 3390 23276
rect 4893 23273 4905 23276
rect 4939 23273 4951 23307
rect 5629 23307 5687 23313
rect 5629 23304 5641 23307
rect 4893 23267 4951 23273
rect 5184 23276 5641 23304
rect 5184 23236 5212 23276
rect 5629 23273 5641 23276
rect 5675 23273 5687 23307
rect 5629 23267 5687 23273
rect 7098 23264 7104 23316
rect 7156 23264 7162 23316
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 7926 23304 7932 23316
rect 7248 23276 7932 23304
rect 7248 23264 7254 23276
rect 7926 23264 7932 23276
rect 7984 23264 7990 23316
rect 8757 23307 8815 23313
rect 8757 23273 8769 23307
rect 8803 23304 8815 23307
rect 8846 23304 8852 23316
rect 8803 23276 8852 23304
rect 8803 23273 8815 23276
rect 8757 23267 8815 23273
rect 3344 23208 5212 23236
rect 1210 23128 1216 23180
rect 1268 23168 1274 23180
rect 3344 23177 3372 23208
rect 6362 23196 6368 23248
rect 6420 23196 6426 23248
rect 6730 23196 6736 23248
rect 6788 23196 6794 23248
rect 1857 23171 1915 23177
rect 1857 23168 1869 23171
rect 1268 23140 1869 23168
rect 1268 23128 1274 23140
rect 1857 23137 1869 23140
rect 1903 23137 1915 23171
rect 3329 23171 3387 23177
rect 3329 23168 3341 23171
rect 1857 23131 1915 23137
rect 2746 23140 3341 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 2746 23100 2774 23140
rect 3329 23137 3341 23140
rect 3375 23137 3387 23171
rect 3329 23131 3387 23137
rect 3513 23171 3571 23177
rect 3513 23137 3525 23171
rect 3559 23168 3571 23171
rect 3602 23168 3608 23180
rect 3559 23140 3608 23168
rect 3559 23137 3571 23140
rect 3513 23131 3571 23137
rect 3602 23128 3608 23140
rect 3660 23128 3666 23180
rect 4157 23171 4215 23177
rect 4157 23168 4169 23171
rect 3712 23140 4169 23168
rect 1627 23072 2774 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 3234 23060 3240 23112
rect 3292 23060 3298 23112
rect 2130 22992 2136 23044
rect 2188 23032 2194 23044
rect 3712 23032 3740 23140
rect 4157 23137 4169 23140
rect 4203 23137 4215 23171
rect 4614 23168 4620 23180
rect 4157 23131 4215 23137
rect 4412 23140 4620 23168
rect 4062 23060 4068 23112
rect 4120 23100 4126 23112
rect 4412 23109 4440 23140
rect 4614 23128 4620 23140
rect 4672 23168 4678 23180
rect 5902 23168 5908 23180
rect 4672 23140 5111 23168
rect 4672 23128 4678 23140
rect 4249 23103 4307 23109
rect 4249 23100 4261 23103
rect 4120 23072 4261 23100
rect 4120 23060 4126 23072
rect 4249 23069 4261 23072
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 4397 23103 4455 23109
rect 4397 23069 4409 23103
rect 4443 23069 4455 23103
rect 4397 23063 4455 23069
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23069 4583 23103
rect 4525 23063 4583 23069
rect 2188 23004 3740 23032
rect 2188 22992 2194 23004
rect 3252 22976 3280 23004
rect 3786 22992 3792 23044
rect 3844 22992 3850 23044
rect 3973 23035 4031 23041
rect 3973 23001 3985 23035
rect 4019 23001 4031 23035
rect 4540 23032 4568 23063
rect 4706 23060 4712 23112
rect 4764 23109 4770 23112
rect 5083 23109 5111 23140
rect 5276 23140 5672 23168
rect 5276 23109 5304 23140
rect 4764 23100 4772 23109
rect 4985 23103 5043 23109
rect 4764 23072 4809 23100
rect 4764 23063 4772 23072
rect 4985 23069 4997 23103
rect 5031 23100 5043 23103
rect 5078 23103 5136 23109
rect 5031 23069 5044 23100
rect 4985 23063 5044 23069
rect 5078 23069 5090 23103
rect 5124 23069 5136 23103
rect 5078 23063 5136 23069
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5450 23103 5508 23109
rect 5450 23069 5462 23103
rect 5496 23069 5508 23103
rect 5450 23063 5508 23069
rect 4764 23060 4770 23063
rect 3973 22995 4031 23001
rect 4264 23004 4568 23032
rect 1578 22924 1584 22976
rect 1636 22964 1642 22976
rect 3050 22964 3056 22976
rect 1636 22936 3056 22964
rect 1636 22924 1642 22936
rect 3050 22924 3056 22936
rect 3108 22924 3114 22976
rect 3234 22924 3240 22976
rect 3292 22924 3298 22976
rect 3510 22924 3516 22976
rect 3568 22964 3574 22976
rect 3988 22964 4016 22995
rect 4264 22976 4292 23004
rect 4614 22992 4620 23044
rect 4672 22992 4678 23044
rect 3568 22936 4016 22964
rect 3568 22924 3574 22936
rect 4246 22924 4252 22976
rect 4304 22924 4310 22976
rect 5016 22964 5044 23063
rect 5368 22976 5396 23063
rect 5465 23032 5493 23063
rect 5644 23044 5672 23140
rect 5736 23140 5908 23168
rect 5736 23109 5764 23140
rect 5902 23128 5908 23140
rect 5960 23128 5966 23180
rect 6748 23168 6776 23196
rect 6104 23140 6776 23168
rect 7116 23168 7144 23264
rect 8021 23239 8079 23245
rect 8021 23205 8033 23239
rect 8067 23236 8079 23239
rect 8662 23236 8668 23248
rect 8067 23208 8668 23236
rect 8067 23205 8079 23208
rect 8021 23199 8079 23205
rect 8662 23196 8668 23208
rect 8720 23236 8726 23248
rect 8772 23236 8800 23267
rect 8846 23264 8852 23276
rect 8904 23304 8910 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 8904 23276 9137 23304
rect 8904 23264 8910 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10870 23304 10876 23316
rect 9732 23276 10876 23304
rect 9732 23264 9738 23276
rect 10870 23264 10876 23276
rect 10928 23264 10934 23316
rect 11330 23264 11336 23316
rect 11388 23304 11394 23316
rect 11388 23276 12204 23304
rect 11388 23264 11394 23276
rect 8720 23208 8800 23236
rect 8720 23196 8726 23208
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 10744 23208 11560 23236
rect 10744 23196 10750 23208
rect 11422 23168 11428 23180
rect 7116 23140 7236 23168
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23069 5779 23103
rect 5721 23063 5779 23069
rect 5810 23060 5816 23112
rect 5868 23100 5874 23112
rect 6104 23109 6132 23140
rect 6089 23103 6147 23109
rect 5868 23072 5913 23100
rect 5868 23060 5874 23072
rect 6089 23069 6101 23103
rect 6135 23069 6147 23103
rect 6089 23063 6147 23069
rect 6186 23103 6244 23109
rect 6186 23069 6198 23103
rect 6232 23069 6244 23103
rect 6186 23063 6244 23069
rect 5465 23004 5580 23032
rect 5166 22964 5172 22976
rect 5016 22936 5172 22964
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 5350 22924 5356 22976
rect 5408 22924 5414 22976
rect 5552 22964 5580 23004
rect 5626 22992 5632 23044
rect 5684 23032 5690 23044
rect 5997 23035 6055 23041
rect 5997 23032 6009 23035
rect 5684 23004 6009 23032
rect 5684 22992 5690 23004
rect 5997 23001 6009 23004
rect 6043 23001 6055 23035
rect 5997 22995 6055 23001
rect 6197 22964 6225 23063
rect 6730 23060 6736 23112
rect 6788 23100 6794 23112
rect 6917 23103 6975 23109
rect 6917 23100 6929 23103
rect 6788 23072 6929 23100
rect 6788 23060 6794 23072
rect 6917 23069 6929 23072
rect 6963 23069 6975 23103
rect 6917 23063 6975 23069
rect 7010 23103 7068 23109
rect 7010 23069 7022 23103
rect 7056 23100 7068 23103
rect 7098 23100 7104 23112
rect 7056 23072 7104 23100
rect 7056 23069 7068 23072
rect 7010 23063 7068 23069
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 7208 23109 7236 23140
rect 11164 23140 11428 23168
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 7374 23060 7380 23112
rect 7432 23109 7438 23112
rect 7432 23100 7440 23109
rect 9309 23103 9367 23109
rect 7432 23072 7477 23100
rect 7432 23063 7440 23072
rect 9309 23069 9321 23103
rect 9355 23100 9367 23103
rect 10594 23100 10600 23112
rect 9355 23072 10600 23100
rect 9355 23069 9367 23072
rect 9309 23063 9367 23069
rect 7432 23060 7438 23063
rect 10594 23060 10600 23072
rect 10652 23060 10658 23112
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 7285 23035 7343 23041
rect 7285 23032 7297 23035
rect 6932 23004 7297 23032
rect 6932 22976 6960 23004
rect 7285 23001 7297 23004
rect 7331 23001 7343 23035
rect 7285 22995 7343 23001
rect 9576 23035 9634 23041
rect 9576 23001 9588 23035
rect 9622 23032 9634 23035
rect 10318 23032 10324 23044
rect 9622 23004 10324 23032
rect 9622 23001 9634 23004
rect 9576 22995 9634 23001
rect 10318 22992 10324 23004
rect 10376 22992 10382 23044
rect 10796 23032 10824 23063
rect 11054 23060 11060 23112
rect 11112 23100 11118 23112
rect 11164 23100 11192 23140
rect 11422 23128 11428 23140
rect 11480 23128 11486 23180
rect 11532 23177 11560 23208
rect 11882 23196 11888 23248
rect 11940 23196 11946 23248
rect 11517 23171 11575 23177
rect 11517 23137 11529 23171
rect 11563 23137 11575 23171
rect 11900 23168 11928 23196
rect 11900 23140 12021 23168
rect 11517 23131 11575 23137
rect 11112 23072 11192 23100
rect 11112 23060 11118 23072
rect 11238 23060 11244 23112
rect 11296 23060 11302 23112
rect 11606 23060 11612 23112
rect 11664 23060 11670 23112
rect 11993 23109 12021 23140
rect 12176 23109 12204 23276
rect 14826 23264 14832 23316
rect 14884 23304 14890 23316
rect 15654 23304 15660 23316
rect 14884 23276 15660 23304
rect 14884 23264 14890 23276
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16209 23307 16267 23313
rect 16209 23273 16221 23307
rect 16255 23304 16267 23307
rect 17034 23304 17040 23316
rect 16255 23276 17040 23304
rect 16255 23273 16267 23276
rect 16209 23267 16267 23273
rect 17034 23264 17040 23276
rect 17092 23264 17098 23316
rect 17129 23307 17187 23313
rect 17129 23273 17141 23307
rect 17175 23273 17187 23307
rect 17129 23267 17187 23273
rect 14734 23236 14740 23248
rect 14568 23208 14740 23236
rect 12434 23109 12440 23112
rect 11885 23103 11943 23109
rect 11885 23069 11897 23103
rect 11931 23069 11943 23103
rect 11885 23063 11943 23069
rect 11978 23103 12036 23109
rect 11978 23069 11990 23103
rect 12024 23069 12036 23103
rect 11978 23063 12036 23069
rect 12161 23103 12219 23109
rect 12161 23069 12173 23103
rect 12207 23069 12219 23103
rect 12391 23103 12440 23109
rect 12391 23100 12403 23103
rect 12347 23072 12403 23100
rect 12161 23063 12219 23069
rect 12391 23069 12403 23072
rect 12437 23069 12440 23103
rect 12391 23063 12440 23069
rect 11900 23032 11928 23063
rect 12434 23060 12440 23063
rect 12492 23060 12498 23112
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13078 23100 13084 23112
rect 13035 23072 13084 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 13262 23060 13268 23112
rect 13320 23060 13326 23112
rect 14568 23109 14596 23208
rect 14734 23196 14740 23208
rect 14792 23236 14798 23248
rect 17144 23236 17172 23267
rect 17218 23264 17224 23316
rect 17276 23304 17282 23316
rect 17589 23307 17647 23313
rect 17589 23304 17601 23307
rect 17276 23276 17601 23304
rect 17276 23264 17282 23276
rect 17589 23273 17601 23276
rect 17635 23273 17647 23307
rect 18322 23304 18328 23316
rect 17589 23267 17647 23273
rect 17696 23276 18328 23304
rect 17310 23236 17316 23248
rect 14792 23208 15332 23236
rect 17144 23208 17316 23236
rect 14792 23196 14798 23208
rect 15304 23168 15332 23208
rect 17310 23196 17316 23208
rect 17368 23196 17374 23248
rect 17221 23171 17279 23177
rect 17221 23168 17233 23171
rect 15304 23140 17233 23168
rect 17221 23137 17233 23140
rect 17267 23168 17279 23171
rect 17696 23168 17724 23276
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 18509 23307 18567 23313
rect 18509 23273 18521 23307
rect 18555 23304 18567 23307
rect 18966 23304 18972 23316
rect 18555 23276 18972 23304
rect 18555 23273 18567 23276
rect 18509 23267 18567 23273
rect 18966 23264 18972 23276
rect 19024 23304 19030 23316
rect 19242 23304 19248 23316
rect 19024 23276 19248 23304
rect 19024 23264 19030 23276
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 19886 23264 19892 23316
rect 19944 23264 19950 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 21358 23304 21364 23316
rect 20128 23276 21364 23304
rect 20128 23264 20134 23276
rect 21358 23264 21364 23276
rect 21416 23304 21422 23316
rect 21416 23276 21680 23304
rect 21416 23264 21422 23276
rect 19610 23236 19616 23248
rect 17267 23140 17724 23168
rect 17972 23208 19616 23236
rect 17267 23137 17279 23140
rect 17221 23131 17279 23137
rect 14553 23103 14611 23109
rect 14553 23069 14565 23103
rect 14599 23069 14611 23103
rect 14553 23063 14611 23069
rect 15102 23060 15108 23112
rect 15160 23060 15166 23112
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17405 23103 17463 23109
rect 17405 23100 17417 23103
rect 16816 23072 17417 23100
rect 16816 23060 16822 23072
rect 17405 23069 17417 23072
rect 17451 23069 17463 23103
rect 17405 23063 17463 23069
rect 17770 23060 17776 23112
rect 17828 23060 17834 23112
rect 10796 23004 11192 23032
rect 11900 23004 12204 23032
rect 6362 22964 6368 22976
rect 5552 22936 6368 22964
rect 6362 22924 6368 22936
rect 6420 22924 6426 22976
rect 6546 22924 6552 22976
rect 6604 22964 6610 22976
rect 6641 22967 6699 22973
rect 6641 22964 6653 22967
rect 6604 22936 6653 22964
rect 6604 22924 6610 22936
rect 6641 22933 6653 22936
rect 6687 22933 6699 22967
rect 6641 22927 6699 22933
rect 6914 22924 6920 22976
rect 6972 22924 6978 22976
rect 7558 22924 7564 22976
rect 7616 22924 7622 22976
rect 7650 22924 7656 22976
rect 7708 22964 7714 22976
rect 8110 22964 8116 22976
rect 7708 22936 8116 22964
rect 7708 22924 7714 22936
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 8297 22967 8355 22973
rect 8297 22964 8309 22967
rect 8260 22936 8309 22964
rect 8260 22924 8266 22936
rect 8297 22933 8309 22936
rect 8343 22933 8355 22967
rect 8297 22927 8355 22933
rect 10689 22967 10747 22973
rect 10689 22933 10701 22967
rect 10735 22964 10747 22967
rect 10778 22964 10784 22976
rect 10735 22936 10784 22964
rect 10735 22933 10747 22936
rect 10689 22927 10747 22933
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 10873 22967 10931 22973
rect 10873 22933 10885 22967
rect 10919 22964 10931 22967
rect 11054 22964 11060 22976
rect 10919 22936 11060 22964
rect 10919 22933 10931 22936
rect 10873 22927 10931 22933
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 11164 22964 11192 23004
rect 12066 22964 12072 22976
rect 11164 22936 12072 22964
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 12176 22964 12204 23004
rect 12250 22992 12256 23044
rect 12308 23032 12314 23044
rect 12308 23004 12350 23032
rect 12406 23004 12655 23032
rect 12308 22992 12314 23004
rect 12406 22964 12434 23004
rect 12176 22936 12434 22964
rect 12526 22924 12532 22976
rect 12584 22924 12590 22976
rect 12627 22964 12655 23004
rect 12802 22992 12808 23044
rect 12860 22992 12866 23044
rect 12894 22992 12900 23044
rect 12952 22992 12958 23044
rect 13354 22992 13360 23044
rect 13412 23032 13418 23044
rect 13541 23035 13599 23041
rect 13541 23032 13553 23035
rect 13412 23004 13553 23032
rect 13412 22992 13418 23004
rect 13541 23001 13553 23004
rect 13587 23001 13599 23035
rect 13541 22995 13599 23001
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 14056 23004 14381 23032
rect 14056 22992 14062 23004
rect 14369 23001 14381 23004
rect 14415 23032 14427 23035
rect 15120 23032 15148 23060
rect 14415 23004 15148 23032
rect 14415 23001 14427 23004
rect 14369 22995 14427 23001
rect 16574 22992 16580 23044
rect 16632 23032 16638 23044
rect 17034 23032 17040 23044
rect 16632 23004 17040 23032
rect 16632 22992 16638 23004
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 17129 23035 17187 23041
rect 17129 23001 17141 23035
rect 17175 23032 17187 23035
rect 17972 23032 18000 23208
rect 19610 23196 19616 23208
rect 19668 23196 19674 23248
rect 20438 23236 20444 23248
rect 19720 23208 20444 23236
rect 19720 23168 19748 23208
rect 20438 23196 20444 23208
rect 20496 23196 20502 23248
rect 20714 23196 20720 23248
rect 20772 23196 20778 23248
rect 21542 23236 21548 23248
rect 21008 23208 21548 23236
rect 20732 23168 20760 23196
rect 18064 23140 18644 23168
rect 18064 23109 18092 23140
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 18233 23103 18291 23109
rect 18233 23100 18245 23103
rect 18095 23072 18245 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 18233 23069 18245 23072
rect 18279 23069 18291 23103
rect 18233 23063 18291 23069
rect 18414 23060 18420 23112
rect 18472 23109 18478 23112
rect 18472 23103 18487 23109
rect 18475 23100 18487 23103
rect 18475 23072 18552 23100
rect 18475 23069 18487 23072
rect 18472 23063 18487 23069
rect 18472 23060 18478 23063
rect 17175 23004 18000 23032
rect 17175 23001 17187 23004
rect 17129 22995 17187 23001
rect 18322 22992 18328 23044
rect 18380 22992 18386 23044
rect 18524 23041 18552 23072
rect 18509 23035 18567 23041
rect 18509 23001 18521 23035
rect 18555 23001 18567 23035
rect 18616 23032 18644 23140
rect 18708 23140 19748 23168
rect 20364 23140 20760 23168
rect 18708 23109 18736 23140
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23069 18751 23103
rect 18693 23063 18751 23069
rect 18782 23060 18788 23112
rect 18840 23060 18846 23112
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19061 23103 19119 23109
rect 19061 23069 19073 23103
rect 19107 23094 19119 23103
rect 19260 23094 19288 23140
rect 19107 23069 19288 23094
rect 19061 23066 19288 23069
rect 19061 23063 19119 23066
rect 18800 23032 18828 23060
rect 18616 23004 18828 23032
rect 18892 23032 18920 23063
rect 19334 23060 19340 23112
rect 19392 23060 19398 23112
rect 19886 23060 19892 23112
rect 19944 23100 19950 23112
rect 19981 23103 20039 23109
rect 19981 23100 19993 23103
rect 19944 23072 19993 23100
rect 19944 23060 19950 23072
rect 19981 23069 19993 23072
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 20162 23060 20168 23112
rect 20220 23060 20226 23112
rect 20364 23109 20392 23140
rect 20530 23109 20536 23112
rect 20349 23103 20407 23109
rect 20349 23069 20361 23103
rect 20395 23069 20407 23103
rect 20349 23063 20407 23069
rect 20487 23103 20536 23109
rect 20487 23069 20499 23103
rect 20533 23069 20536 23103
rect 20487 23063 20536 23069
rect 20364 23032 20392 23063
rect 20530 23060 20536 23063
rect 20588 23060 20594 23112
rect 20622 23060 20628 23112
rect 20680 23060 20686 23112
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20809 23103 20867 23109
rect 20809 23069 20821 23103
rect 20855 23100 20867 23103
rect 20898 23100 20904 23112
rect 20855 23072 20904 23100
rect 20855 23069 20867 23072
rect 20809 23063 20867 23069
rect 20732 23032 20760 23063
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21008 23109 21036 23208
rect 21542 23196 21548 23208
rect 21600 23196 21606 23248
rect 21652 23168 21680 23276
rect 21910 23264 21916 23316
rect 21968 23264 21974 23316
rect 22097 23307 22155 23313
rect 22097 23273 22109 23307
rect 22143 23273 22155 23307
rect 22097 23267 22155 23273
rect 22281 23307 22339 23313
rect 22281 23273 22293 23307
rect 22327 23304 22339 23307
rect 22922 23304 22928 23316
rect 22327 23276 22928 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 21928 23168 21956 23264
rect 22112 23236 22140 23267
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 23290 23264 23296 23316
rect 23348 23304 23354 23316
rect 23934 23304 23940 23316
rect 23348 23276 23940 23304
rect 23348 23264 23354 23276
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 25130 23264 25136 23316
rect 25188 23304 25194 23316
rect 27338 23304 27344 23316
rect 25188 23276 27344 23304
rect 25188 23264 25194 23276
rect 27338 23264 27344 23276
rect 27396 23264 27402 23316
rect 28074 23264 28080 23316
rect 28132 23264 28138 23316
rect 32398 23264 32404 23316
rect 32456 23264 32462 23316
rect 32493 23307 32551 23313
rect 32493 23273 32505 23307
rect 32539 23304 32551 23307
rect 33134 23304 33140 23316
rect 32539 23276 33140 23304
rect 32539 23273 32551 23276
rect 32493 23267 32551 23273
rect 33134 23264 33140 23276
rect 33192 23264 33198 23316
rect 33594 23264 33600 23316
rect 33652 23264 33658 23316
rect 22112 23208 22324 23236
rect 22296 23180 22324 23208
rect 24872 23208 25176 23236
rect 21652 23140 21772 23168
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21174 23060 21180 23112
rect 21232 23100 21238 23112
rect 21545 23103 21603 23109
rect 21545 23100 21557 23103
rect 21232 23072 21557 23100
rect 21232 23060 21238 23072
rect 21545 23069 21557 23072
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21744 23109 21772 23140
rect 21836 23140 21956 23168
rect 21836 23109 21864 23140
rect 22278 23128 22284 23180
rect 22336 23128 22342 23180
rect 24872 23168 24900 23208
rect 22664 23140 24900 23168
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 21910 23060 21916 23112
rect 21968 23100 21974 23112
rect 22664 23109 22692 23140
rect 25038 23128 25044 23180
rect 25096 23128 25102 23180
rect 25148 23168 25176 23208
rect 25406 23196 25412 23248
rect 25464 23236 25470 23248
rect 28092 23236 28120 23264
rect 32416 23236 32444 23264
rect 32677 23239 32735 23245
rect 32677 23236 32689 23239
rect 25464 23208 26188 23236
rect 25464 23196 25470 23208
rect 26050 23168 26056 23180
rect 25148 23140 26056 23168
rect 26050 23128 26056 23140
rect 26108 23128 26114 23180
rect 26160 23168 26188 23208
rect 27632 23208 28120 23236
rect 28276 23208 28856 23236
rect 32416 23208 32689 23236
rect 27632 23177 27660 23208
rect 27617 23171 27675 23177
rect 26160 23140 26832 23168
rect 22005 23103 22063 23109
rect 22005 23100 22017 23103
rect 21968 23072 22017 23100
rect 21968 23060 21974 23072
rect 22005 23069 22017 23072
rect 22051 23069 22063 23103
rect 22005 23063 22063 23069
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23069 22707 23103
rect 22649 23063 22707 23069
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23100 23259 23103
rect 23474 23100 23480 23112
rect 23247 23072 23480 23100
rect 23247 23069 23259 23072
rect 23201 23063 23259 23069
rect 21928 23032 21956 23060
rect 18892 23004 19304 23032
rect 18509 22995 18567 23001
rect 13173 22967 13231 22973
rect 13173 22964 13185 22967
rect 12627 22936 13185 22964
rect 13173 22933 13185 22936
rect 13219 22933 13231 22967
rect 13173 22927 13231 22933
rect 14645 22967 14703 22973
rect 14645 22933 14657 22967
rect 14691 22964 14703 22967
rect 15194 22964 15200 22976
rect 14691 22936 15200 22964
rect 14691 22933 14703 22936
rect 14645 22927 14703 22933
rect 15194 22924 15200 22936
rect 15252 22924 15258 22976
rect 15381 22967 15439 22973
rect 15381 22933 15393 22967
rect 15427 22964 15439 22967
rect 15562 22964 15568 22976
rect 15427 22936 15568 22964
rect 15427 22933 15439 22936
rect 15381 22927 15439 22933
rect 15562 22924 15568 22936
rect 15620 22964 15626 22976
rect 17310 22964 17316 22976
rect 15620 22936 17316 22964
rect 15620 22924 15626 22936
rect 17310 22924 17316 22936
rect 17368 22924 17374 22976
rect 17494 22924 17500 22976
rect 17552 22964 17558 22976
rect 17865 22967 17923 22973
rect 17865 22964 17877 22967
rect 17552 22936 17877 22964
rect 17552 22924 17558 22936
rect 17865 22933 17877 22936
rect 17911 22933 17923 22967
rect 17865 22927 17923 22933
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18104 22936 18981 22964
rect 18104 22924 18110 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 19276 22964 19304 23004
rect 19966 23004 20392 23032
rect 20456 23004 21956 23032
rect 19966 22964 19994 23004
rect 19276 22936 19994 22964
rect 20073 22967 20131 22973
rect 18969 22927 19027 22933
rect 20073 22933 20085 22967
rect 20119 22964 20131 22967
rect 20456 22964 20484 23004
rect 20119 22936 20484 22964
rect 20119 22933 20131 22936
rect 20073 22927 20131 22933
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 21177 22967 21235 22973
rect 21177 22964 21189 22967
rect 20588 22936 21189 22964
rect 20588 22924 20594 22936
rect 21177 22933 21189 22936
rect 21223 22933 21235 22967
rect 21177 22927 21235 22933
rect 21266 22924 21272 22976
rect 21324 22964 21330 22976
rect 21726 22964 21732 22976
rect 21324 22936 21732 22964
rect 21324 22924 21330 22936
rect 21726 22924 21732 22936
rect 21784 22924 21790 22976
rect 22002 22924 22008 22976
rect 22060 22964 22066 22976
rect 22112 22964 22140 23063
rect 23474 23060 23480 23072
rect 23532 23060 23538 23112
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23069 23719 23103
rect 25133 23103 25191 23109
rect 25133 23100 25145 23103
rect 23661 23063 23719 23069
rect 24964 23072 25145 23100
rect 23676 23032 23704 23063
rect 24964 23044 24992 23072
rect 25133 23069 25145 23072
rect 25179 23100 25191 23103
rect 25682 23100 25688 23112
rect 25179 23072 25688 23100
rect 25179 23069 25191 23072
rect 25133 23063 25191 23069
rect 25682 23060 25688 23072
rect 25740 23060 25746 23112
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23069 25835 23103
rect 25777 23063 25835 23069
rect 23308 23004 23704 23032
rect 23937 23035 23995 23041
rect 23308 22976 23336 23004
rect 23937 23001 23949 23035
rect 23983 23032 23995 23035
rect 24118 23032 24124 23044
rect 23983 23004 24124 23032
rect 23983 23001 23995 23004
rect 23937 22995 23995 23001
rect 22060 22936 22140 22964
rect 22925 22967 22983 22973
rect 22060 22924 22066 22936
rect 22925 22933 22937 22967
rect 22971 22964 22983 22967
rect 23106 22964 23112 22976
rect 22971 22936 23112 22964
rect 22971 22933 22983 22936
rect 22925 22927 22983 22933
rect 23106 22924 23112 22936
rect 23164 22924 23170 22976
rect 23290 22924 23296 22976
rect 23348 22924 23354 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 23952 22964 23980 22995
rect 24118 22992 24124 23004
rect 24176 23032 24182 23044
rect 24762 23032 24768 23044
rect 24176 23004 24768 23032
rect 24176 22992 24182 23004
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 24854 22992 24860 23044
rect 24912 22992 24918 23044
rect 24946 22992 24952 23044
rect 25004 22992 25010 23044
rect 25792 23032 25820 23063
rect 25866 23060 25872 23112
rect 25924 23100 25930 23112
rect 25924 23072 25969 23100
rect 25924 23060 25930 23072
rect 26068 23041 26096 23128
rect 26160 23109 26188 23140
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 26283 23103 26341 23109
rect 26283 23069 26295 23103
rect 26329 23100 26341 23103
rect 26418 23100 26424 23112
rect 26329 23072 26424 23100
rect 26329 23069 26341 23072
rect 26283 23063 26341 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 26513 23103 26571 23109
rect 26513 23069 26525 23103
rect 26559 23100 26571 23103
rect 26602 23100 26608 23112
rect 26559 23072 26608 23100
rect 26559 23069 26571 23072
rect 26513 23063 26571 23069
rect 26602 23060 26608 23072
rect 26660 23060 26666 23112
rect 26694 23060 26700 23112
rect 26752 23060 26758 23112
rect 26804 23109 26832 23140
rect 27617 23137 27629 23171
rect 27663 23137 27675 23171
rect 28276 23168 28304 23208
rect 27617 23131 27675 23137
rect 28000 23140 28304 23168
rect 28353 23171 28411 23177
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23100 26939 23103
rect 26970 23100 26976 23112
rect 26927 23072 26976 23100
rect 26927 23069 26939 23072
rect 26881 23063 26939 23069
rect 26970 23060 26976 23072
rect 27028 23100 27034 23112
rect 27430 23100 27436 23112
rect 27028 23072 27436 23100
rect 27028 23060 27034 23072
rect 27430 23060 27436 23072
rect 27488 23100 27494 23112
rect 27798 23100 27804 23112
rect 27488 23072 27804 23100
rect 27488 23060 27494 23072
rect 27798 23060 27804 23072
rect 27856 23100 27862 23112
rect 28000 23109 28028 23140
rect 28353 23137 28365 23171
rect 28399 23168 28411 23171
rect 28534 23168 28540 23180
rect 28399 23140 28540 23168
rect 28399 23137 28411 23140
rect 28353 23131 28411 23137
rect 28534 23128 28540 23140
rect 28592 23128 28598 23180
rect 28828 23177 28856 23208
rect 32677 23205 32689 23208
rect 32723 23205 32735 23239
rect 32677 23199 32735 23205
rect 33045 23239 33103 23245
rect 33045 23205 33057 23239
rect 33091 23236 33103 23239
rect 33612 23236 33640 23264
rect 33091 23208 33640 23236
rect 33091 23205 33103 23208
rect 33045 23199 33103 23205
rect 28813 23171 28871 23177
rect 28813 23137 28825 23171
rect 28859 23137 28871 23171
rect 28813 23131 28871 23137
rect 32306 23128 32312 23180
rect 32364 23168 32370 23180
rect 32401 23171 32459 23177
rect 32401 23168 32413 23171
rect 32364 23140 32413 23168
rect 32364 23128 32370 23140
rect 32401 23137 32413 23140
rect 32447 23137 32459 23171
rect 32401 23131 32459 23137
rect 27985 23103 28043 23109
rect 27985 23100 27997 23103
rect 27856 23072 27997 23100
rect 27856 23060 27862 23072
rect 27985 23069 27997 23072
rect 28031 23069 28043 23103
rect 27985 23063 28043 23069
rect 28077 23103 28135 23109
rect 28077 23069 28089 23103
rect 28123 23100 28135 23103
rect 28258 23100 28264 23112
rect 28123 23072 28264 23100
rect 28123 23069 28135 23072
rect 28077 23063 28135 23069
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 28721 23103 28779 23109
rect 28721 23100 28733 23103
rect 28368 23072 28733 23100
rect 26053 23035 26111 23041
rect 25792 23004 25912 23032
rect 23624 22936 23980 22964
rect 23624 22924 23630 22936
rect 25130 22924 25136 22976
rect 25188 22964 25194 22976
rect 25317 22967 25375 22973
rect 25317 22964 25329 22967
rect 25188 22936 25329 22964
rect 25188 22924 25194 22936
rect 25317 22933 25329 22936
rect 25363 22933 25375 22967
rect 25884 22964 25912 23004
rect 26053 23001 26065 23035
rect 26099 23001 26111 23035
rect 26053 22995 26111 23001
rect 28368 22976 28396 23072
rect 28721 23069 28733 23072
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 32125 23103 32183 23109
rect 32125 23069 32137 23103
rect 32171 23100 32183 23103
rect 33060 23100 33088 23199
rect 32171 23072 33088 23100
rect 32171 23069 32183 23072
rect 32125 23063 32183 23069
rect 26234 22964 26240 22976
rect 25884 22936 26240 22964
rect 25317 22927 25375 22933
rect 26234 22924 26240 22936
rect 26292 22924 26298 22976
rect 26418 22924 26424 22976
rect 26476 22924 26482 22976
rect 27065 22967 27123 22973
rect 27065 22933 27077 22967
rect 27111 22964 27123 22967
rect 27154 22964 27160 22976
rect 27111 22936 27160 22964
rect 27111 22933 27123 22936
rect 27065 22927 27123 22933
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 28261 22967 28319 22973
rect 28261 22964 28273 22967
rect 27764 22936 28273 22964
rect 27764 22924 27770 22936
rect 28261 22933 28273 22936
rect 28307 22933 28319 22967
rect 28261 22927 28319 22933
rect 28350 22924 28356 22976
rect 28408 22924 28414 22976
rect 28442 22924 28448 22976
rect 28500 22964 28506 22976
rect 28997 22967 29055 22973
rect 28997 22964 29009 22967
rect 28500 22936 29009 22964
rect 28500 22924 28506 22936
rect 28997 22933 29009 22936
rect 29043 22933 29055 22967
rect 28997 22927 29055 22933
rect 1104 22874 43884 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 43884 22874
rect 1104 22800 43884 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3513 22763 3571 22769
rect 3513 22760 3525 22763
rect 3200 22732 3525 22760
rect 3200 22720 3206 22732
rect 3513 22729 3525 22732
rect 3559 22729 3571 22763
rect 3513 22723 3571 22729
rect 3878 22720 3884 22772
rect 3936 22760 3942 22772
rect 6546 22760 6552 22772
rect 3936 22732 6552 22760
rect 3936 22720 3942 22732
rect 3970 22652 3976 22704
rect 4028 22692 4034 22704
rect 4028 22664 4661 22692
rect 4028 22652 4034 22664
rect 1664 22627 1722 22633
rect 1664 22593 1676 22627
rect 1710 22624 1722 22627
rect 3878 22624 3884 22636
rect 1710 22596 3884 22624
rect 1710 22593 1722 22596
rect 1664 22587 1722 22593
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 4633 22633 4661 22664
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22593 4583 22627
rect 4525 22587 4583 22593
rect 4618 22627 4676 22633
rect 4618 22593 4630 22627
rect 4664 22593 4676 22627
rect 4618 22587 4676 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 1412 22420 1440 22519
rect 2958 22516 2964 22568
rect 3016 22516 3022 22568
rect 3694 22516 3700 22568
rect 3752 22516 3758 22568
rect 4540 22556 4568 22587
rect 4724 22556 4752 22732
rect 6546 22720 6552 22732
rect 6604 22720 6610 22772
rect 8941 22763 8999 22769
rect 6656 22732 7328 22760
rect 6656 22704 6684 22732
rect 5644 22664 6592 22692
rect 5644 22636 5672 22664
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 5074 22633 5080 22636
rect 4893 22627 4951 22633
rect 4893 22593 4905 22627
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 5031 22627 5080 22633
rect 5031 22593 5043 22627
rect 5077 22593 5080 22627
rect 5031 22587 5080 22593
rect 4540 22528 4752 22556
rect 4908 22556 4936 22587
rect 5074 22584 5080 22587
rect 5132 22584 5138 22636
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 5626 22584 5632 22636
rect 5684 22584 5690 22636
rect 5718 22584 5724 22636
rect 5776 22624 5782 22636
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5776 22596 5825 22624
rect 5776 22584 5782 22596
rect 5813 22593 5825 22596
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 5902 22584 5908 22636
rect 5960 22584 5966 22636
rect 5997 22627 6055 22633
rect 5997 22593 6009 22627
rect 6043 22624 6055 22627
rect 6270 22624 6276 22636
rect 6043 22596 6276 22624
rect 6043 22593 6055 22596
rect 5997 22587 6055 22593
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 6564 22624 6592 22664
rect 6638 22652 6644 22704
rect 6696 22652 6702 22704
rect 7190 22652 7196 22704
rect 7248 22652 7254 22704
rect 7300 22701 7328 22732
rect 7576 22732 8202 22760
rect 7285 22695 7343 22701
rect 7285 22661 7297 22695
rect 7331 22661 7343 22695
rect 7285 22655 7343 22661
rect 6822 22624 6828 22636
rect 6564 22596 6828 22624
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 6914 22584 6920 22636
rect 6972 22584 6978 22636
rect 7098 22634 7104 22636
rect 7025 22633 7104 22634
rect 7010 22627 7104 22633
rect 7010 22593 7022 22627
rect 7056 22606 7104 22627
rect 7056 22593 7068 22606
rect 7010 22587 7068 22593
rect 7098 22584 7104 22606
rect 7156 22624 7162 22636
rect 7156 22596 7328 22624
rect 7156 22584 7162 22596
rect 6638 22556 6644 22568
rect 4908 22528 6644 22556
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7300 22556 7328 22596
rect 7374 22584 7380 22636
rect 7432 22633 7438 22636
rect 7432 22627 7481 22633
rect 7432 22593 7435 22627
rect 7469 22624 7481 22627
rect 7576 22624 7604 22732
rect 7926 22652 7932 22704
rect 7984 22652 7990 22704
rect 8018 22652 8024 22704
rect 8076 22652 8082 22704
rect 8174 22692 8202 22732
rect 8941 22729 8953 22763
rect 8987 22760 8999 22763
rect 8987 22732 10272 22760
rect 8987 22729 8999 22732
rect 8941 22723 8999 22729
rect 9309 22695 9367 22701
rect 8174 22664 8892 22692
rect 7469 22596 7604 22624
rect 7469 22593 7481 22596
rect 7432 22587 7481 22593
rect 7432 22584 7438 22587
rect 7650 22584 7656 22636
rect 7708 22584 7714 22636
rect 8174 22633 8202 22664
rect 8864 22636 8892 22664
rect 9309 22661 9321 22695
rect 9355 22692 9367 22695
rect 10042 22692 10048 22704
rect 9355 22664 10048 22692
rect 9355 22661 9367 22664
rect 9309 22655 9367 22661
rect 10042 22652 10048 22664
rect 10100 22652 10106 22704
rect 10244 22692 10272 22732
rect 10318 22720 10324 22772
rect 10376 22720 10382 22772
rect 10870 22760 10876 22772
rect 10520 22732 10876 22760
rect 10520 22692 10548 22732
rect 10870 22720 10876 22732
rect 10928 22720 10934 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 12342 22760 12348 22772
rect 11112 22732 12348 22760
rect 11112 22720 11118 22732
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 13173 22763 13231 22769
rect 13173 22729 13185 22763
rect 13219 22760 13231 22763
rect 13262 22760 13268 22772
rect 13219 22732 13268 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13262 22720 13268 22732
rect 13320 22760 13326 22772
rect 13814 22760 13820 22772
rect 13320 22732 13820 22760
rect 13320 22720 13326 22732
rect 13814 22720 13820 22732
rect 13872 22720 13878 22772
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15378 22760 15384 22772
rect 15160 22732 15384 22760
rect 15160 22720 15166 22732
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 15565 22763 15623 22769
rect 15565 22729 15577 22763
rect 15611 22760 15623 22763
rect 15838 22760 15844 22772
rect 15611 22732 15844 22760
rect 15611 22729 15623 22732
rect 15565 22723 15623 22729
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 16114 22720 16120 22772
rect 16172 22760 16178 22772
rect 17313 22763 17371 22769
rect 17313 22760 17325 22763
rect 16172 22732 17325 22760
rect 16172 22720 16178 22732
rect 17313 22729 17325 22732
rect 17359 22729 17371 22763
rect 17313 22723 17371 22729
rect 18046 22720 18052 22772
rect 18104 22720 18110 22772
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 19242 22760 19248 22772
rect 19116 22732 19248 22760
rect 19116 22720 19122 22732
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 19518 22720 19524 22772
rect 19576 22760 19582 22772
rect 19889 22763 19947 22769
rect 19889 22760 19901 22763
rect 19576 22732 19901 22760
rect 19576 22720 19582 22732
rect 19889 22729 19901 22732
rect 19935 22760 19947 22763
rect 20162 22760 20168 22772
rect 19935 22732 20168 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 20714 22760 20720 22772
rect 20272 22732 20720 22760
rect 11238 22692 11244 22704
rect 10244 22664 10548 22692
rect 10612 22664 11244 22692
rect 7801 22627 7859 22633
rect 7801 22593 7813 22627
rect 7847 22624 7859 22627
rect 8159 22627 8217 22633
rect 7847 22596 7972 22624
rect 7847 22593 7859 22596
rect 7801 22587 7859 22593
rect 7944 22556 7972 22596
rect 8159 22593 8171 22627
rect 8205 22593 8217 22627
rect 8159 22587 8217 22593
rect 8478 22584 8484 22636
rect 8536 22624 8542 22636
rect 8757 22627 8815 22633
rect 8757 22624 8769 22627
rect 8536 22596 8769 22624
rect 8536 22584 8542 22596
rect 8757 22593 8769 22596
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 7300 22528 7972 22556
rect 2777 22491 2835 22497
rect 2777 22457 2789 22491
rect 2823 22488 2835 22491
rect 3142 22488 3148 22500
rect 2823 22460 3148 22488
rect 2823 22457 2835 22460
rect 2777 22451 2835 22457
rect 3142 22448 3148 22460
rect 3200 22488 3206 22500
rect 3712 22488 3740 22516
rect 3200 22460 3740 22488
rect 3200 22448 3206 22460
rect 4062 22448 4068 22500
rect 4120 22488 4126 22500
rect 4120 22460 5212 22488
rect 4120 22448 4126 22460
rect 1762 22420 1768 22432
rect 1412 22392 1768 22420
rect 1762 22380 1768 22392
rect 1820 22380 1826 22432
rect 2406 22380 2412 22432
rect 2464 22420 2470 22432
rect 4249 22423 4307 22429
rect 4249 22420 4261 22423
rect 2464 22392 4261 22420
rect 2464 22380 2470 22392
rect 4249 22389 4261 22392
rect 4295 22420 4307 22423
rect 4890 22420 4896 22432
rect 4295 22392 4896 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4890 22380 4896 22392
rect 4948 22380 4954 22432
rect 5184 22429 5212 22460
rect 5442 22448 5448 22500
rect 5500 22488 5506 22500
rect 5994 22488 6000 22500
rect 5500 22460 6000 22488
rect 5500 22448 5506 22460
rect 5994 22448 6000 22460
rect 6052 22448 6058 22500
rect 6822 22448 6828 22500
rect 6880 22488 6886 22500
rect 7834 22488 7840 22500
rect 6880 22460 7840 22488
rect 6880 22448 6886 22460
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 7944 22488 7972 22528
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22556 8723 22559
rect 8956 22556 8984 22587
rect 9030 22584 9036 22636
rect 9088 22584 9094 22636
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9217 22627 9275 22633
rect 9217 22624 9229 22627
rect 9180 22596 9229 22624
rect 9180 22584 9186 22596
rect 9217 22593 9229 22596
rect 9263 22593 9275 22627
rect 9217 22587 9275 22593
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 9490 22584 9496 22636
rect 9548 22584 9554 22636
rect 10612 22633 10640 22664
rect 11238 22652 11244 22664
rect 11296 22692 11302 22704
rect 12161 22695 12219 22701
rect 12161 22692 12173 22695
rect 11296 22664 12173 22692
rect 11296 22652 11302 22664
rect 12161 22661 12173 22664
rect 12207 22661 12219 22695
rect 12161 22655 12219 22661
rect 12802 22652 12808 22704
rect 12860 22692 12866 22704
rect 17954 22692 17960 22704
rect 12860 22664 17960 22692
rect 12860 22652 12866 22664
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 9600 22596 10425 22624
rect 9508 22556 9536 22584
rect 8711 22528 9536 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 9600 22497 9628 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10413 22587 10471 22593
rect 10561 22627 10640 22633
rect 10561 22593 10573 22627
rect 10607 22596 10640 22627
rect 10689 22627 10747 22633
rect 10607 22593 10619 22596
rect 10561 22587 10619 22593
rect 10689 22593 10701 22627
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 10704 22556 10732 22587
rect 10778 22584 10784 22636
rect 10836 22584 10842 22636
rect 10878 22627 10936 22633
rect 10878 22593 10890 22627
rect 10924 22593 10936 22627
rect 10878 22587 10936 22593
rect 10612 22528 10732 22556
rect 10612 22500 10640 22528
rect 9585 22491 9643 22497
rect 7944 22460 9168 22488
rect 9140 22432 9168 22460
rect 9585 22457 9597 22491
rect 9631 22457 9643 22491
rect 9585 22451 9643 22457
rect 10226 22448 10232 22500
rect 10284 22488 10290 22500
rect 10594 22488 10600 22500
rect 10284 22460 10600 22488
rect 10284 22448 10290 22460
rect 10594 22448 10600 22460
rect 10652 22448 10658 22500
rect 5169 22423 5227 22429
rect 5169 22389 5181 22423
rect 5215 22389 5227 22423
rect 5169 22383 5227 22389
rect 6086 22380 6092 22432
rect 6144 22420 6150 22432
rect 6181 22423 6239 22429
rect 6181 22420 6193 22423
rect 6144 22392 6193 22420
rect 6144 22380 6150 22392
rect 6181 22389 6193 22392
rect 6227 22389 6239 22423
rect 6181 22383 6239 22389
rect 6730 22380 6736 22432
rect 6788 22420 6794 22432
rect 7006 22420 7012 22432
rect 6788 22392 7012 22420
rect 6788 22380 6794 22392
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 7558 22380 7564 22432
rect 7616 22380 7622 22432
rect 8294 22380 8300 22432
rect 8352 22380 8358 22432
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 9950 22420 9956 22432
rect 9732 22392 9956 22420
rect 9732 22380 9738 22392
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 10893 22420 10921 22587
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 12621 22627 12679 22633
rect 12621 22624 12633 22627
rect 11204 22596 12633 22624
rect 11204 22584 11210 22596
rect 12621 22593 12633 22596
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11020 22528 11529 22556
rect 11020 22516 11026 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11517 22519 11575 22525
rect 11606 22516 11612 22568
rect 11664 22556 11670 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11664 22528 12449 22556
rect 11664 22516 11670 22528
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 12529 22559 12587 22565
rect 12529 22525 12541 22559
rect 12575 22525 12587 22559
rect 12529 22519 12587 22525
rect 12342 22448 12348 22500
rect 12400 22488 12406 22500
rect 12544 22488 12572 22519
rect 12710 22516 12716 22568
rect 12768 22516 12774 22568
rect 13372 22500 13400 22587
rect 13722 22584 13728 22636
rect 13780 22584 13786 22636
rect 13906 22584 13912 22636
rect 13964 22584 13970 22636
rect 14476 22633 14504 22664
rect 17954 22652 17960 22664
rect 18012 22652 18018 22704
rect 18064 22692 18092 22720
rect 18693 22695 18751 22701
rect 18064 22664 18276 22692
rect 14461 22627 14519 22633
rect 14461 22593 14473 22627
rect 14507 22593 14519 22627
rect 14461 22587 14519 22593
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 14734 22584 14740 22636
rect 14792 22584 14798 22636
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15010 22624 15016 22636
rect 14967 22596 15016 22624
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22593 15531 22627
rect 15473 22587 15531 22593
rect 13630 22516 13636 22568
rect 13688 22556 13694 22568
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 13688 22528 15117 22556
rect 13688 22516 13694 22528
rect 15105 22525 15117 22528
rect 15151 22525 15163 22559
rect 15105 22519 15163 22525
rect 15378 22516 15384 22568
rect 15436 22556 15442 22568
rect 15488 22556 15516 22587
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 15620 22596 15669 22624
rect 15620 22584 15626 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 15657 22587 15715 22593
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16390 22624 16396 22636
rect 16071 22596 16396 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16040 22556 16068 22587
rect 16390 22584 16396 22596
rect 16448 22584 16454 22636
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22624 16727 22627
rect 17218 22624 17224 22636
rect 16715 22596 17224 22624
rect 16715 22593 16727 22596
rect 16669 22587 16727 22593
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 17678 22584 17684 22636
rect 17736 22584 17742 22636
rect 18248 22633 18276 22664
rect 18693 22661 18705 22695
rect 18739 22692 18751 22695
rect 18739 22664 19564 22692
rect 18739 22661 18751 22664
rect 18693 22655 18751 22661
rect 19536 22636 19564 22664
rect 19610 22652 19616 22704
rect 19668 22692 19674 22704
rect 19668 22664 20116 22692
rect 19668 22652 19674 22664
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22593 18291 22627
rect 18233 22587 18291 22593
rect 15436 22528 16068 22556
rect 15436 22516 15442 22528
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17037 22559 17095 22565
rect 17037 22556 17049 22559
rect 16816 22528 17049 22556
rect 16816 22516 16822 22528
rect 17037 22525 17049 22528
rect 17083 22525 17095 22559
rect 17037 22519 17095 22525
rect 17310 22516 17316 22568
rect 17368 22516 17374 22568
rect 17696 22556 17724 22584
rect 18064 22556 18092 22587
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 18472 22596 18920 22624
rect 18472 22584 18478 22596
rect 18506 22556 18512 22568
rect 17696 22528 18512 22556
rect 18506 22516 18512 22528
rect 18564 22516 18570 22568
rect 18785 22559 18843 22565
rect 18785 22525 18797 22559
rect 18831 22525 18843 22559
rect 18785 22519 18843 22525
rect 12400 22460 12572 22488
rect 12400 22448 12406 22460
rect 13078 22448 13084 22500
rect 13136 22448 13142 22500
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 13412 22460 15516 22488
rect 13412 22448 13418 22460
rect 10376 22392 10921 22420
rect 11057 22423 11115 22429
rect 10376 22380 10382 22392
rect 11057 22389 11069 22423
rect 11103 22420 11115 22423
rect 11606 22420 11612 22432
rect 11103 22392 11612 22420
rect 11103 22389 11115 22392
rect 11057 22383 11115 22389
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 12253 22423 12311 22429
rect 12253 22420 12265 22423
rect 11848 22392 12265 22420
rect 11848 22380 11854 22392
rect 12253 22389 12265 22392
rect 12299 22389 12311 22423
rect 13096 22420 13124 22448
rect 15488 22432 15516 22460
rect 16666 22448 16672 22500
rect 16724 22488 16730 22500
rect 16945 22491 17003 22497
rect 16945 22488 16957 22491
rect 16724 22460 16957 22488
rect 16724 22448 16730 22460
rect 16945 22457 16957 22460
rect 16991 22457 17003 22491
rect 17328 22488 17356 22516
rect 18800 22488 18828 22519
rect 17328 22460 18828 22488
rect 18892 22488 18920 22596
rect 18966 22584 18972 22636
rect 19024 22584 19030 22636
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19334 22584 19340 22636
rect 19392 22584 19398 22636
rect 19426 22584 19432 22636
rect 19484 22584 19490 22636
rect 19518 22584 19524 22636
rect 19576 22584 19582 22636
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22593 19855 22627
rect 19797 22587 19855 22593
rect 19352 22556 19380 22584
rect 19812 22556 19840 22587
rect 19886 22584 19892 22636
rect 19944 22624 19950 22636
rect 20088 22633 20116 22664
rect 20272 22633 20300 22732
rect 20714 22720 20720 22732
rect 20772 22720 20778 22772
rect 21082 22720 21088 22772
rect 21140 22760 21146 22772
rect 21450 22760 21456 22772
rect 21140 22732 21456 22760
rect 21140 22720 21146 22732
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 21542 22720 21548 22772
rect 21600 22720 21606 22772
rect 23474 22720 23480 22772
rect 23532 22720 23538 22772
rect 24394 22720 24400 22772
rect 24452 22720 24458 22772
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 25961 22763 26019 22769
rect 24636 22732 24716 22760
rect 24636 22720 24642 22732
rect 20640 22664 20852 22692
rect 20640 22636 20668 22664
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19944 22596 19993 22624
rect 19944 22584 19950 22596
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 19352 22528 19840 22556
rect 20088 22556 20116 22587
rect 20346 22584 20352 22636
rect 20404 22584 20410 22636
rect 20438 22584 20444 22636
rect 20496 22624 20502 22636
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 20496 22596 20545 22624
rect 20496 22584 20502 22596
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20622 22584 20628 22636
rect 20680 22584 20686 22636
rect 20824 22633 20852 22664
rect 20916 22664 21220 22692
rect 20809 22627 20867 22633
rect 20809 22593 20821 22627
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 20916 22556 20944 22664
rect 21192 22636 21220 22664
rect 21358 22652 21364 22704
rect 21416 22652 21422 22704
rect 21821 22695 21879 22701
rect 21821 22692 21833 22695
rect 21468 22664 21833 22692
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22593 21051 22627
rect 20993 22587 21051 22593
rect 20088 22528 20944 22556
rect 21008 22556 21036 22587
rect 21082 22584 21088 22636
rect 21140 22584 21146 22636
rect 21174 22584 21180 22636
rect 21232 22584 21238 22636
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22624 21327 22627
rect 21376 22624 21404 22652
rect 21315 22596 21404 22624
rect 21315 22593 21327 22596
rect 21269 22587 21327 22593
rect 21358 22556 21364 22568
rect 21008 22528 21364 22556
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 20073 22491 20131 22497
rect 18892 22460 19748 22488
rect 16945 22451 17003 22457
rect 13906 22420 13912 22432
rect 13096 22392 13912 22420
rect 12253 22383 12311 22389
rect 13906 22380 13912 22392
rect 13964 22420 13970 22432
rect 14826 22420 14832 22432
rect 13964 22392 14832 22420
rect 13964 22380 13970 22392
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 16390 22380 16396 22432
rect 16448 22380 16454 22432
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 16834 22423 16892 22429
rect 16834 22420 16846 22423
rect 16632 22392 16846 22420
rect 16632 22380 16638 22392
rect 16834 22389 16846 22392
rect 16880 22420 16892 22423
rect 17126 22420 17132 22432
rect 16880 22392 17132 22420
rect 16880 22389 16892 22392
rect 16834 22383 16892 22389
rect 17126 22380 17132 22392
rect 17184 22380 17190 22432
rect 17586 22380 17592 22432
rect 17644 22420 17650 22432
rect 17865 22423 17923 22429
rect 17865 22420 17877 22423
rect 17644 22392 17877 22420
rect 17644 22380 17650 22392
rect 17865 22389 17877 22392
rect 17911 22389 17923 22423
rect 17865 22383 17923 22389
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18325 22423 18383 22429
rect 18325 22420 18337 22423
rect 18012 22392 18337 22420
rect 18012 22380 18018 22392
rect 18325 22389 18337 22392
rect 18371 22389 18383 22423
rect 18325 22383 18383 22389
rect 18414 22380 18420 22432
rect 18472 22420 18478 22432
rect 18690 22420 18696 22432
rect 18472 22392 18696 22420
rect 18472 22380 18478 22392
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 18782 22380 18788 22432
rect 18840 22420 18846 22432
rect 19153 22423 19211 22429
rect 19153 22420 19165 22423
rect 18840 22392 19165 22420
rect 18840 22380 18846 22392
rect 19153 22389 19165 22392
rect 19199 22389 19211 22423
rect 19153 22383 19211 22389
rect 19610 22380 19616 22432
rect 19668 22380 19674 22432
rect 19720 22420 19748 22460
rect 20073 22457 20085 22491
rect 20119 22488 20131 22491
rect 20898 22488 20904 22500
rect 20119 22460 20904 22488
rect 20119 22457 20131 22460
rect 20073 22451 20131 22457
rect 20898 22448 20904 22460
rect 20956 22448 20962 22500
rect 21082 22448 21088 22500
rect 21140 22488 21146 22500
rect 21468 22488 21496 22664
rect 21821 22661 21833 22664
rect 21867 22661 21879 22695
rect 21821 22655 21879 22661
rect 21910 22652 21916 22704
rect 21968 22692 21974 22704
rect 24412 22692 24440 22720
rect 24688 22701 24716 22732
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26007 22732 27200 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 21968 22664 23980 22692
rect 21968 22652 21974 22664
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 21818 22516 21824 22568
rect 21876 22556 21882 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21876 22528 21925 22556
rect 21876 22516 21882 22528
rect 21913 22525 21925 22528
rect 21959 22525 21971 22559
rect 22278 22556 22284 22568
rect 21913 22519 21971 22525
rect 22112 22528 22284 22556
rect 22112 22488 22140 22528
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22480 22556 22508 22587
rect 22554 22584 22560 22636
rect 22612 22624 22618 22636
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 22612 22596 22661 22624
rect 22612 22584 22618 22596
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 22738 22584 22744 22636
rect 22796 22584 22802 22636
rect 22833 22627 22891 22633
rect 22833 22593 22845 22627
rect 22879 22593 22891 22627
rect 22833 22587 22891 22593
rect 22336 22528 22508 22556
rect 22336 22516 22342 22528
rect 21140 22460 21496 22488
rect 21566 22460 22140 22488
rect 21140 22448 21146 22460
rect 20254 22420 20260 22432
rect 19720 22392 20260 22420
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 20349 22423 20407 22429
rect 20349 22389 20361 22423
rect 20395 22420 20407 22423
rect 20530 22420 20536 22432
rect 20395 22392 20536 22420
rect 20395 22389 20407 22392
rect 20349 22383 20407 22389
rect 20530 22380 20536 22392
rect 20588 22380 20594 22432
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 20809 22423 20867 22429
rect 20809 22420 20821 22423
rect 20772 22392 20821 22420
rect 20772 22380 20778 22392
rect 20809 22389 20821 22392
rect 20855 22420 20867 22423
rect 21566 22420 21594 22460
rect 22186 22448 22192 22500
rect 22244 22488 22250 22500
rect 22756 22488 22784 22584
rect 22244 22460 22784 22488
rect 22848 22556 22876 22587
rect 22922 22584 22928 22636
rect 22980 22624 22986 22636
rect 23201 22627 23259 22633
rect 23201 22624 23213 22627
rect 22980 22596 23213 22624
rect 22980 22584 22986 22596
rect 23201 22593 23213 22596
rect 23247 22593 23259 22627
rect 23201 22587 23259 22593
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 23952 22633 23980 22664
rect 24228 22664 24440 22692
rect 24673 22695 24731 22701
rect 24228 22633 24256 22664
rect 24673 22661 24685 22695
rect 24719 22661 24731 22695
rect 24673 22655 24731 22661
rect 25130 22652 25136 22704
rect 25188 22692 25194 22704
rect 25501 22695 25559 22701
rect 25501 22692 25513 22695
rect 25188 22664 25513 22692
rect 25188 22652 25194 22664
rect 25501 22661 25513 22664
rect 25547 22661 25559 22695
rect 25501 22655 25559 22661
rect 26878 22652 26884 22704
rect 26936 22652 26942 22704
rect 27172 22701 27200 22732
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 28169 22763 28227 22769
rect 27488 22732 28028 22760
rect 27488 22720 27494 22732
rect 27157 22695 27215 22701
rect 27157 22661 27169 22695
rect 27203 22661 27215 22695
rect 27157 22655 27215 22661
rect 27341 22695 27399 22701
rect 27341 22661 27353 22695
rect 27387 22692 27399 22695
rect 27706 22692 27712 22704
rect 27387 22664 27712 22692
rect 27387 22661 27399 22664
rect 27341 22655 27399 22661
rect 27706 22652 27712 22664
rect 27764 22652 27770 22704
rect 27890 22652 27896 22704
rect 27948 22652 27954 22704
rect 23845 22627 23903 22633
rect 23845 22624 23857 22627
rect 23808 22596 23857 22624
rect 23808 22584 23814 22596
rect 23845 22593 23857 22596
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22593 24179 22627
rect 24121 22587 24179 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 23290 22556 23296 22568
rect 22848 22528 23296 22556
rect 22244 22448 22250 22460
rect 20855 22392 21594 22420
rect 20855 22389 20867 22392
rect 20809 22383 20867 22389
rect 21634 22380 21640 22432
rect 21692 22420 21698 22432
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21692 22392 21833 22420
rect 21692 22380 21698 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 22278 22380 22284 22432
rect 22336 22380 22342 22432
rect 22646 22380 22652 22432
rect 22704 22420 22710 22432
rect 22848 22420 22876 22528
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 24136 22556 24164 22587
rect 24394 22584 24400 22636
rect 24452 22584 24458 22636
rect 24486 22584 24492 22636
rect 24544 22624 24550 22636
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 24544 22596 24593 22624
rect 24544 22584 24550 22596
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 25777 22627 25835 22633
rect 25516 22596 25728 22624
rect 25516 22556 25544 22596
rect 23532 22528 24164 22556
rect 24780 22528 25544 22556
rect 25593 22559 25651 22565
rect 23532 22516 23538 22528
rect 23017 22491 23075 22497
rect 23017 22457 23029 22491
rect 23063 22488 23075 22491
rect 23566 22488 23572 22500
rect 23063 22460 23572 22488
rect 23063 22457 23075 22460
rect 23017 22451 23075 22457
rect 23566 22448 23572 22460
rect 23624 22448 23630 22500
rect 24780 22488 24808 22528
rect 25593 22525 25605 22559
rect 25639 22525 25651 22559
rect 25700 22556 25728 22596
rect 25777 22593 25789 22627
rect 25823 22624 25835 22627
rect 26234 22624 26240 22636
rect 25823 22596 26240 22624
rect 25823 22593 25835 22596
rect 25777 22587 25835 22593
rect 26234 22584 26240 22596
rect 26292 22624 26298 22636
rect 26896 22624 26924 22652
rect 26292 22596 26924 22624
rect 26292 22584 26298 22596
rect 27614 22584 27620 22636
rect 27672 22584 27678 22636
rect 28000 22633 28028 22732
rect 28169 22729 28181 22763
rect 28215 22729 28227 22763
rect 28169 22723 28227 22729
rect 28074 22652 28080 22704
rect 28132 22692 28138 22704
rect 28184 22692 28212 22723
rect 28534 22720 28540 22772
rect 28592 22720 28598 22772
rect 29089 22695 29147 22701
rect 29089 22692 29101 22695
rect 28132 22664 29101 22692
rect 28132 22652 28138 22664
rect 29089 22661 29101 22664
rect 29135 22661 29147 22695
rect 29089 22655 29147 22661
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 26602 22556 26608 22568
rect 25700 22528 26608 22556
rect 25593 22519 25651 22525
rect 25608 22488 25636 22519
rect 26602 22516 26608 22528
rect 26660 22516 26666 22568
rect 27816 22556 27844 22587
rect 28258 22584 28264 22636
rect 28316 22584 28322 22636
rect 28350 22584 28356 22636
rect 28408 22624 28414 22636
rect 28445 22627 28503 22633
rect 28445 22624 28457 22627
rect 28408 22596 28457 22624
rect 28408 22584 28414 22596
rect 28445 22593 28457 22596
rect 28491 22593 28503 22627
rect 28445 22587 28503 22593
rect 28626 22584 28632 22636
rect 28684 22584 28690 22636
rect 28905 22627 28963 22633
rect 28905 22593 28917 22627
rect 28951 22593 28963 22627
rect 28905 22587 28963 22593
rect 28644 22556 28672 22584
rect 27816 22528 28672 22556
rect 23676 22460 24808 22488
rect 24872 22460 25636 22488
rect 23676 22429 23704 22460
rect 24872 22432 24900 22460
rect 25866 22448 25872 22500
rect 25924 22448 25930 22500
rect 27982 22488 27988 22500
rect 27448 22460 27988 22488
rect 22704 22392 22876 22420
rect 23661 22423 23719 22429
rect 22704 22380 22710 22392
rect 23661 22389 23673 22423
rect 23707 22389 23719 22423
rect 23661 22383 23719 22389
rect 24854 22380 24860 22432
rect 24912 22380 24918 22432
rect 24946 22380 24952 22432
rect 25004 22380 25010 22432
rect 25774 22380 25780 22432
rect 25832 22380 25838 22432
rect 25884 22420 25912 22448
rect 27448 22432 27476 22460
rect 27982 22448 27988 22460
rect 28040 22488 28046 22500
rect 28920 22488 28948 22587
rect 28040 22460 28948 22488
rect 28040 22448 28046 22460
rect 26142 22420 26148 22432
rect 25884 22392 26148 22420
rect 26142 22380 26148 22392
rect 26200 22380 26206 22432
rect 27430 22380 27436 22432
rect 27488 22380 27494 22432
rect 27525 22423 27583 22429
rect 27525 22389 27537 22423
rect 27571 22420 27583 22423
rect 27614 22420 27620 22432
rect 27571 22392 27620 22420
rect 27571 22389 27583 22392
rect 27525 22383 27583 22389
rect 27614 22380 27620 22392
rect 27672 22380 27678 22432
rect 27890 22380 27896 22432
rect 27948 22420 27954 22432
rect 28442 22420 28448 22432
rect 27948 22392 28448 22420
rect 27948 22380 27954 22392
rect 28442 22380 28448 22392
rect 28500 22380 28506 22432
rect 28626 22380 28632 22432
rect 28684 22420 28690 22432
rect 29273 22423 29331 22429
rect 29273 22420 29285 22423
rect 28684 22392 29285 22420
rect 28684 22380 28690 22392
rect 29273 22389 29285 22392
rect 29319 22389 29331 22423
rect 29273 22383 29331 22389
rect 1104 22330 43884 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 43884 22330
rect 1104 22256 43884 22278
rect 2866 22176 2872 22228
rect 2924 22216 2930 22228
rect 3605 22219 3663 22225
rect 3605 22216 3617 22219
rect 2924 22188 3617 22216
rect 2924 22176 2930 22188
rect 3605 22185 3617 22188
rect 3651 22185 3663 22219
rect 4706 22216 4712 22228
rect 3605 22179 3663 22185
rect 3804 22188 4712 22216
rect 3694 22148 3700 22160
rect 3068 22120 3700 22148
rect 1210 22040 1216 22092
rect 1268 22080 1274 22092
rect 1857 22083 1915 22089
rect 1857 22080 1869 22083
rect 1268 22052 1869 22080
rect 1268 22040 1274 22052
rect 1857 22049 1869 22052
rect 1903 22049 1915 22083
rect 1857 22043 1915 22049
rect 1578 21972 1584 22024
rect 1636 21972 1642 22024
rect 3068 22021 3096 22120
rect 3694 22108 3700 22120
rect 3752 22108 3758 22160
rect 3418 22040 3424 22092
rect 3476 22040 3482 22092
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 21981 3111 22015
rect 3053 21975 3111 21981
rect 3436 21944 3464 22040
rect 3804 22021 3832 22188
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 5350 22176 5356 22228
rect 5408 22176 5414 22228
rect 5626 22176 5632 22228
rect 5684 22176 5690 22228
rect 7926 22216 7932 22228
rect 5736 22188 7932 22216
rect 4614 22108 4620 22160
rect 4672 22148 4678 22160
rect 5644 22148 5672 22176
rect 4672 22120 5672 22148
rect 4672 22108 4678 22120
rect 5736 22092 5764 22188
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 8110 22176 8116 22228
rect 8168 22216 8174 22228
rect 8389 22219 8447 22225
rect 8389 22216 8401 22219
rect 8168 22188 8401 22216
rect 8168 22176 8174 22188
rect 8389 22185 8401 22188
rect 8435 22185 8447 22219
rect 8389 22179 8447 22185
rect 9217 22219 9275 22225
rect 9217 22185 9229 22219
rect 9263 22216 9275 22219
rect 9398 22216 9404 22228
rect 9263 22188 9404 22216
rect 9263 22185 9275 22188
rect 9217 22179 9275 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 9824 22188 10241 22216
rect 9824 22176 9830 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 10229 22179 10287 22185
rect 11057 22219 11115 22225
rect 11057 22185 11069 22219
rect 11103 22216 11115 22219
rect 11146 22216 11152 22228
rect 11103 22188 11152 22216
rect 11103 22185 11115 22188
rect 11057 22179 11115 22185
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11514 22176 11520 22228
rect 11572 22216 11578 22228
rect 12342 22216 12348 22228
rect 11572 22188 12348 22216
rect 11572 22176 11578 22188
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 13906 22216 13912 22228
rect 13648 22188 13912 22216
rect 5902 22108 5908 22160
rect 5960 22148 5966 22160
rect 5997 22151 6055 22157
rect 5997 22148 6009 22151
rect 5960 22120 6009 22148
rect 5960 22108 5966 22120
rect 5997 22117 6009 22120
rect 6043 22117 6055 22151
rect 5997 22111 6055 22117
rect 6380 22120 6675 22148
rect 4157 22083 4215 22089
rect 4157 22049 4169 22083
rect 4203 22080 4215 22083
rect 4338 22080 4344 22092
rect 4203 22052 4344 22080
rect 4203 22049 4215 22052
rect 4157 22043 4215 22049
rect 4338 22040 4344 22052
rect 4396 22080 4402 22092
rect 5258 22080 5264 22092
rect 4396 22052 5264 22080
rect 4396 22040 4402 22052
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 5718 22080 5724 22092
rect 5644 22052 5724 22080
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3789 21975 3847 21981
rect 3896 21984 3985 22012
rect 3896 21944 3924 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4798 21972 4804 22024
rect 4856 21972 4862 22024
rect 5074 21972 5080 22024
rect 5132 21972 5138 22024
rect 5169 22015 5227 22021
rect 5169 21981 5181 22015
rect 5215 22012 5227 22015
rect 5350 22012 5356 22024
rect 5215 21984 5356 22012
rect 5215 21981 5227 21984
rect 5169 21975 5227 21981
rect 5350 21972 5356 21984
rect 5408 22012 5414 22024
rect 5644 22021 5672 22052
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 6270 22080 6276 22092
rect 5828 22052 6276 22080
rect 5828 22021 5856 22052
rect 6270 22040 6276 22052
rect 6328 22040 6334 22092
rect 5445 22015 5503 22021
rect 5445 22012 5457 22015
rect 5408 21984 5457 22012
rect 5408 21972 5414 21984
rect 5445 21981 5457 21984
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5813 22015 5871 22021
rect 5813 21981 5825 22015
rect 5859 21981 5871 22015
rect 5813 21975 5871 21981
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6086 21972 6092 22024
rect 6144 21972 6150 22024
rect 6182 22015 6240 22021
rect 6182 21981 6194 22015
rect 6228 21981 6240 22015
rect 6380 22012 6408 22120
rect 6454 22040 6460 22092
rect 6512 22080 6518 22092
rect 6647 22080 6675 22120
rect 6730 22108 6736 22160
rect 6788 22108 6794 22160
rect 7098 22108 7104 22160
rect 7156 22108 7162 22160
rect 8846 22108 8852 22160
rect 8904 22148 8910 22160
rect 8904 22120 9858 22148
rect 8904 22108 8910 22120
rect 7116 22080 7144 22108
rect 8018 22080 8024 22092
rect 6512 22052 6592 22080
rect 6647 22052 7144 22080
rect 7760 22052 8024 22080
rect 6512 22040 6518 22052
rect 6564 22021 6592 22052
rect 6564 22015 6631 22021
rect 6380 21984 6500 22012
rect 6564 21984 6585 22015
rect 6182 21975 6240 21981
rect 3436 21916 3924 21944
rect 4430 21904 4436 21956
rect 4488 21944 4494 21956
rect 4709 21947 4767 21953
rect 4709 21944 4721 21947
rect 4488 21916 4721 21944
rect 4488 21904 4494 21916
rect 4709 21913 4721 21916
rect 4755 21913 4767 21947
rect 4709 21907 4767 21913
rect 4982 21904 4988 21956
rect 5040 21904 5046 21956
rect 5258 21904 5264 21956
rect 5316 21944 5322 21956
rect 5721 21947 5779 21953
rect 5316 21916 5580 21944
rect 5316 21904 5322 21916
rect 3973 21879 4031 21885
rect 3973 21845 3985 21879
rect 4019 21876 4031 21879
rect 5442 21876 5448 21888
rect 4019 21848 5448 21876
rect 4019 21845 4031 21848
rect 3973 21839 4031 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 5552 21876 5580 21916
rect 5721 21913 5733 21947
rect 5767 21944 5779 21947
rect 6012 21944 6040 21972
rect 6197 21944 6225 21975
rect 6472 21953 6500 21984
rect 6573 21981 6585 21984
rect 6619 21981 6631 22015
rect 7374 22012 7380 22024
rect 6573 21975 6631 21981
rect 6749 21984 7380 22012
rect 5767 21916 5948 21944
rect 6012 21916 6225 21944
rect 6365 21947 6423 21953
rect 5767 21913 5779 21916
rect 5721 21907 5779 21913
rect 5810 21876 5816 21888
rect 5552 21848 5816 21876
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 5920 21876 5948 21916
rect 6365 21913 6377 21947
rect 6411 21913 6423 21947
rect 6365 21907 6423 21913
rect 6457 21947 6515 21953
rect 6457 21913 6469 21947
rect 6503 21913 6515 21947
rect 6457 21907 6515 21913
rect 6178 21876 6184 21888
rect 5920 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 6380 21876 6408 21907
rect 6749 21876 6777 21984
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 7760 22012 7788 22052
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 8352 22052 9076 22080
rect 8352 22040 8358 22052
rect 9048 22024 9076 22052
rect 9122 22040 9128 22092
rect 9180 22080 9186 22092
rect 9180 22052 9444 22080
rect 9180 22040 9186 22052
rect 9416 22024 9444 22052
rect 9490 22040 9496 22092
rect 9548 22080 9554 22092
rect 9548 22052 9628 22080
rect 9548 22040 9554 22052
rect 7489 21984 7788 22012
rect 7837 22015 7895 22021
rect 6822 21904 6828 21956
rect 6880 21904 6886 21956
rect 7098 21904 7104 21956
rect 7156 21944 7162 21956
rect 7489 21944 7517 21984
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 22012 8263 22015
rect 8386 22012 8392 22024
rect 8251 21984 8392 22012
rect 8251 21981 8263 21984
rect 8205 21975 8263 21981
rect 7156 21916 7517 21944
rect 7156 21904 7162 21916
rect 7558 21904 7564 21956
rect 7616 21904 7622 21956
rect 7852 21888 7880 21975
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 8478 21972 8484 22024
rect 8536 22012 8542 22024
rect 8573 22015 8631 22021
rect 8573 22012 8585 22015
rect 8536 21984 8585 22012
rect 8536 21972 8542 21984
rect 8573 21981 8585 21984
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 7926 21904 7932 21956
rect 7984 21944 7990 21956
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 7984 21916 8033 21944
rect 7984 21904 7990 21916
rect 8021 21913 8033 21916
rect 8067 21913 8079 21947
rect 8021 21907 8079 21913
rect 8110 21904 8116 21956
rect 8168 21904 8174 21956
rect 8588 21944 8616 21975
rect 8662 21972 8668 22024
rect 8720 22012 8726 22024
rect 8757 22015 8815 22021
rect 8757 22012 8769 22015
rect 8720 21984 8769 22012
rect 8720 21972 8726 21984
rect 8757 21981 8769 21984
rect 8803 21981 8815 22015
rect 8757 21975 8815 21981
rect 9030 21972 9036 22024
rect 9088 21972 9094 22024
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 9324 21944 9352 21975
rect 9398 21972 9404 22024
rect 9456 22012 9462 22024
rect 9600 22021 9628 22052
rect 9830 22021 9858 22120
rect 9950 22108 9956 22160
rect 10008 22108 10014 22160
rect 10962 22148 10968 22160
rect 10434 22120 10968 22148
rect 10434 22021 10462 22120
rect 10962 22108 10968 22120
rect 11020 22148 11026 22160
rect 11885 22151 11943 22157
rect 11020 22120 11836 22148
rect 11020 22108 11026 22120
rect 11808 22092 11836 22120
rect 11885 22117 11897 22151
rect 11931 22117 11943 22151
rect 11885 22111 11943 22117
rect 10594 22040 10600 22092
rect 10652 22040 10658 22092
rect 10873 22083 10931 22089
rect 10873 22049 10885 22083
rect 10919 22080 10931 22083
rect 11238 22080 11244 22092
rect 10919 22052 11244 22080
rect 10919 22049 10931 22052
rect 10873 22043 10931 22049
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 11790 22040 11796 22092
rect 11848 22040 11854 22092
rect 11900 22080 11928 22111
rect 11974 22108 11980 22160
rect 12032 22148 12038 22160
rect 12032 22120 12480 22148
rect 12032 22108 12038 22120
rect 11900 22052 12020 22080
rect 9585 22015 9643 22021
rect 9456 21984 9501 22012
rect 9456 21972 9462 21984
rect 9585 21981 9597 22015
rect 9631 21981 9643 22015
rect 9585 21975 9643 21981
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 9815 22015 9873 22021
rect 9815 21981 9827 22015
rect 9861 21981 9873 22015
rect 9815 21975 9873 21981
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 21981 10471 22015
rect 10413 21975 10471 21981
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 10612 22012 10640 22040
rect 10715 22015 10773 22021
rect 10715 22012 10727 22015
rect 10612 21984 10727 22012
rect 10505 21975 10563 21981
rect 10715 21981 10727 21984
rect 10761 21981 10773 22015
rect 10715 21975 10773 21981
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 21981 11023 22015
rect 10965 21975 11023 21981
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 22012 11207 22015
rect 11256 22012 11284 22040
rect 11195 21984 11284 22012
rect 11333 22015 11391 22021
rect 11195 21981 11207 21984
rect 11149 21975 11207 21981
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 11422 22012 11428 22024
rect 11379 21984 11428 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 9490 21944 9496 21956
rect 8588 21916 8984 21944
rect 9324 21916 9496 21944
rect 6380 21848 6777 21876
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7834 21876 7840 21888
rect 6972 21848 7840 21876
rect 6972 21836 6978 21848
rect 7834 21836 7840 21848
rect 7892 21876 7898 21888
rect 8202 21876 8208 21888
rect 7892 21848 8208 21876
rect 7892 21836 7898 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 8757 21879 8815 21885
rect 8757 21845 8769 21879
rect 8803 21876 8815 21879
rect 8846 21876 8852 21888
rect 8803 21848 8852 21876
rect 8803 21845 8815 21848
rect 8757 21839 8815 21845
rect 8846 21836 8852 21848
rect 8904 21836 8910 21888
rect 8956 21876 8984 21916
rect 9490 21904 9496 21916
rect 9548 21904 9554 21956
rect 9692 21888 9720 21975
rect 9398 21876 9404 21888
rect 8956 21848 9404 21876
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 9830 21876 9858 21975
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10530 21944 10558 21975
rect 10192 21916 10558 21944
rect 10192 21904 10198 21916
rect 10594 21904 10600 21956
rect 10652 21904 10658 21956
rect 10410 21876 10416 21888
rect 9830 21848 10416 21876
rect 10410 21836 10416 21848
rect 10468 21836 10474 21888
rect 10502 21836 10508 21888
rect 10560 21876 10566 21888
rect 10980 21876 11008 21975
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 11701 22015 11759 22021
rect 11701 21981 11713 22015
rect 11747 22012 11759 22015
rect 11882 22012 11888 22024
rect 11747 21984 11888 22012
rect 11747 21981 11759 21984
rect 11701 21975 11759 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 11992 22021 12020 22052
rect 12176 22021 12204 22120
rect 12342 22040 12348 22092
rect 12400 22040 12406 22092
rect 12452 22080 12480 22120
rect 13170 22108 13176 22160
rect 13228 22148 13234 22160
rect 13446 22148 13452 22160
rect 13228 22120 13452 22148
rect 13228 22108 13234 22120
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 12452 22052 13400 22080
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12125 22015 12204 22021
rect 12125 21981 12137 22015
rect 12171 21984 12204 22015
rect 12253 22015 12311 22021
rect 12171 21981 12183 21984
rect 12125 21975 12183 21981
rect 12253 21981 12265 22015
rect 12299 22012 12311 22015
rect 12360 22012 12388 22040
rect 13372 22024 13400 22052
rect 12299 21984 12388 22012
rect 12299 21981 12311 21984
rect 12253 21975 12311 21981
rect 12434 21972 12440 22024
rect 12492 22021 12498 22024
rect 12492 22015 12541 22021
rect 12492 21981 12495 22015
rect 12529 22012 12541 22015
rect 12529 21984 13032 22012
rect 12529 21981 12541 21984
rect 12492 21975 12541 21981
rect 12492 21972 12498 21975
rect 11514 21904 11520 21956
rect 11572 21904 11578 21956
rect 11609 21947 11667 21953
rect 11609 21913 11621 21947
rect 11655 21944 11667 21947
rect 11790 21944 11796 21956
rect 11655 21916 11796 21944
rect 11655 21913 11667 21916
rect 11609 21907 11667 21913
rect 11790 21904 11796 21916
rect 11848 21904 11854 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12268 21916 12357 21944
rect 12268 21888 12296 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 13004 21944 13032 21984
rect 13262 21972 13268 22024
rect 13320 21972 13326 22024
rect 13354 21972 13360 22024
rect 13412 22012 13418 22024
rect 13412 21984 13457 22012
rect 13412 21972 13418 21984
rect 13538 21972 13544 22024
rect 13596 21972 13602 22024
rect 13648 22021 13676 22188
rect 13906 22176 13912 22188
rect 13964 22176 13970 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 14642 22216 14648 22228
rect 14332 22188 14648 22216
rect 14332 22176 14338 22188
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 16482 22176 16488 22228
rect 16540 22176 16546 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 16853 22219 16911 22225
rect 16853 22216 16865 22219
rect 16632 22188 16865 22216
rect 16632 22176 16638 22188
rect 16853 22185 16865 22188
rect 16899 22185 16911 22219
rect 16853 22179 16911 22185
rect 16942 22176 16948 22228
rect 17000 22216 17006 22228
rect 17000 22188 18000 22216
rect 17000 22176 17006 22188
rect 13722 22108 13728 22160
rect 13780 22148 13786 22160
rect 13780 22120 13952 22148
rect 13780 22108 13786 22120
rect 13740 22021 13768 22108
rect 13924 22080 13952 22120
rect 15286 22108 15292 22160
rect 15344 22148 15350 22160
rect 16500 22148 16528 22176
rect 17310 22148 17316 22160
rect 15344 22120 16436 22148
rect 16500 22120 17316 22148
rect 15344 22108 15350 22120
rect 15565 22083 15623 22089
rect 15565 22080 15577 22083
rect 13924 22052 15577 22080
rect 15565 22049 15577 22052
rect 15611 22049 15623 22083
rect 16298 22080 16304 22092
rect 15565 22043 15623 22049
rect 16040 22052 16304 22080
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 21981 13691 22015
rect 13633 21975 13691 21981
rect 13730 22015 13788 22021
rect 13730 21981 13742 22015
rect 13776 21981 13788 22015
rect 13730 21975 13788 21981
rect 13740 21944 13768 21975
rect 14090 21972 14096 22024
rect 14148 21972 14154 22024
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 14918 22012 14924 22024
rect 14700 21984 14924 22012
rect 14700 21972 14706 21984
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15010 21972 15016 22024
rect 15068 22012 15074 22024
rect 16040 22021 16068 22052
rect 16298 22040 16304 22052
rect 16356 22040 16362 22092
rect 16408 22080 16436 22120
rect 17310 22108 17316 22120
rect 17368 22108 17374 22160
rect 17972 22148 18000 22188
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18601 22219 18659 22225
rect 18601 22216 18613 22219
rect 18288 22188 18613 22216
rect 18288 22176 18294 22188
rect 18601 22185 18613 22188
rect 18647 22185 18659 22219
rect 18601 22179 18659 22185
rect 19429 22219 19487 22225
rect 19429 22185 19441 22219
rect 19475 22185 19487 22219
rect 19429 22179 19487 22185
rect 18509 22151 18567 22157
rect 18509 22148 18521 22151
rect 17420 22120 17908 22148
rect 17972 22120 18521 22148
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16408 22052 16957 22080
rect 16592 22024 16620 22052
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17420 22024 17448 22120
rect 17678 22040 17684 22092
rect 17736 22040 17742 22092
rect 17880 22089 17908 22120
rect 18509 22117 18521 22120
rect 18555 22117 18567 22151
rect 19061 22151 19119 22157
rect 19061 22148 19073 22151
rect 18509 22111 18567 22117
rect 18616 22120 19073 22148
rect 17865 22083 17923 22089
rect 17865 22049 17877 22083
rect 17911 22049 17923 22083
rect 17865 22043 17923 22049
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 15068 21984 15117 22012
rect 15068 21972 15074 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15105 21975 15163 21981
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 21981 15439 22015
rect 15381 21975 15439 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 14108 21944 14136 21972
rect 13004 21916 13768 21944
rect 13832 21916 14136 21944
rect 12345 21907 12403 21913
rect 10560 21848 11008 21876
rect 10560 21836 10566 21848
rect 12250 21836 12256 21888
rect 12308 21836 12314 21888
rect 12618 21836 12624 21888
rect 12676 21836 12682 21888
rect 13173 21879 13231 21885
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13832 21876 13860 21916
rect 13219 21848 13860 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13906 21836 13912 21888
rect 13964 21836 13970 21888
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14550 21876 14556 21888
rect 14056 21848 14556 21876
rect 14056 21836 14062 21848
rect 14550 21836 14556 21848
rect 14608 21836 14614 21888
rect 15212 21876 15240 21975
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 15396 21944 15424 21975
rect 16574 21972 16580 22024
rect 16632 21972 16638 22024
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 21981 17187 22015
rect 17129 21975 17187 21981
rect 16485 21947 16543 21953
rect 15344 21916 16436 21944
rect 15344 21904 15350 21916
rect 16408 21888 16436 21916
rect 16485 21913 16497 21947
rect 16531 21913 16543 21947
rect 16485 21907 16543 21913
rect 16853 21947 16911 21953
rect 16853 21913 16865 21947
rect 16899 21944 16911 21947
rect 16942 21944 16948 21956
rect 16899 21916 16948 21944
rect 16899 21913 16911 21916
rect 16853 21907 16911 21913
rect 15746 21876 15752 21888
rect 15212 21848 15752 21876
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 16209 21879 16267 21885
rect 16209 21876 16221 21879
rect 15988 21848 16221 21876
rect 15988 21836 15994 21848
rect 16209 21845 16221 21848
rect 16255 21845 16267 21879
rect 16209 21839 16267 21845
rect 16390 21836 16396 21888
rect 16448 21836 16454 21888
rect 16500 21876 16528 21907
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17144 21944 17172 21975
rect 17402 21972 17408 22024
rect 17460 21972 17466 22024
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 22012 17831 22015
rect 18414 22012 18420 22024
rect 17819 21984 18420 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18616 22012 18644 22120
rect 19061 22117 19073 22120
rect 19107 22117 19119 22151
rect 19444 22148 19472 22179
rect 19518 22176 19524 22228
rect 19576 22216 19582 22228
rect 19797 22219 19855 22225
rect 19797 22216 19809 22219
rect 19576 22188 19809 22216
rect 19576 22176 19582 22188
rect 19797 22185 19809 22188
rect 19843 22185 19855 22219
rect 19797 22179 19855 22185
rect 19978 22176 19984 22228
rect 20036 22176 20042 22228
rect 20257 22219 20315 22225
rect 20257 22185 20269 22219
rect 20303 22216 20315 22219
rect 20303 22188 20944 22216
rect 20303 22185 20315 22188
rect 20257 22179 20315 22185
rect 19996 22148 20024 22176
rect 20438 22148 20444 22160
rect 19444 22120 20024 22148
rect 20088 22120 20444 22148
rect 19061 22111 19119 22117
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 19334 22080 19340 22092
rect 18831 22052 19340 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19426 22040 19432 22092
rect 19484 22040 19490 22092
rect 19521 22083 19579 22089
rect 19521 22049 19533 22083
rect 19567 22080 19579 22083
rect 19794 22080 19800 22092
rect 19567 22052 19800 22080
rect 19567 22049 19579 22052
rect 19521 22043 19579 22049
rect 19794 22040 19800 22052
rect 19852 22040 19858 22092
rect 18524 21984 18644 22012
rect 17494 21944 17500 21956
rect 17144 21916 17500 21944
rect 17494 21904 17500 21916
rect 17552 21944 17558 21956
rect 17678 21944 17684 21956
rect 17552 21916 17684 21944
rect 17552 21904 17558 21916
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 18524 21944 18552 21984
rect 18874 21972 18880 22024
rect 18932 21972 18938 22024
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19116 21984 19257 22012
rect 19116 21972 19122 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19444 22012 19472 22040
rect 20088 22012 20116 22120
rect 20438 22108 20444 22120
rect 20496 22108 20502 22160
rect 20806 22108 20812 22160
rect 20864 22108 20870 22160
rect 20916 22148 20944 22188
rect 20990 22176 20996 22228
rect 21048 22216 21054 22228
rect 21085 22219 21143 22225
rect 21085 22216 21097 22219
rect 21048 22188 21097 22216
rect 21048 22176 21054 22188
rect 21085 22185 21097 22188
rect 21131 22216 21143 22219
rect 21634 22216 21640 22228
rect 21131 22188 21640 22216
rect 21131 22185 21143 22188
rect 21085 22179 21143 22185
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 24210 22176 24216 22228
rect 24268 22176 24274 22228
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 25777 22219 25835 22225
rect 24452 22188 25544 22216
rect 24452 22176 24458 22188
rect 21358 22148 21364 22160
rect 20916 22120 21364 22148
rect 21358 22108 21364 22120
rect 21416 22148 21422 22160
rect 24228 22148 24256 22176
rect 24578 22148 24584 22160
rect 21416 22120 24190 22148
rect 24228 22120 24584 22148
rect 21416 22108 21422 22120
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22080 20223 22083
rect 20714 22080 20720 22092
rect 20211 22052 20720 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 19444 21984 20116 22012
rect 19245 21975 19303 21981
rect 17788 21916 18552 21944
rect 18601 21947 18659 21953
rect 17788 21876 17816 21916
rect 18601 21913 18613 21947
rect 18647 21944 18659 21947
rect 19150 21944 19156 21956
rect 18647 21916 19156 21944
rect 18647 21913 18659 21916
rect 18601 21907 18659 21913
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 19981 21947 20039 21953
rect 19981 21913 19993 21947
rect 20027 21913 20039 21947
rect 20088 21944 20116 21984
rect 20254 21972 20260 22024
rect 20312 21972 20318 22024
rect 20824 22021 20852 22108
rect 20993 22083 21051 22089
rect 20993 22049 21005 22083
rect 21039 22080 21051 22083
rect 21174 22080 21180 22092
rect 21039 22052 21180 22080
rect 21039 22049 21051 22052
rect 20993 22043 21051 22049
rect 20625 22015 20683 22021
rect 20625 21981 20637 22015
rect 20671 21981 20683 22015
rect 20625 21975 20683 21981
rect 20803 22015 20861 22021
rect 20803 21981 20815 22015
rect 20849 21981 20861 22015
rect 20803 21975 20861 21981
rect 20640 21944 20668 21975
rect 20898 21972 20904 22024
rect 20956 21972 20962 22024
rect 20088 21916 20668 21944
rect 20717 21947 20775 21953
rect 19981 21907 20039 21913
rect 20717 21913 20729 21947
rect 20763 21944 20775 21947
rect 21008 21944 21036 22043
rect 21174 22040 21180 22052
rect 21232 22040 21238 22092
rect 21453 22083 21511 22089
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21726 22080 21732 22092
rect 21499 22052 21732 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 21726 22040 21732 22052
rect 21784 22080 21790 22092
rect 22186 22080 22192 22092
rect 21784 22052 22192 22080
rect 21784 22040 21790 22052
rect 22186 22040 22192 22052
rect 22244 22040 22250 22092
rect 23750 22080 23756 22092
rect 22480 22052 23244 22080
rect 21266 21972 21272 22024
rect 21324 22012 21330 22024
rect 21361 22015 21419 22021
rect 21361 22012 21373 22015
rect 21324 21984 21373 22012
rect 21324 21972 21330 21984
rect 21361 21981 21373 21984
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21542 21972 21548 22024
rect 21600 21972 21606 22024
rect 22480 22012 22508 22052
rect 21652 21984 22508 22012
rect 20763 21916 21036 21944
rect 20763 21913 20775 21916
rect 20717 21907 20775 21913
rect 16500 21848 17816 21876
rect 18046 21836 18052 21888
rect 18104 21876 18110 21888
rect 19610 21876 19616 21888
rect 18104 21848 19616 21876
rect 18104 21836 18110 21848
rect 19610 21836 19616 21848
rect 19668 21876 19674 21888
rect 19996 21876 20024 21907
rect 21082 21904 21088 21956
rect 21140 21944 21146 21956
rect 21652 21944 21680 21984
rect 22554 21972 22560 22024
rect 22612 21972 22618 22024
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 22012 22707 22015
rect 22738 22012 22744 22024
rect 22695 21984 22744 22012
rect 22695 21981 22707 21984
rect 22649 21975 22707 21981
rect 22738 21972 22744 21984
rect 22796 22012 22802 22024
rect 23106 22012 23112 22024
rect 22796 21984 23112 22012
rect 22796 21972 22802 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23216 22021 23244 22052
rect 23400 22052 23756 22080
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 21140 21916 21680 21944
rect 22572 21944 22600 21972
rect 23400 21956 23428 22052
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 24162 22080 24190 22120
rect 24578 22108 24584 22120
rect 24636 22108 24642 22160
rect 24670 22108 24676 22160
rect 24728 22148 24734 22160
rect 24728 22120 25269 22148
rect 24728 22108 24734 22120
rect 24162 22052 24624 22080
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 22012 23627 22015
rect 23658 22012 23664 22024
rect 23615 21984 23664 22012
rect 23615 21981 23627 21984
rect 23569 21975 23627 21981
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 22925 21947 22983 21953
rect 22925 21944 22937 21947
rect 22572 21916 22937 21944
rect 21140 21904 21146 21916
rect 22925 21913 22937 21916
rect 22971 21944 22983 21947
rect 23382 21944 23388 21956
rect 22971 21916 23388 21944
rect 22971 21913 22983 21916
rect 22925 21907 22983 21913
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21913 23535 21947
rect 23768 21944 23796 22040
rect 23842 21972 23848 22024
rect 23900 22012 23906 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23900 21984 24409 22012
rect 23900 21972 23906 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24490 22015 24548 22021
rect 24490 21981 24502 22015
rect 24536 21981 24548 22015
rect 24596 22012 24624 22052
rect 24762 22012 24768 22024
rect 24596 21984 24768 22012
rect 24490 21975 24548 21981
rect 23768 21916 23981 21944
rect 23477 21907 23535 21913
rect 19668 21848 20024 21876
rect 19668 21836 19674 21848
rect 20438 21836 20444 21888
rect 20496 21836 20502 21888
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 21269 21879 21327 21885
rect 21269 21876 21281 21879
rect 21232 21848 21281 21876
rect 21232 21836 21238 21848
rect 21269 21845 21281 21848
rect 21315 21845 21327 21879
rect 21269 21839 21327 21845
rect 21634 21836 21640 21888
rect 21692 21876 21698 21888
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 21692 21848 21833 21876
rect 21692 21836 21698 21848
rect 21821 21845 21833 21848
rect 21867 21845 21879 21879
rect 21821 21839 21879 21845
rect 22554 21836 22560 21888
rect 22612 21836 22618 21888
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 23492 21876 23520 21907
rect 23348 21848 23520 21876
rect 23348 21836 23354 21848
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 23753 21879 23811 21885
rect 23753 21876 23765 21879
rect 23716 21848 23765 21876
rect 23716 21836 23722 21848
rect 23753 21845 23765 21848
rect 23799 21845 23811 21879
rect 23953 21876 23981 21916
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24505 21944 24533 21975
rect 24762 21972 24768 21984
rect 24820 21972 24826 22024
rect 24862 22015 24920 22021
rect 24862 21981 24874 22015
rect 24908 21981 24920 22015
rect 24862 21975 24920 21981
rect 24084 21916 24533 21944
rect 24084 21904 24090 21916
rect 24670 21904 24676 21956
rect 24728 21904 24734 21956
rect 24877 21944 24905 21975
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25241 22021 25269 22120
rect 25516 22021 25544 22188
rect 25777 22185 25789 22219
rect 25823 22216 25835 22219
rect 25823 22188 25912 22216
rect 25823 22185 25835 22188
rect 25777 22179 25835 22185
rect 25590 22108 25596 22160
rect 25648 22108 25654 22160
rect 25884 22148 25912 22188
rect 26694 22176 26700 22228
rect 26752 22176 26758 22228
rect 27433 22219 27491 22225
rect 27433 22185 27445 22219
rect 27479 22216 27491 22219
rect 27890 22216 27896 22228
rect 27479 22188 27896 22216
rect 27479 22185 27491 22188
rect 27433 22179 27491 22185
rect 27890 22176 27896 22188
rect 27948 22176 27954 22228
rect 27985 22219 28043 22225
rect 27985 22185 27997 22219
rect 28031 22216 28043 22219
rect 28074 22216 28080 22228
rect 28031 22188 28080 22216
rect 28031 22185 28043 22188
rect 27985 22179 28043 22185
rect 28074 22176 28080 22188
rect 28132 22176 28138 22228
rect 28721 22219 28779 22225
rect 28721 22185 28733 22219
rect 28767 22185 28779 22219
rect 28721 22179 28779 22185
rect 26050 22148 26056 22160
rect 25884 22120 26056 22148
rect 26050 22108 26056 22120
rect 26108 22148 26114 22160
rect 28736 22148 28764 22179
rect 26108 22120 26740 22148
rect 26108 22108 26114 22120
rect 25608 22080 25636 22108
rect 25608 22052 26005 22080
rect 25226 22015 25284 22021
rect 25226 21981 25238 22015
rect 25272 21981 25284 22015
rect 25226 21975 25284 21981
rect 25501 22015 25559 22021
rect 25501 21981 25513 22015
rect 25547 21981 25559 22015
rect 25501 21975 25559 21981
rect 25590 21972 25596 22024
rect 25648 22021 25654 22024
rect 25648 22012 25656 22021
rect 25648 21984 25693 22012
rect 25648 21975 25656 21984
rect 25648 21972 25654 21975
rect 25774 21972 25780 22024
rect 25832 22012 25838 22024
rect 25977 22021 26005 22052
rect 26142 22040 26148 22092
rect 26200 22080 26206 22092
rect 26712 22089 26740 22120
rect 27264 22120 27844 22148
rect 26697 22083 26755 22089
rect 26200 22052 26280 22080
rect 26200 22040 26206 22052
rect 26252 22021 26280 22052
rect 26697 22049 26709 22083
rect 26743 22049 26755 22083
rect 27264 22080 27292 22120
rect 26697 22043 26755 22049
rect 26896 22052 27292 22080
rect 27341 22083 27399 22089
rect 25869 22015 25927 22021
rect 25869 22012 25881 22015
rect 25832 21984 25881 22012
rect 25832 21972 25838 21984
rect 25869 21981 25881 21984
rect 25915 21981 25927 22015
rect 25869 21975 25927 21981
rect 25962 22015 26020 22021
rect 25962 21981 25974 22015
rect 26008 21981 26020 22015
rect 25962 21975 26020 21981
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 26326 21972 26332 22024
rect 26384 22021 26390 22024
rect 26384 22012 26392 22021
rect 26384 21984 26429 22012
rect 26384 21975 26392 21984
rect 26384 21972 26390 21975
rect 26602 21972 26608 22024
rect 26660 21972 26666 22024
rect 26786 21972 26792 22024
rect 26844 22012 26850 22024
rect 26896 22021 26924 22052
rect 27341 22049 27353 22083
rect 27387 22080 27399 22083
rect 27430 22080 27436 22092
rect 27387 22052 27436 22080
rect 27387 22049 27399 22052
rect 27341 22043 27399 22049
rect 27430 22040 27436 22052
rect 27488 22040 27494 22092
rect 27816 22089 27844 22120
rect 28092 22120 28764 22148
rect 28092 22092 28120 22120
rect 27801 22083 27859 22089
rect 27801 22049 27813 22083
rect 27847 22049 27859 22083
rect 27801 22043 27859 22049
rect 28074 22040 28080 22092
rect 28132 22040 28138 22092
rect 26881 22015 26939 22021
rect 26881 22012 26893 22015
rect 26844 21984 26893 22012
rect 26844 21972 26850 21984
rect 26881 21981 26893 21984
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 26970 21972 26976 22024
rect 27028 22012 27034 22024
rect 27249 22015 27307 22021
rect 27249 22012 27261 22015
rect 27028 21984 27261 22012
rect 27028 21972 27034 21984
rect 27249 21981 27261 21984
rect 27295 21981 27307 22015
rect 27249 21975 27307 21981
rect 27706 21972 27712 22024
rect 27764 21972 27770 22024
rect 27985 22015 28043 22021
rect 27985 21981 27997 22015
rect 28031 22012 28043 22015
rect 28092 22012 28120 22040
rect 28031 21984 28120 22012
rect 28261 22015 28319 22021
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 28261 21981 28273 22015
rect 28307 22012 28319 22015
rect 28350 22012 28356 22024
rect 28307 21984 28356 22012
rect 28307 21981 28319 21984
rect 28261 21975 28319 21981
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 28445 22015 28503 22021
rect 28445 21981 28457 22015
rect 28491 21981 28503 22015
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 28445 21975 28503 21981
rect 28552 21984 28733 22012
rect 24780 21916 24905 21944
rect 25409 21947 25467 21953
rect 24780 21888 24808 21916
rect 25409 21913 25421 21947
rect 25455 21944 25467 21947
rect 26142 21944 26148 21956
rect 25455 21916 26148 21944
rect 25455 21913 25467 21916
rect 25409 21907 25467 21913
rect 26142 21904 26148 21916
rect 26200 21904 26206 21956
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 28460 21944 28488 21975
rect 28552 21956 28580 21984
rect 28721 21981 28733 21984
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 28810 21972 28816 22024
rect 28868 21972 28874 22024
rect 27396 21916 28488 21944
rect 27396 21904 27402 21916
rect 28534 21904 28540 21956
rect 28592 21904 28598 21956
rect 24486 21876 24492 21888
rect 23953 21848 24492 21876
rect 23753 21839 23811 21845
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24762 21836 24768 21888
rect 24820 21836 24826 21888
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25866 21876 25872 21888
rect 25087 21848 25872 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 26513 21879 26571 21885
rect 26513 21845 26525 21879
rect 26559 21876 26571 21879
rect 26878 21876 26884 21888
rect 26559 21848 26884 21876
rect 26559 21845 26571 21848
rect 26513 21839 26571 21845
rect 26878 21836 26884 21848
rect 26936 21836 26942 21888
rect 27062 21836 27068 21888
rect 27120 21836 27126 21888
rect 27614 21836 27620 21888
rect 27672 21836 27678 21888
rect 27982 21836 27988 21888
rect 28040 21876 28046 21888
rect 28169 21879 28227 21885
rect 28169 21876 28181 21879
rect 28040 21848 28181 21876
rect 28040 21836 28046 21848
rect 28169 21845 28181 21848
rect 28215 21845 28227 21879
rect 28169 21839 28227 21845
rect 28258 21836 28264 21888
rect 28316 21876 28322 21888
rect 28442 21876 28448 21888
rect 28316 21848 28448 21876
rect 28316 21836 28322 21848
rect 28442 21836 28448 21848
rect 28500 21876 28506 21888
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 28500 21848 28641 21876
rect 28500 21836 28506 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 29086 21836 29092 21888
rect 29144 21836 29150 21888
rect 1104 21786 43884 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 43884 21786
rect 1104 21712 43884 21734
rect 1489 21675 1547 21681
rect 1489 21641 1501 21675
rect 1535 21672 1547 21675
rect 2866 21672 2872 21684
rect 1535 21644 2544 21672
rect 1535 21641 1547 21644
rect 1489 21635 1547 21641
rect 1946 21564 1952 21616
rect 2004 21564 2010 21616
rect 2406 21564 2412 21616
rect 2464 21564 2470 21616
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2424 21536 2452 21564
rect 1903 21508 2452 21536
rect 2516 21536 2544 21644
rect 2746 21644 2872 21672
rect 2584 21607 2642 21613
rect 2584 21573 2596 21607
rect 2630 21604 2642 21607
rect 2746 21604 2774 21644
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 3694 21632 3700 21684
rect 3752 21672 3758 21684
rect 3789 21675 3847 21681
rect 3789 21672 3801 21675
rect 3752 21644 3801 21672
rect 3752 21632 3758 21644
rect 3789 21641 3801 21644
rect 3835 21641 3847 21675
rect 3789 21635 3847 21641
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 4488 21644 5111 21672
rect 4488 21632 4494 21644
rect 2630 21576 2774 21604
rect 3896 21576 4752 21604
rect 2630 21573 2642 21576
rect 2584 21567 2642 21573
rect 3896 21536 3924 21576
rect 2516 21508 3924 21536
rect 3973 21539 4031 21545
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 3973 21505 3985 21539
rect 4019 21505 4031 21539
rect 3973 21499 4031 21505
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 2130 21428 2136 21480
rect 2188 21428 2194 21480
rect 2317 21471 2375 21477
rect 2317 21437 2329 21471
rect 2363 21437 2375 21471
rect 2317 21431 2375 21437
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2332 21332 2360 21431
rect 3510 21428 3516 21480
rect 3568 21468 3574 21480
rect 3878 21468 3884 21480
rect 3568 21440 3884 21468
rect 3568 21428 3574 21440
rect 3878 21428 3884 21440
rect 3936 21468 3942 21480
rect 3988 21468 4016 21499
rect 3936 21440 4016 21468
rect 4080 21468 4108 21499
rect 4154 21496 4160 21548
rect 4212 21496 4218 21548
rect 4246 21496 4252 21548
rect 4304 21545 4310 21548
rect 4304 21539 4333 21545
rect 4321 21505 4333 21539
rect 4304 21499 4333 21505
rect 4304 21496 4310 21499
rect 4430 21496 4436 21548
rect 4488 21496 4494 21548
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 4724 21545 4752 21576
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21505 4767 21539
rect 4709 21499 4767 21505
rect 4982 21496 4988 21548
rect 5040 21496 5046 21548
rect 5083 21545 5111 21644
rect 5442 21632 5448 21684
rect 5500 21632 5506 21684
rect 5626 21632 5632 21684
rect 5684 21632 5690 21684
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 5813 21675 5871 21681
rect 5813 21672 5825 21675
rect 5776 21644 5825 21672
rect 5776 21632 5782 21644
rect 5813 21641 5825 21644
rect 5859 21641 5871 21675
rect 5813 21635 5871 21641
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 5994 21672 6000 21684
rect 5951 21644 6000 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 8018 21672 8024 21684
rect 7760 21644 8024 21672
rect 5258 21564 5264 21616
rect 5316 21564 5322 21616
rect 5460 21604 5488 21632
rect 5460 21576 5780 21604
rect 5078 21539 5136 21545
rect 5078 21505 5090 21539
rect 5124 21505 5136 21539
rect 5078 21499 5136 21505
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 5752 21545 5780 21576
rect 6270 21564 6276 21616
rect 6328 21604 6334 21616
rect 7193 21607 7251 21613
rect 7193 21604 7205 21607
rect 6328 21576 7205 21604
rect 6328 21564 6334 21576
rect 7193 21573 7205 21576
rect 7239 21573 7251 21607
rect 7193 21567 7251 21573
rect 7282 21564 7288 21616
rect 7340 21604 7346 21616
rect 7760 21613 7788 21644
rect 8018 21632 8024 21644
rect 8076 21672 8082 21684
rect 8076 21644 8432 21672
rect 8076 21632 8082 21644
rect 7745 21607 7803 21613
rect 7340 21576 7604 21604
rect 7340 21564 7346 21576
rect 5450 21539 5508 21545
rect 5450 21505 5462 21539
rect 5496 21536 5508 21539
rect 5721 21539 5780 21545
rect 5496 21526 5580 21536
rect 5496 21508 5673 21526
rect 5496 21505 5508 21508
rect 5450 21499 5508 21505
rect 5552 21498 5673 21508
rect 5721 21505 5733 21539
rect 5767 21508 5780 21539
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 5645 21468 5673 21498
rect 5810 21496 5816 21548
rect 5868 21536 5874 21548
rect 6457 21539 6515 21545
rect 5868 21508 6224 21536
rect 5868 21496 5874 21508
rect 4080 21440 4660 21468
rect 5645 21440 5948 21468
rect 3936 21428 3942 21440
rect 3697 21403 3755 21409
rect 3697 21369 3709 21403
rect 3743 21400 3755 21403
rect 4338 21400 4344 21412
rect 3743 21372 4344 21400
rect 3743 21369 3755 21372
rect 3697 21363 3755 21369
rect 4338 21360 4344 21372
rect 4396 21360 4402 21412
rect 4522 21360 4528 21412
rect 4580 21360 4586 21412
rect 4632 21400 4660 21440
rect 5813 21403 5871 21409
rect 5813 21400 5825 21403
rect 4632 21372 5825 21400
rect 5813 21369 5825 21372
rect 5859 21369 5871 21403
rect 5920 21400 5948 21440
rect 6086 21428 6092 21480
rect 6144 21428 6150 21480
rect 6196 21468 6224 21508
rect 6457 21505 6469 21539
rect 6503 21536 6515 21539
rect 6822 21536 6828 21548
rect 6503 21508 6828 21536
rect 6503 21505 6515 21508
rect 6457 21499 6515 21505
rect 6822 21496 6828 21508
rect 6880 21536 6886 21548
rect 7374 21536 7380 21548
rect 6880 21508 7380 21536
rect 6880 21496 6886 21508
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7576 21536 7604 21576
rect 7745 21573 7757 21607
rect 7791 21573 7803 21607
rect 8294 21604 8300 21616
rect 7745 21567 7803 21573
rect 7963 21576 8300 21604
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7576 21508 7665 21536
rect 7469 21499 7527 21505
rect 7653 21505 7665 21508
rect 7699 21536 7711 21539
rect 7699 21508 7788 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 7006 21468 7012 21480
rect 6196 21440 7012 21468
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 6362 21400 6368 21412
rect 5920 21372 6368 21400
rect 5813 21363 5871 21369
rect 6362 21360 6368 21372
rect 6420 21400 6426 21412
rect 7190 21400 7196 21412
rect 6420 21372 7196 21400
rect 6420 21360 6426 21372
rect 7190 21360 7196 21372
rect 7248 21360 7254 21412
rect 7484 21400 7512 21499
rect 7650 21400 7656 21412
rect 7484 21372 7656 21400
rect 7650 21360 7656 21372
rect 7708 21360 7714 21412
rect 7760 21400 7788 21508
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 7963 21400 7991 21576
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 8404 21613 8432 21644
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 9214 21672 9220 21684
rect 8904 21644 9220 21672
rect 8904 21632 8910 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 9490 21632 9496 21684
rect 9548 21632 9554 21684
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 10873 21675 10931 21681
rect 10873 21672 10885 21675
rect 10652 21644 10885 21672
rect 10652 21632 10658 21644
rect 10873 21641 10885 21644
rect 10919 21641 10931 21675
rect 10873 21635 10931 21641
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11333 21675 11391 21681
rect 11333 21641 11345 21675
rect 11379 21672 11391 21675
rect 11422 21672 11428 21684
rect 11379 21644 11428 21672
rect 11379 21641 11391 21644
rect 11333 21635 11391 21641
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 11572 21644 11827 21672
rect 11572 21632 11578 21644
rect 8389 21607 8447 21613
rect 8389 21573 8401 21607
rect 8435 21604 8447 21607
rect 10042 21604 10048 21616
rect 8435 21576 10048 21604
rect 8435 21573 8447 21576
rect 8389 21567 8447 21573
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 10137 21607 10195 21613
rect 10137 21573 10149 21607
rect 10183 21604 10195 21607
rect 10505 21607 10563 21613
rect 10505 21604 10517 21607
rect 10183 21576 10517 21604
rect 10183 21573 10195 21576
rect 10137 21567 10195 21573
rect 10505 21573 10517 21576
rect 10551 21604 10563 21607
rect 10778 21604 10784 21616
rect 10551 21576 10784 21604
rect 10551 21573 10563 21576
rect 10505 21567 10563 21573
rect 10778 21564 10784 21576
rect 10836 21604 10842 21616
rect 11701 21607 11759 21613
rect 11701 21604 11713 21607
rect 10836 21576 11713 21604
rect 10836 21564 10842 21576
rect 11701 21573 11713 21576
rect 11747 21573 11759 21607
rect 11799 21604 11827 21644
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 13078 21672 13084 21684
rect 11940 21644 13084 21672
rect 11940 21632 11946 21644
rect 13078 21632 13084 21644
rect 13136 21632 13142 21684
rect 13262 21632 13268 21684
rect 13320 21632 13326 21684
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 14553 21675 14611 21681
rect 13412 21644 13865 21672
rect 13412 21632 13418 21644
rect 12802 21604 12808 21616
rect 11799 21576 12808 21604
rect 11701 21567 11759 21573
rect 12802 21564 12808 21576
rect 12860 21604 12866 21616
rect 12897 21607 12955 21613
rect 12897 21604 12909 21607
rect 12860 21576 12909 21604
rect 12860 21564 12866 21576
rect 12897 21573 12909 21576
rect 12943 21573 12955 21607
rect 12897 21567 12955 21573
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21536 8171 21539
rect 8202 21536 8208 21548
rect 8159 21508 8208 21536
rect 8159 21505 8171 21508
rect 8113 21499 8171 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21536 8539 21539
rect 8662 21536 8668 21548
rect 8527 21508 8668 21536
rect 8527 21505 8539 21508
rect 8481 21499 8539 21505
rect 8662 21496 8668 21508
rect 8720 21536 8726 21548
rect 8941 21539 8999 21545
rect 8941 21536 8953 21539
rect 8720 21508 8953 21536
rect 8720 21496 8726 21508
rect 8941 21505 8953 21508
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21505 9183 21539
rect 9125 21499 9183 21505
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 9140 21468 9168 21499
rect 8904 21440 9168 21468
rect 8904 21428 8910 21440
rect 7760 21372 7991 21400
rect 8386 21360 8392 21412
rect 8444 21400 8450 21412
rect 8864 21400 8892 21428
rect 8444 21372 8892 21400
rect 8444 21360 8450 21372
rect 8938 21360 8944 21412
rect 8996 21400 9002 21412
rect 9232 21400 9260 21499
rect 9306 21496 9312 21548
rect 9364 21545 9370 21548
rect 9364 21539 9413 21545
rect 9364 21505 9367 21539
rect 9401 21536 9413 21539
rect 9401 21508 9536 21536
rect 9401 21505 9413 21508
rect 9364 21499 9413 21505
rect 9364 21496 9370 21499
rect 9508 21480 9536 21508
rect 10870 21496 10876 21548
rect 10928 21536 10934 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10928 21508 10977 21536
rect 10928 21496 10934 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 11054 21496 11060 21548
rect 11112 21496 11118 21548
rect 11882 21536 11888 21548
rect 11164 21508 11888 21536
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 11164 21468 11192 21508
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 13096 21545 13124 21632
rect 13630 21564 13636 21616
rect 13688 21564 13694 21616
rect 13837 21604 13865 21644
rect 14553 21641 14565 21675
rect 14599 21672 14611 21675
rect 14826 21672 14832 21684
rect 14599 21644 14832 21672
rect 14599 21641 14611 21644
rect 14553 21635 14611 21641
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15470 21632 15476 21684
rect 15528 21632 15534 21684
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 15930 21672 15936 21684
rect 15620 21644 15936 21672
rect 15620 21632 15626 21644
rect 15930 21632 15936 21644
rect 15988 21632 15994 21684
rect 16298 21632 16304 21684
rect 16356 21632 16362 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 17129 21675 17187 21681
rect 17129 21672 17141 21675
rect 16448 21644 17141 21672
rect 16448 21632 16454 21644
rect 17129 21641 17141 21644
rect 17175 21641 17187 21675
rect 17129 21635 17187 21641
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 17681 21675 17739 21681
rect 17681 21672 17693 21675
rect 17552 21644 17693 21672
rect 17552 21632 17558 21644
rect 17681 21641 17693 21644
rect 17727 21641 17739 21675
rect 18877 21675 18935 21681
rect 18877 21672 18889 21675
rect 17681 21635 17739 21641
rect 17788 21644 18889 21672
rect 13837 21576 14412 21604
rect 13538 21545 13544 21548
rect 12713 21539 12771 21545
rect 12713 21536 12725 21539
rect 12676 21508 12725 21536
rect 12676 21496 12682 21508
rect 12713 21505 12725 21508
rect 12759 21536 12771 21539
rect 12989 21539 13047 21545
rect 12759 21508 12940 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 12912 21480 12940 21508
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13505 21539 13544 21545
rect 13505 21505 13517 21539
rect 13505 21499 13544 21505
rect 9548 21440 11192 21468
rect 11333 21471 11391 21477
rect 9548 21428 9554 21440
rect 11333 21437 11345 21471
rect 11379 21468 11391 21471
rect 11379 21440 12756 21468
rect 11379 21437 11391 21440
rect 11333 21431 11391 21437
rect 12728 21412 12756 21440
rect 12894 21428 12900 21480
rect 12952 21428 12958 21480
rect 8996 21372 9260 21400
rect 8996 21360 9002 21372
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 11974 21400 11980 21412
rect 10652 21372 11980 21400
rect 10652 21360 10658 21372
rect 11974 21360 11980 21372
rect 12032 21360 12038 21412
rect 12066 21360 12072 21412
rect 12124 21400 12130 21412
rect 12124 21372 12572 21400
rect 12124 21360 12130 21372
rect 2498 21332 2504 21344
rect 1912 21304 2504 21332
rect 1912 21292 1918 21304
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 4430 21332 4436 21344
rect 3476 21304 4436 21332
rect 3476 21292 3482 21304
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 4540 21332 4568 21360
rect 4893 21335 4951 21341
rect 4893 21332 4905 21335
rect 4540 21304 4905 21332
rect 4893 21301 4905 21304
rect 4939 21301 4951 21335
rect 4893 21295 4951 21301
rect 7282 21292 7288 21344
rect 7340 21332 7346 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7340 21304 8033 21332
rect 7340 21292 7346 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8665 21335 8723 21341
rect 8665 21301 8677 21335
rect 8711 21332 8723 21335
rect 8846 21332 8852 21344
rect 8711 21304 8852 21332
rect 8711 21301 8723 21304
rect 8665 21295 8723 21301
rect 8846 21292 8852 21304
rect 8904 21292 8910 21344
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9766 21332 9772 21344
rect 9088 21304 9772 21332
rect 9088 21292 9094 21304
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 10410 21292 10416 21344
rect 10468 21332 10474 21344
rect 12434 21332 12440 21344
rect 10468 21304 12440 21332
rect 10468 21292 10474 21304
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 12544 21332 12572 21372
rect 12710 21360 12716 21412
rect 12768 21360 12774 21412
rect 12802 21332 12808 21344
rect 12544 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 13004 21332 13032 21499
rect 13372 21400 13400 21499
rect 13538 21496 13544 21499
rect 13596 21496 13602 21548
rect 13837 21545 13865 21576
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21505 13783 21539
rect 13725 21499 13783 21505
rect 13822 21539 13880 21545
rect 13822 21505 13834 21539
rect 13868 21505 13880 21539
rect 13822 21499 13880 21505
rect 13740 21468 13768 21499
rect 13998 21496 14004 21548
rect 14056 21496 14062 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21536 14151 21539
rect 14274 21536 14280 21548
rect 14139 21508 14280 21536
rect 14139 21505 14151 21508
rect 14093 21499 14151 21505
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 14384 21545 14412 21576
rect 14918 21564 14924 21616
rect 14976 21604 14982 21616
rect 14976 21576 15424 21604
rect 14976 21564 14982 21576
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21536 14427 21539
rect 15010 21536 15016 21548
rect 14415 21508 15016 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 15102 21496 15108 21548
rect 15160 21496 15166 21548
rect 15396 21545 15424 21576
rect 15488 21545 15516 21632
rect 15841 21607 15899 21613
rect 15841 21573 15853 21607
rect 15887 21604 15899 21607
rect 17788 21604 17816 21644
rect 18877 21641 18889 21644
rect 18923 21641 18935 21675
rect 18877 21635 18935 21641
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 21082 21672 21088 21684
rect 19392 21644 21088 21672
rect 19392 21632 19398 21644
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 21269 21675 21327 21681
rect 21269 21641 21281 21675
rect 21315 21672 21327 21675
rect 21358 21672 21364 21684
rect 21315 21644 21364 21672
rect 21315 21641 21327 21644
rect 21269 21635 21327 21641
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 21928 21644 24532 21672
rect 15887 21576 17816 21604
rect 15887 21573 15899 21576
rect 15841 21567 15899 21573
rect 18046 21564 18052 21616
rect 18104 21604 18110 21616
rect 20438 21604 20444 21616
rect 18104 21576 18184 21604
rect 18104 21564 18110 21576
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 16390 21536 16396 21548
rect 16163 21508 16396 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 14016 21468 14044 21496
rect 13740 21440 14044 21468
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21468 14243 21471
rect 14734 21468 14740 21480
rect 14231 21440 14740 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 15212 21468 15240 21499
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16632 21508 16681 21536
rect 16632 21496 16638 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16816 21508 16957 21536
rect 16816 21496 16822 21508
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 17184 21508 17233 21536
rect 17184 21496 17190 21508
rect 17221 21505 17233 21508
rect 17267 21536 17279 21539
rect 17497 21539 17555 21545
rect 17267 21508 17439 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 16025 21471 16083 21477
rect 15212 21440 15424 21468
rect 15286 21400 15292 21412
rect 13372 21372 15292 21400
rect 15286 21360 15292 21372
rect 15344 21360 15350 21412
rect 15396 21400 15424 21440
rect 16025 21437 16037 21471
rect 16071 21468 16083 21471
rect 16298 21468 16304 21480
rect 16071 21440 16304 21468
rect 16071 21437 16083 21440
rect 16025 21431 16083 21437
rect 16298 21428 16304 21440
rect 16356 21428 16362 21480
rect 16408 21468 16436 21496
rect 16776 21468 16804 21496
rect 16408 21440 16804 21468
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21468 16911 21471
rect 17236 21468 17264 21499
rect 16899 21440 17264 21468
rect 17313 21471 17371 21477
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 17313 21437 17325 21471
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 15746 21400 15752 21412
rect 15396 21372 15752 21400
rect 15746 21360 15752 21372
rect 15804 21400 15810 21412
rect 17034 21400 17040 21412
rect 15804 21372 17040 21400
rect 15804 21360 15810 21372
rect 17034 21360 17040 21372
rect 17092 21360 17098 21412
rect 17126 21360 17132 21412
rect 17184 21400 17190 21412
rect 17328 21400 17356 21431
rect 17184 21372 17356 21400
rect 17184 21360 17190 21372
rect 13630 21332 13636 21344
rect 13004 21304 13636 21332
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 13998 21292 14004 21344
rect 14056 21292 14062 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14734 21332 14740 21344
rect 14424 21304 14740 21332
rect 14424 21292 14430 21304
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 14918 21292 14924 21344
rect 14976 21292 14982 21344
rect 15194 21292 15200 21344
rect 15252 21332 15258 21344
rect 15841 21335 15899 21341
rect 15841 21332 15853 21335
rect 15252 21304 15853 21332
rect 15252 21292 15258 21304
rect 15841 21301 15853 21304
rect 15887 21301 15899 21335
rect 15841 21295 15899 21301
rect 16666 21292 16672 21344
rect 16724 21292 16730 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 17411 21332 17439 21508
rect 17497 21505 17509 21539
rect 17543 21536 17555 21539
rect 17678 21536 17684 21548
rect 17543 21508 17684 21536
rect 17543 21505 17555 21508
rect 17497 21499 17555 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 18156 21545 18184 21576
rect 18524 21576 18828 21604
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21505 18199 21539
rect 18141 21499 18199 21505
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 17972 21400 18000 21499
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18432 21468 18460 21499
rect 18524 21477 18552 21576
rect 18800 21548 18828 21576
rect 18892 21576 19472 21604
rect 18690 21496 18696 21548
rect 18748 21496 18754 21548
rect 18782 21496 18788 21548
rect 18840 21496 18846 21548
rect 18104 21440 18460 21468
rect 18509 21471 18567 21477
rect 18104 21428 18110 21440
rect 18509 21437 18521 21471
rect 18555 21437 18567 21471
rect 18509 21431 18567 21437
rect 18892 21400 18920 21576
rect 18966 21496 18972 21548
rect 19024 21496 19030 21548
rect 19150 21496 19156 21548
rect 19208 21496 19214 21548
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21536 19303 21539
rect 19291 21508 19380 21536
rect 19291 21505 19303 21508
rect 19245 21499 19303 21505
rect 19150 21400 19156 21412
rect 17972 21372 18920 21400
rect 19076 21372 19156 21400
rect 17368 21304 17439 21332
rect 17368 21292 17374 21304
rect 17494 21292 17500 21344
rect 17552 21292 17558 21344
rect 17954 21292 17960 21344
rect 18012 21292 18018 21344
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 18325 21335 18383 21341
rect 18325 21332 18337 21335
rect 18104 21304 18337 21332
rect 18104 21292 18110 21304
rect 18325 21301 18337 21304
rect 18371 21301 18383 21335
rect 18325 21295 18383 21301
rect 18506 21292 18512 21344
rect 18564 21292 18570 21344
rect 19076 21341 19104 21372
rect 19150 21360 19156 21372
rect 19208 21360 19214 21412
rect 19352 21344 19380 21508
rect 19444 21409 19472 21576
rect 20180 21576 20444 21604
rect 19610 21496 19616 21548
rect 19668 21536 19674 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19668 21508 19717 21536
rect 19668 21496 19674 21508
rect 19705 21505 19717 21508
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20006 21542 20064 21545
rect 20180 21542 20208 21576
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 20806 21564 20812 21616
rect 20864 21604 20870 21616
rect 20864 21576 21404 21604
rect 20864 21564 20870 21576
rect 21376 21548 21404 21576
rect 21818 21564 21824 21616
rect 21876 21604 21882 21616
rect 21928 21604 21956 21644
rect 21876 21576 21956 21604
rect 21876 21564 21882 21576
rect 22462 21564 22468 21616
rect 22520 21564 22526 21616
rect 22646 21604 22652 21616
rect 22572 21576 22652 21604
rect 20006 21539 20208 21542
rect 20006 21505 20018 21539
rect 20052 21514 20208 21539
rect 20257 21539 20315 21545
rect 20052 21505 20064 21514
rect 20006 21499 20064 21505
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 19429 21403 19487 21409
rect 19429 21369 19441 21403
rect 19475 21369 19487 21403
rect 20272 21400 20300 21499
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21536 20683 21539
rect 21082 21536 21088 21548
rect 20671 21508 21088 21536
rect 20671 21505 20683 21508
rect 20625 21499 20683 21505
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 20548 21468 20576 21496
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20548 21440 20821 21468
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 21192 21468 21220 21499
rect 21358 21496 21364 21548
rect 21416 21496 21422 21548
rect 21542 21496 21548 21548
rect 21600 21496 21606 21548
rect 21910 21496 21916 21548
rect 21968 21496 21974 21548
rect 22186 21496 22192 21548
rect 22244 21496 22250 21548
rect 22572 21545 22600 21576
rect 22646 21564 22652 21576
rect 22704 21604 22710 21616
rect 22704 21576 23244 21604
rect 22704 21564 22710 21576
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 21560 21468 21588 21496
rect 20809 21431 20867 21437
rect 21008 21440 21588 21468
rect 22388 21468 22416 21499
rect 22830 21496 22836 21548
rect 22888 21545 22894 21548
rect 22888 21539 22911 21545
rect 22899 21505 22911 21539
rect 22888 21499 22911 21505
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 22888 21496 22894 21499
rect 22462 21468 22468 21480
rect 22388 21440 22468 21468
rect 19429 21363 19487 21369
rect 20088 21372 20300 21400
rect 20441 21403 20499 21409
rect 19061 21335 19119 21341
rect 19061 21301 19073 21335
rect 19107 21301 19119 21335
rect 19061 21295 19119 21301
rect 19334 21292 19340 21344
rect 19392 21292 19398 21344
rect 19705 21335 19763 21341
rect 19705 21301 19717 21335
rect 19751 21332 19763 21335
rect 19794 21332 19800 21344
rect 19751 21304 19800 21332
rect 19751 21301 19763 21304
rect 19705 21295 19763 21301
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 19886 21292 19892 21344
rect 19944 21332 19950 21344
rect 20088 21332 20116 21372
rect 20441 21369 20453 21403
rect 20487 21400 20499 21403
rect 21008 21400 21036 21440
rect 22462 21428 22468 21440
rect 22520 21468 22526 21480
rect 22738 21468 22744 21480
rect 22520 21440 22744 21468
rect 22520 21428 22526 21440
rect 22738 21428 22744 21440
rect 22796 21468 22802 21480
rect 23032 21468 23060 21499
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23216 21545 23244 21576
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 23842 21604 23848 21616
rect 23624 21576 23848 21604
rect 23624 21564 23630 21576
rect 23842 21564 23848 21576
rect 23900 21604 23906 21616
rect 24504 21613 24532 21644
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25590 21672 25596 21684
rect 24820 21644 25596 21672
rect 24820 21632 24826 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 26605 21675 26663 21681
rect 26007 21644 26188 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 24489 21607 24547 21613
rect 23900 21576 24072 21604
rect 23900 21564 23906 21576
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21505 23259 21539
rect 23201 21499 23259 21505
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21505 23719 21539
rect 23937 21539 23995 21545
rect 23937 21536 23949 21539
rect 23661 21499 23719 21505
rect 23861 21508 23949 21536
rect 22796 21440 23060 21468
rect 22796 21428 22802 21440
rect 20487 21372 21036 21400
rect 20487 21369 20499 21372
rect 20441 21363 20499 21369
rect 19944 21304 20116 21332
rect 19944 21292 19950 21304
rect 20254 21292 20260 21344
rect 20312 21292 20318 21344
rect 22002 21292 22008 21344
rect 22060 21292 22066 21344
rect 22741 21335 22799 21341
rect 22741 21301 22753 21335
rect 22787 21332 22799 21335
rect 22922 21332 22928 21344
rect 22787 21304 22928 21332
rect 22787 21301 22799 21304
rect 22741 21295 22799 21301
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23124 21332 23152 21496
rect 23072 21304 23152 21332
rect 23216 21332 23244 21499
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 23676 21468 23704 21499
rect 23861 21480 23889 21508
rect 23937 21505 23949 21508
rect 23983 21505 23995 21539
rect 23937 21499 23995 21505
rect 23624 21440 23704 21468
rect 23624 21428 23630 21440
rect 23750 21428 23756 21480
rect 23808 21428 23814 21480
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 23385 21403 23443 21409
rect 23385 21369 23397 21403
rect 23431 21400 23443 21403
rect 23861 21400 23889 21428
rect 23431 21372 23889 21400
rect 23431 21369 23443 21372
rect 23385 21363 23443 21369
rect 23842 21332 23848 21344
rect 23216 21304 23848 21332
rect 23072 21292 23078 21304
rect 23842 21292 23848 21304
rect 23900 21292 23906 21344
rect 23937 21335 23995 21341
rect 23937 21301 23949 21335
rect 23983 21332 23995 21335
rect 24044 21332 24072 21576
rect 24489 21573 24501 21607
rect 24535 21573 24547 21607
rect 24489 21567 24547 21573
rect 24578 21564 24584 21616
rect 24636 21564 24642 21616
rect 25501 21607 25559 21613
rect 25501 21573 25513 21607
rect 25547 21604 25559 21607
rect 26050 21604 26056 21616
rect 25547 21576 26056 21604
rect 25547 21573 25559 21576
rect 25501 21567 25559 21573
rect 26050 21564 26056 21576
rect 26108 21564 26114 21616
rect 26160 21613 26188 21644
rect 26605 21641 26617 21675
rect 26651 21672 26663 21675
rect 26970 21672 26976 21684
rect 26651 21644 26976 21672
rect 26651 21641 26663 21644
rect 26605 21635 26663 21641
rect 26970 21632 26976 21644
rect 27028 21632 27034 21684
rect 27062 21632 27068 21684
rect 27120 21672 27126 21684
rect 27338 21672 27344 21684
rect 27120 21644 27344 21672
rect 27120 21632 27126 21644
rect 27338 21632 27344 21644
rect 27396 21632 27402 21684
rect 26145 21607 26203 21613
rect 26145 21573 26157 21607
rect 26191 21573 26203 21607
rect 26145 21567 26203 21573
rect 26326 21564 26332 21616
rect 26384 21564 26390 21616
rect 26620 21576 27292 21604
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 24305 21539 24363 21545
rect 24305 21536 24317 21539
rect 24176 21508 24317 21536
rect 24176 21496 24182 21508
rect 24305 21505 24317 21508
rect 24351 21505 24363 21539
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 24305 21499 24363 21505
rect 24504 21508 24685 21536
rect 24504 21480 24532 21508
rect 24673 21505 24685 21508
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 25774 21496 25780 21548
rect 25832 21496 25838 21548
rect 25866 21496 25872 21548
rect 25924 21536 25930 21548
rect 26344 21536 26372 21564
rect 26620 21548 26648 21576
rect 26421 21539 26479 21545
rect 26421 21536 26433 21539
rect 25924 21508 26433 21536
rect 25924 21496 25930 21508
rect 26421 21505 26433 21508
rect 26467 21505 26479 21539
rect 26421 21499 26479 21505
rect 26602 21496 26608 21548
rect 26660 21496 26666 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27264 21545 27292 21576
rect 27908 21576 28764 21604
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 27430 21496 27436 21548
rect 27488 21536 27494 21548
rect 27908 21545 27936 21576
rect 28736 21548 28764 21576
rect 27709 21539 27767 21545
rect 27709 21536 27721 21539
rect 27488 21508 27721 21536
rect 27488 21496 27494 21508
rect 27709 21505 27721 21508
rect 27755 21505 27767 21539
rect 27709 21499 27767 21505
rect 27893 21539 27951 21545
rect 27893 21505 27905 21539
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 27985 21539 28043 21545
rect 27985 21505 27997 21539
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 24486 21428 24492 21480
rect 24544 21428 24550 21480
rect 24854 21428 24860 21480
rect 24912 21428 24918 21480
rect 24946 21428 24952 21480
rect 25004 21468 25010 21480
rect 25593 21471 25651 21477
rect 25593 21468 25605 21471
rect 25004 21440 25605 21468
rect 25004 21428 25010 21440
rect 25593 21437 25605 21440
rect 25639 21437 25651 21471
rect 25593 21431 25651 21437
rect 26329 21471 26387 21477
rect 26329 21437 26341 21471
rect 26375 21468 26387 21471
rect 26786 21468 26792 21480
rect 26375 21440 26792 21468
rect 26375 21437 26387 21440
rect 26329 21431 26387 21437
rect 26786 21428 26792 21440
rect 26844 21428 26850 21480
rect 27065 21471 27123 21477
rect 27065 21437 27077 21471
rect 27111 21437 27123 21471
rect 28000 21468 28028 21499
rect 28258 21496 28264 21548
rect 28316 21545 28322 21548
rect 28316 21536 28324 21545
rect 28445 21539 28503 21545
rect 28316 21508 28361 21536
rect 28316 21499 28324 21508
rect 28445 21505 28457 21539
rect 28491 21536 28503 21539
rect 28626 21536 28632 21548
rect 28491 21508 28632 21536
rect 28491 21505 28503 21508
rect 28445 21499 28503 21505
rect 28316 21496 28322 21499
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 28718 21496 28724 21548
rect 28776 21496 28782 21548
rect 28534 21468 28540 21480
rect 28000 21440 28540 21468
rect 27065 21431 27123 21437
rect 24121 21403 24179 21409
rect 24121 21369 24133 21403
rect 24167 21369 24179 21403
rect 24872 21400 24900 21428
rect 26694 21400 26700 21412
rect 24121 21363 24179 21369
rect 24786 21372 24900 21400
rect 25700 21372 26700 21400
rect 23983 21304 24072 21332
rect 24136 21332 24164 21363
rect 24786 21332 24814 21372
rect 24136 21304 24814 21332
rect 24857 21335 24915 21341
rect 23983 21301 23995 21304
rect 23937 21295 23995 21301
rect 24857 21301 24869 21335
rect 24903 21332 24915 21335
rect 25700 21332 25728 21372
rect 26694 21360 26700 21372
rect 26752 21400 26758 21412
rect 27080 21400 27108 21431
rect 28534 21428 28540 21440
rect 28592 21428 28598 21480
rect 28350 21400 28356 21412
rect 26752 21372 27108 21400
rect 28000 21372 28356 21400
rect 26752 21360 26758 21372
rect 24903 21304 25728 21332
rect 25777 21335 25835 21341
rect 24903 21301 24915 21304
rect 24857 21295 24915 21301
rect 25777 21301 25789 21335
rect 25823 21332 25835 21335
rect 25866 21332 25872 21344
rect 25823 21304 25872 21332
rect 25823 21301 25835 21304
rect 25777 21295 25835 21301
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 26418 21292 26424 21344
rect 26476 21292 26482 21344
rect 27154 21292 27160 21344
rect 27212 21292 27218 21344
rect 27433 21335 27491 21341
rect 27433 21301 27445 21335
rect 27479 21332 27491 21335
rect 27706 21332 27712 21344
rect 27479 21304 27712 21332
rect 27479 21301 27491 21304
rect 27433 21295 27491 21301
rect 27706 21292 27712 21304
rect 27764 21292 27770 21344
rect 28000 21341 28028 21372
rect 28350 21360 28356 21372
rect 28408 21400 28414 21412
rect 28629 21403 28687 21409
rect 28629 21400 28641 21403
rect 28408 21372 28641 21400
rect 28408 21360 28414 21372
rect 28629 21369 28641 21372
rect 28675 21369 28687 21403
rect 28629 21363 28687 21369
rect 27985 21335 28043 21341
rect 27985 21301 27997 21335
rect 28031 21301 28043 21335
rect 27985 21295 28043 21301
rect 28166 21292 28172 21344
rect 28224 21292 28230 21344
rect 28445 21335 28503 21341
rect 28445 21301 28457 21335
rect 28491 21332 28503 21335
rect 29178 21332 29184 21344
rect 28491 21304 29184 21332
rect 28491 21301 28503 21304
rect 28445 21295 28503 21301
rect 29178 21292 29184 21304
rect 29236 21292 29242 21344
rect 1104 21242 43884 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 43884 21242
rect 1104 21168 43884 21190
rect 2130 21088 2136 21140
rect 2188 21128 2194 21140
rect 2774 21128 2780 21140
rect 2188 21100 2780 21128
rect 2188 21088 2194 21100
rect 2774 21088 2780 21100
rect 2832 21088 2838 21140
rect 2958 21088 2964 21140
rect 3016 21128 3022 21140
rect 3605 21131 3663 21137
rect 3605 21128 3617 21131
rect 3016 21100 3617 21128
rect 3016 21088 3022 21100
rect 3605 21097 3617 21100
rect 3651 21097 3663 21131
rect 5353 21131 5411 21137
rect 5353 21128 5365 21131
rect 3605 21091 3663 21097
rect 5000 21100 5365 21128
rect 5000 21060 5028 21100
rect 5353 21097 5365 21100
rect 5399 21097 5411 21131
rect 5353 21091 5411 21097
rect 5457 21100 5764 21128
rect 5457 21060 5485 21100
rect 3068 21032 5028 21060
rect 5093 21032 5485 21060
rect 1210 20952 1216 21004
rect 1268 20992 1274 21004
rect 1857 20995 1915 21001
rect 1857 20992 1869 20995
rect 1268 20964 1869 20992
rect 1268 20952 1274 20964
rect 1857 20961 1869 20964
rect 1903 20961 1915 20995
rect 1857 20955 1915 20961
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 1946 20924 1952 20936
rect 1627 20896 1952 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 3068 20933 3096 21032
rect 3602 20992 3608 21004
rect 3436 20964 3608 20992
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20893 3111 20927
rect 3053 20887 3111 20893
rect 3234 20884 3240 20936
rect 3292 20884 3298 20936
rect 3326 20884 3332 20936
rect 3384 20884 3390 20936
rect 3436 20933 3464 20964
rect 3602 20952 3608 20964
rect 3660 20952 3666 21004
rect 4341 20995 4399 21001
rect 4341 20992 4353 20995
rect 3712 20964 4353 20992
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 1670 20816 1676 20868
rect 1728 20816 1734 20868
rect 3344 20856 3372 20884
rect 3712 20856 3740 20964
rect 4341 20961 4353 20964
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4706 20952 4712 21004
rect 4764 20992 4770 21004
rect 4801 20995 4859 21001
rect 4801 20992 4813 20995
rect 4764 20964 4813 20992
rect 4764 20952 4770 20964
rect 4801 20961 4813 20964
rect 4847 20992 4859 20995
rect 5093 20992 5121 21032
rect 5534 21020 5540 21072
rect 5592 21020 5598 21072
rect 5626 21020 5632 21072
rect 5684 21020 5690 21072
rect 5736 21060 5764 21100
rect 5994 21088 6000 21140
rect 6052 21128 6058 21140
rect 6730 21128 6736 21140
rect 6052 21100 6736 21128
rect 6052 21088 6058 21100
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 6914 21128 6920 21140
rect 6840 21100 6920 21128
rect 6270 21060 6276 21072
rect 5736 21032 6276 21060
rect 6270 21020 6276 21032
rect 6328 21060 6334 21072
rect 6840 21060 6868 21100
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 7282 21128 7288 21140
rect 7024 21100 7288 21128
rect 7024 21060 7052 21100
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 7834 21128 7840 21140
rect 7524 21100 7840 21128
rect 7524 21088 7530 21100
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 7926 21088 7932 21140
rect 7984 21128 7990 21140
rect 8757 21131 8815 21137
rect 8757 21128 8769 21131
rect 7984 21100 8769 21128
rect 7984 21088 7990 21100
rect 8757 21097 8769 21100
rect 8803 21097 8815 21131
rect 10226 21128 10232 21140
rect 8757 21091 8815 21097
rect 9278 21100 10232 21128
rect 6328 21032 6500 21060
rect 6328 21020 6334 21032
rect 4847 20964 5121 20992
rect 5169 20995 5227 21001
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 5169 20961 5181 20995
rect 5215 20992 5227 20995
rect 5350 20992 5356 21004
rect 5215 20964 5356 20992
rect 5215 20961 5227 20964
rect 5169 20955 5227 20961
rect 5350 20952 5356 20964
rect 5408 20992 5414 21004
rect 5552 20992 5580 21020
rect 5408 20964 5580 20992
rect 5644 20992 5672 21020
rect 6365 20995 6423 21001
rect 6365 20992 6377 20995
rect 5644 20964 6377 20992
rect 5408 20952 5414 20964
rect 6365 20961 6377 20964
rect 6411 20961 6423 20995
rect 6365 20955 6423 20961
rect 3786 20884 3792 20936
rect 3844 20884 3850 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 4522 20884 4528 20936
rect 4580 20884 4586 20936
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 4724 20896 4905 20924
rect 3344 20828 3740 20856
rect 3804 20856 3832 20884
rect 4724 20868 4752 20896
rect 4893 20893 4905 20896
rect 4939 20893 4951 20927
rect 5629 20927 5687 20933
rect 5629 20924 5641 20927
rect 5368 20920 5641 20924
rect 4893 20887 4951 20893
rect 4992 20896 5641 20920
rect 4992 20892 5396 20896
rect 5629 20893 5641 20896
rect 5675 20893 5687 20927
rect 4157 20859 4215 20865
rect 4157 20856 4169 20859
rect 3804 20828 4169 20856
rect 4157 20825 4169 20828
rect 4203 20825 4215 20859
rect 4157 20819 4215 20825
rect 1688 20788 1716 20816
rect 3418 20788 3424 20800
rect 1688 20760 3424 20788
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 4172 20788 4200 20819
rect 4706 20816 4712 20868
rect 4764 20816 4770 20868
rect 4992 20788 5020 20892
rect 5629 20887 5687 20893
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6472 20933 6500 21032
rect 6656 21032 6868 21060
rect 6896 21032 7052 21060
rect 6656 20933 6684 21032
rect 6896 20992 6924 21032
rect 7374 21020 7380 21072
rect 7432 21020 7438 21072
rect 9278 21060 9306 21100
rect 10226 21088 10232 21100
rect 10284 21088 10290 21140
rect 10318 21088 10324 21140
rect 10376 21088 10382 21140
rect 10410 21088 10416 21140
rect 10468 21128 10474 21140
rect 10778 21128 10784 21140
rect 10468 21100 10784 21128
rect 10468 21088 10474 21100
rect 10778 21088 10784 21100
rect 10836 21128 10842 21140
rect 11885 21131 11943 21137
rect 10836 21100 11468 21128
rect 10836 21088 10842 21100
rect 10336 21060 10364 21088
rect 7484 21032 9306 21060
rect 9692 21032 11054 21060
rect 7484 20992 7512 21032
rect 6748 20964 6924 20992
rect 7024 20964 7512 20992
rect 7561 20995 7619 21001
rect 6748 20933 6776 20964
rect 7024 20936 7052 20964
rect 7561 20961 7573 20995
rect 7607 20992 7619 20995
rect 7742 20992 7748 21004
rect 7607 20964 7748 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 7742 20952 7748 20964
rect 7800 20952 7806 21004
rect 8018 20952 8024 21004
rect 8076 20952 8082 21004
rect 6914 20934 6920 20936
rect 6840 20933 6920 20934
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 6641 20927 6699 20933
rect 6641 20893 6653 20927
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 6733 20927 6791 20933
rect 6733 20893 6745 20927
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 6826 20927 6920 20933
rect 6826 20893 6838 20927
rect 6872 20906 6920 20927
rect 6872 20893 6884 20906
rect 6826 20887 6884 20893
rect 6914 20884 6920 20906
rect 6972 20884 6978 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 7190 20884 7196 20936
rect 7248 20933 7254 20936
rect 7248 20924 7256 20933
rect 8036 20924 8064 20952
rect 7248 20896 7293 20924
rect 7489 20896 8064 20924
rect 8205 20927 8263 20933
rect 7248 20887 7256 20896
rect 7248 20884 7254 20887
rect 5534 20816 5540 20868
rect 5592 20816 5598 20868
rect 7489 20856 7517 20896
rect 8205 20893 8217 20927
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 5920 20828 7517 20856
rect 5920 20800 5948 20828
rect 8018 20816 8024 20868
rect 8076 20856 8082 20868
rect 8220 20856 8248 20887
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 8481 20927 8539 20933
rect 8481 20926 8493 20927
rect 8408 20924 8493 20926
rect 8352 20898 8493 20924
rect 8352 20896 8436 20898
rect 8352 20884 8358 20896
rect 8481 20893 8493 20898
rect 8527 20893 8539 20927
rect 8481 20887 8539 20893
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 8076 20828 8248 20856
rect 8076 20816 8082 20828
rect 8386 20816 8392 20868
rect 8444 20816 8450 20868
rect 8588 20856 8616 20887
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 8941 20927 8999 20933
rect 8904 20920 8913 20924
rect 8941 20920 8953 20927
rect 8904 20893 8953 20920
rect 8987 20893 8999 20927
rect 8904 20892 8999 20893
rect 8904 20884 8910 20892
rect 8941 20887 8999 20892
rect 9030 20884 9036 20936
rect 9088 20884 9094 20936
rect 9232 20933 9260 21032
rect 9582 20992 9588 21004
rect 9324 20964 9588 20992
rect 9324 20933 9352 20964
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9217 20927 9275 20933
rect 9217 20893 9229 20927
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9398 20884 9404 20936
rect 9456 20933 9462 20936
rect 9456 20924 9464 20933
rect 9692 20924 9720 21032
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 11026 20992 11054 21032
rect 11146 21020 11152 21072
rect 11204 21020 11210 21072
rect 11164 20992 11192 21020
rect 10376 20964 10732 20992
rect 10376 20952 10382 20964
rect 9456 20896 9720 20924
rect 9769 20927 9827 20933
rect 9456 20887 9464 20896
rect 9769 20893 9781 20927
rect 9815 20924 9827 20927
rect 9858 20924 9864 20936
rect 9815 20896 9864 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 9456 20884 9462 20887
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 10042 20884 10048 20936
rect 10100 20884 10106 20936
rect 10704 20933 10732 20964
rect 10893 20964 11192 20992
rect 10893 20933 10921 20964
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20926 10195 20927
rect 10413 20927 10471 20933
rect 10183 20898 10272 20926
rect 10413 20924 10425 20927
rect 10183 20893 10195 20898
rect 10137 20887 10195 20893
rect 10244 20868 10272 20898
rect 10336 20896 10425 20924
rect 9490 20856 9496 20868
rect 8588 20828 9496 20856
rect 9490 20816 9496 20828
rect 9548 20816 9554 20868
rect 9953 20859 10011 20865
rect 9953 20856 9965 20859
rect 9784 20828 9965 20856
rect 9784 20800 9812 20828
rect 9953 20825 9965 20828
rect 9999 20825 10011 20859
rect 9953 20819 10011 20825
rect 10226 20816 10232 20868
rect 10284 20816 10290 20868
rect 4172 20760 5020 20788
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5902 20788 5908 20800
rect 5132 20760 5908 20788
rect 5132 20748 5138 20760
rect 5902 20748 5908 20760
rect 5960 20748 5966 20800
rect 6641 20791 6699 20797
rect 6641 20757 6653 20791
rect 6687 20788 6699 20791
rect 6822 20788 6828 20800
rect 6687 20760 6828 20788
rect 6687 20757 6699 20760
rect 6641 20751 6699 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 6914 20748 6920 20800
rect 6972 20788 6978 20800
rect 7282 20788 7288 20800
rect 6972 20760 7288 20788
rect 6972 20748 6978 20760
rect 7282 20748 7288 20760
rect 7340 20788 7346 20800
rect 8113 20791 8171 20797
rect 8113 20788 8125 20791
rect 7340 20760 8125 20788
rect 7340 20748 7346 20760
rect 8113 20757 8125 20760
rect 8159 20757 8171 20791
rect 8113 20751 8171 20757
rect 9582 20748 9588 20800
rect 9640 20748 9646 20800
rect 9766 20748 9772 20800
rect 9824 20748 9830 20800
rect 10336 20797 10364 20896
rect 10413 20893 10425 20896
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 10561 20927 10619 20933
rect 10561 20893 10573 20927
rect 10607 20924 10619 20927
rect 10689 20927 10747 20933
rect 10607 20893 10640 20924
rect 10561 20887 10640 20893
rect 10689 20893 10701 20927
rect 10735 20893 10747 20927
rect 10689 20887 10747 20893
rect 10878 20927 10936 20933
rect 10878 20893 10890 20927
rect 10924 20893 10936 20927
rect 10878 20887 10936 20893
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20757 10379 20791
rect 10612 20788 10640 20887
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11440 20933 11468 21100
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 12250 21128 12256 21140
rect 11931 21100 12256 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12345 21131 12403 21137
rect 12345 21097 12357 21131
rect 12391 21128 12403 21131
rect 12618 21128 12624 21140
rect 12391 21100 12624 21128
rect 12391 21097 12403 21100
rect 12345 21091 12403 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 12728 21100 16957 21128
rect 12728 20992 12756 21100
rect 16945 21097 16957 21100
rect 16991 21097 17003 21131
rect 16945 21091 17003 21097
rect 17313 21131 17371 21137
rect 17313 21097 17325 21131
rect 17359 21128 17371 21131
rect 17494 21128 17500 21140
rect 17359 21100 17500 21128
rect 17359 21097 17371 21100
rect 17313 21091 17371 21097
rect 17494 21088 17500 21100
rect 17552 21088 17558 21140
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 18748 21100 19564 21128
rect 18748 21088 18754 21100
rect 14737 21063 14795 21069
rect 14737 21060 14749 21063
rect 13096 21032 14749 21060
rect 13096 21004 13124 21032
rect 14737 21029 14749 21032
rect 14783 21029 14795 21063
rect 14737 21023 14795 21029
rect 14918 21020 14924 21072
rect 14976 21020 14982 21072
rect 17218 21020 17224 21072
rect 17276 21060 17282 21072
rect 17957 21063 18015 21069
rect 17957 21060 17969 21063
rect 17276 21032 17969 21060
rect 17276 21020 17282 21032
rect 17957 21029 17969 21032
rect 18003 21029 18015 21063
rect 17957 21023 18015 21029
rect 18233 21063 18291 21069
rect 18233 21029 18245 21063
rect 18279 21029 18291 21063
rect 18233 21023 18291 21029
rect 18325 21063 18383 21069
rect 18325 21029 18337 21063
rect 18371 21060 18383 21063
rect 18506 21060 18512 21072
rect 18371 21032 18512 21060
rect 18371 21029 18383 21032
rect 18325 21023 18383 21029
rect 12452 20964 12756 20992
rect 12897 20995 12955 21001
rect 12452 20933 12480 20964
rect 12897 20961 12909 20995
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 11112 20896 11253 20924
rect 11112 20884 11118 20896
rect 11241 20893 11253 20896
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 10778 20816 10784 20868
rect 10836 20816 10842 20868
rect 11256 20856 11284 20887
rect 12452 20856 12480 20887
rect 12618 20884 12624 20936
rect 12676 20884 12682 20936
rect 12912 20856 12940 20955
rect 13078 20952 13084 21004
rect 13136 20952 13142 21004
rect 14936 20992 14964 21020
rect 16577 20995 16635 21001
rect 16577 20992 16589 20995
rect 13556 20964 14964 20992
rect 15672 20964 16589 20992
rect 12986 20884 12992 20936
rect 13044 20884 13050 20936
rect 13170 20884 13176 20936
rect 13228 20884 13234 20936
rect 13556 20933 13584 20964
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14093 20927 14151 20933
rect 13872 20896 14044 20924
rect 13872 20884 13878 20896
rect 14016 20868 14044 20896
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14645 20927 14703 20933
rect 14139 20896 14228 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14200 20868 14228 20896
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 11256 20828 12480 20856
rect 12544 20828 12940 20856
rect 10962 20788 10968 20800
rect 10612 20760 10968 20788
rect 10321 20751 10379 20757
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11054 20748 11060 20800
rect 11112 20748 11118 20800
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11514 20788 11520 20800
rect 11471 20760 11520 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 11606 20748 11612 20800
rect 11664 20788 11670 20800
rect 12066 20788 12072 20800
rect 11664 20760 12072 20788
rect 11664 20748 11670 20760
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 12158 20748 12164 20800
rect 12216 20788 12222 20800
rect 12544 20797 12572 20828
rect 13998 20816 14004 20868
rect 14056 20816 14062 20868
rect 14182 20816 14188 20868
rect 14240 20816 14246 20868
rect 14369 20859 14427 20865
rect 14369 20825 14381 20859
rect 14415 20856 14427 20859
rect 14458 20856 14464 20868
rect 14415 20828 14464 20856
rect 14415 20825 14427 20828
rect 14369 20819 14427 20825
rect 14458 20816 14464 20828
rect 14516 20816 14522 20868
rect 14660 20856 14688 20887
rect 14826 20884 14832 20936
rect 14884 20884 14890 20936
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 15672 20933 15700 20964
rect 16577 20961 16589 20964
rect 16623 20961 16635 20995
rect 17586 20992 17592 21004
rect 16577 20955 16635 20961
rect 17236 20964 17592 20992
rect 17236 20936 17264 20964
rect 17586 20952 17592 20964
rect 17644 20992 17650 21004
rect 17644 20964 17908 20992
rect 17644 20952 17650 20964
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 15488 20856 15516 20887
rect 16022 20884 16028 20936
rect 16080 20884 16086 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 16114 20856 16120 20868
rect 14660 20828 14964 20856
rect 15488 20828 16120 20856
rect 14936 20800 14964 20828
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16298 20816 16304 20868
rect 16356 20856 16362 20868
rect 16482 20856 16488 20868
rect 16356 20828 16488 20856
rect 16356 20816 16362 20828
rect 16482 20816 16488 20828
rect 16540 20856 16546 20868
rect 16669 20859 16727 20865
rect 16669 20856 16681 20859
rect 16540 20828 16681 20856
rect 16540 20816 16546 20828
rect 16669 20825 16681 20828
rect 16715 20825 16727 20859
rect 16669 20819 16727 20825
rect 12529 20791 12587 20797
rect 12529 20788 12541 20791
rect 12216 20760 12541 20788
rect 12216 20748 12222 20760
rect 12529 20757 12541 20760
rect 12575 20757 12587 20791
rect 12529 20751 12587 20757
rect 12710 20748 12716 20800
rect 12768 20748 12774 20800
rect 12894 20748 12900 20800
rect 12952 20788 12958 20800
rect 13357 20791 13415 20797
rect 13357 20788 13369 20791
rect 12952 20760 13369 20788
rect 12952 20748 12958 20760
rect 13357 20757 13369 20760
rect 13403 20757 13415 20791
rect 13357 20751 13415 20757
rect 13725 20791 13783 20797
rect 13725 20757 13737 20791
rect 13771 20788 13783 20791
rect 13814 20788 13820 20800
rect 13771 20760 13820 20788
rect 13771 20757 13783 20760
rect 13725 20751 13783 20757
rect 13814 20748 13820 20760
rect 13872 20788 13878 20800
rect 14826 20788 14832 20800
rect 13872 20760 14832 20788
rect 13872 20748 13878 20760
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 14918 20748 14924 20800
rect 14976 20748 14982 20800
rect 15010 20748 15016 20800
rect 15068 20748 15074 20800
rect 15381 20791 15439 20797
rect 15381 20757 15393 20791
rect 15427 20788 15439 20791
rect 15841 20791 15899 20797
rect 15841 20788 15853 20791
rect 15427 20760 15853 20788
rect 15427 20757 15439 20760
rect 15381 20751 15439 20757
rect 15841 20757 15853 20760
rect 15887 20788 15899 20791
rect 15930 20788 15936 20800
rect 15887 20760 15936 20788
rect 15887 20757 15899 20760
rect 15841 20751 15899 20757
rect 15930 20748 15936 20760
rect 15988 20748 15994 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 16868 20788 16896 20887
rect 17218 20884 17224 20936
rect 17276 20884 17282 20936
rect 17880 20933 17908 20964
rect 18046 20952 18052 21004
rect 18104 20952 18110 21004
rect 18248 20992 18276 21023
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 19536 21060 19564 21100
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 20533 21131 20591 21137
rect 20533 21128 20545 21131
rect 19720 21100 20545 21128
rect 19720 21060 19748 21100
rect 20533 21097 20545 21100
rect 20579 21128 20591 21131
rect 21726 21128 21732 21140
rect 20579 21100 20760 21128
rect 20579 21097 20591 21100
rect 20533 21091 20591 21097
rect 20732 21069 20760 21100
rect 20824 21100 21732 21128
rect 19536 21032 19748 21060
rect 20717 21063 20775 21069
rect 20717 21029 20729 21063
rect 20763 21029 20775 21063
rect 20717 21023 20775 21029
rect 18248 20964 19104 20992
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 17773 20927 17831 20933
rect 17543 20896 17724 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 17328 20856 17356 20887
rect 17328 20828 17632 20856
rect 17604 20800 17632 20828
rect 16632 20760 16896 20788
rect 16632 20748 16638 20760
rect 17586 20748 17592 20800
rect 17644 20748 17650 20800
rect 17696 20788 17724 20896
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 18064 20924 18092 20952
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 18064 20896 18245 20924
rect 17865 20887 17923 20893
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18233 20887 18291 20893
rect 18340 20896 18705 20924
rect 17788 20856 17816 20887
rect 18046 20856 18052 20868
rect 17788 20828 18052 20856
rect 18046 20816 18052 20828
rect 18104 20816 18110 20868
rect 18138 20816 18144 20868
rect 18196 20856 18202 20868
rect 18340 20856 18368 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 18782 20884 18788 20936
rect 18840 20884 18846 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 18966 20924 18972 20936
rect 18923 20896 18972 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19076 20924 19104 20964
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 20073 20995 20131 21001
rect 20073 20992 20085 20995
rect 19484 20964 20085 20992
rect 19484 20952 19490 20964
rect 20073 20961 20085 20964
rect 20119 20992 20131 20995
rect 20824 20992 20852 21100
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 21818 21088 21824 21140
rect 21876 21088 21882 21140
rect 22002 21088 22008 21140
rect 22060 21088 22066 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 23109 21131 23167 21137
rect 22244 21100 22968 21128
rect 22244 21088 22250 21100
rect 20990 21020 20996 21072
rect 21048 21060 21054 21072
rect 21453 21063 21511 21069
rect 21453 21060 21465 21063
rect 21048 21032 21465 21060
rect 21048 21020 21054 21032
rect 21453 21029 21465 21032
rect 21499 21029 21511 21063
rect 21453 21023 21511 21029
rect 21174 20992 21180 21004
rect 20119 20964 20852 20992
rect 21008 20964 21180 20992
rect 20119 20961 20131 20964
rect 20073 20955 20131 20961
rect 19334 20924 19340 20936
rect 19076 20896 19340 20924
rect 19334 20884 19340 20896
rect 19392 20924 19398 20936
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19392 20896 19533 20924
rect 19392 20884 19398 20896
rect 19521 20893 19533 20896
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19713 20924 19771 20927
rect 19713 20921 19840 20924
rect 19713 20887 19725 20921
rect 19759 20896 19840 20921
rect 19759 20887 19771 20896
rect 19713 20881 19771 20887
rect 18196 20828 18368 20856
rect 18509 20859 18567 20865
rect 18196 20816 18202 20828
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 18598 20856 18604 20868
rect 18555 20828 18604 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 18598 20816 18604 20828
rect 18656 20856 18662 20868
rect 19812 20856 19840 20896
rect 19886 20884 19892 20936
rect 19944 20924 19950 20936
rect 20165 20927 20223 20933
rect 20165 20924 20177 20927
rect 19944 20896 20177 20924
rect 19944 20884 19950 20896
rect 20165 20893 20177 20896
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20622 20884 20628 20936
rect 20680 20884 20686 20936
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20924 20959 20927
rect 21008 20924 21036 20964
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 21376 20964 21680 20992
rect 21376 20924 21404 20964
rect 20947 20896 21036 20924
rect 21100 20896 21404 20924
rect 21453 20927 21511 20933
rect 20947 20893 20959 20896
rect 20901 20887 20959 20893
rect 20254 20856 20260 20868
rect 18656 20828 19656 20856
rect 19812 20828 20260 20856
rect 18656 20816 18662 20828
rect 18414 20788 18420 20800
rect 17696 20760 18420 20788
rect 18414 20748 18420 20760
rect 18472 20788 18478 20800
rect 18966 20788 18972 20800
rect 18472 20760 18972 20788
rect 18472 20748 18478 20760
rect 18966 20748 18972 20760
rect 19024 20788 19030 20800
rect 19518 20788 19524 20800
rect 19024 20760 19524 20788
rect 19024 20748 19030 20760
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 19628 20788 19656 20828
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 21100 20856 21128 20896
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 21542 20924 21548 20936
rect 21499 20896 21548 20924
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 21652 20933 21680 20964
rect 22020 20933 22048 21088
rect 22830 21020 22836 21072
rect 22888 21020 22894 21072
rect 22738 20952 22744 21004
rect 22796 20952 22802 21004
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22186 20924 22192 20936
rect 22143 20896 22192 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 22186 20884 22192 20896
rect 22244 20884 22250 20936
rect 22278 20884 22284 20936
rect 22336 20884 22342 20936
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20893 22431 20927
rect 22373 20887 22431 20893
rect 20732 20828 21128 20856
rect 19794 20788 19800 20800
rect 19628 20760 19800 20788
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 20070 20748 20076 20800
rect 20128 20788 20134 20800
rect 20622 20788 20628 20800
rect 20128 20760 20628 20788
rect 20128 20748 20134 20760
rect 20622 20748 20628 20760
rect 20680 20788 20686 20800
rect 20732 20788 20760 20828
rect 21174 20816 21180 20868
rect 21232 20856 21238 20868
rect 22388 20856 22416 20887
rect 22462 20884 22468 20936
rect 22520 20884 22526 20936
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 22756 20924 22784 20952
rect 22848 20933 22876 21020
rect 22940 20992 22968 21100
rect 23109 21097 23121 21131
rect 23155 21128 23167 21131
rect 23290 21128 23296 21140
rect 23155 21100 23296 21128
rect 23155 21097 23167 21100
rect 23109 21091 23167 21097
rect 23290 21088 23296 21100
rect 23348 21128 23354 21140
rect 23474 21128 23480 21140
rect 23348 21100 23480 21128
rect 23348 21088 23354 21100
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 24029 21131 24087 21137
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24394 21128 24400 21140
rect 24075 21100 24400 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 24826 21100 25176 21128
rect 23492 21060 23520 21088
rect 24826 21060 24854 21100
rect 23492 21032 24854 21060
rect 22940 20964 23520 20992
rect 22603 20896 22784 20924
rect 22833 20927 22891 20933
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 22833 20893 22845 20927
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 22925 20927 22983 20933
rect 22925 20893 22937 20927
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 21232 20828 22416 20856
rect 22480 20856 22508 20884
rect 22741 20859 22799 20865
rect 22741 20856 22753 20859
rect 22480 20828 22753 20856
rect 21232 20816 21238 20828
rect 22741 20825 22753 20828
rect 22787 20825 22799 20859
rect 22741 20819 22799 20825
rect 22940 20856 22968 20887
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 23164 20896 23213 20924
rect 23164 20884 23170 20896
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 23492 20933 23520 20964
rect 23860 20964 24926 20992
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 23584 20856 23612 20887
rect 23860 20868 23888 20964
rect 24898 20936 24926 20964
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23992 20896 24409 20924
rect 23992 20884 23998 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 24490 20927 24548 20933
rect 24490 20893 24502 20927
rect 24536 20893 24548 20927
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24490 20887 24548 20893
rect 24596 20896 24777 20924
rect 23842 20856 23848 20868
rect 22940 20828 23848 20856
rect 20680 20760 20760 20788
rect 20680 20748 20686 20760
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21085 20791 21143 20797
rect 21085 20788 21097 20791
rect 20864 20760 21097 20788
rect 20864 20748 20870 20760
rect 21085 20757 21097 20760
rect 21131 20757 21143 20791
rect 21085 20751 21143 20757
rect 22278 20748 22284 20800
rect 22336 20788 22342 20800
rect 22940 20788 22968 20828
rect 23842 20816 23848 20828
rect 23900 20816 23906 20868
rect 24026 20816 24032 20868
rect 24084 20865 24090 20868
rect 24084 20859 24103 20865
rect 24091 20825 24103 20859
rect 24505 20856 24533 20887
rect 24084 20819 24103 20825
rect 24136 20828 24533 20856
rect 24084 20816 24090 20819
rect 22336 20760 22968 20788
rect 22336 20748 22342 20760
rect 23658 20748 23664 20800
rect 23716 20788 23722 20800
rect 23753 20791 23811 20797
rect 23753 20788 23765 20791
rect 23716 20760 23765 20788
rect 23716 20748 23722 20760
rect 23753 20757 23765 20760
rect 23799 20757 23811 20791
rect 23753 20751 23811 20757
rect 23934 20748 23940 20800
rect 23992 20788 23998 20800
rect 24136 20788 24164 20828
rect 23992 20760 24164 20788
rect 23992 20748 23998 20760
rect 24210 20748 24216 20800
rect 24268 20748 24274 20800
rect 24486 20748 24492 20800
rect 24544 20788 24550 20800
rect 24596 20788 24624 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24854 20884 24860 20936
rect 24912 20933 24926 20936
rect 25148 20933 25176 21100
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 26513 21131 26571 21137
rect 26513 21128 26525 21131
rect 26252 21100 26525 21128
rect 25866 21020 25872 21072
rect 25924 21060 25930 21072
rect 26252 21060 26280 21100
rect 26513 21097 26525 21100
rect 26559 21097 26571 21131
rect 26513 21091 26571 21097
rect 27246 21088 27252 21140
rect 27304 21088 27310 21140
rect 27338 21088 27344 21140
rect 27396 21128 27402 21140
rect 27396 21100 27481 21128
rect 27396 21088 27402 21100
rect 26878 21060 26884 21072
rect 25924 21032 26280 21060
rect 26390 21032 26884 21060
rect 25924 21020 25930 21032
rect 26390 20992 26418 21032
rect 26878 21020 26884 21032
rect 26936 21060 26942 21072
rect 26936 21032 27292 21060
rect 26936 21020 26942 21032
rect 27264 21004 27292 21032
rect 25792 20964 26188 20992
rect 24912 20927 24959 20933
rect 24912 20893 24913 20927
rect 24947 20893 24959 20927
rect 24912 20887 24959 20893
rect 25133 20927 25191 20933
rect 25133 20893 25145 20927
rect 25179 20893 25191 20927
rect 25133 20887 25191 20893
rect 24912 20884 24918 20887
rect 25222 20884 25228 20936
rect 25280 20924 25286 20936
rect 25317 20927 25375 20933
rect 25317 20924 25329 20927
rect 25280 20896 25329 20924
rect 25280 20884 25286 20896
rect 25317 20893 25329 20896
rect 25363 20893 25375 20927
rect 25317 20887 25375 20893
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20924 25467 20927
rect 25498 20924 25504 20936
rect 25455 20896 25504 20924
rect 25455 20893 25467 20896
rect 25409 20887 25467 20893
rect 25498 20884 25504 20896
rect 25556 20884 25562 20936
rect 24670 20816 24676 20868
rect 24728 20856 24734 20868
rect 25792 20856 25820 20964
rect 26160 20936 26188 20964
rect 26344 20964 26418 20992
rect 26050 20884 26056 20936
rect 26108 20884 26114 20936
rect 26142 20884 26148 20936
rect 26200 20884 26206 20936
rect 26344 20933 26372 20964
rect 26602 20952 26608 21004
rect 26660 20952 26666 21004
rect 27246 20952 27252 21004
rect 27304 20952 27310 21004
rect 27341 20995 27399 21001
rect 27341 20961 27353 20995
rect 27387 20961 27399 20995
rect 27453 20992 27481 21100
rect 28074 21088 28080 21140
rect 28132 21088 28138 21140
rect 28166 21088 28172 21140
rect 28224 21088 28230 21140
rect 28261 21131 28319 21137
rect 28261 21097 28273 21131
rect 28307 21128 28319 21131
rect 28445 21131 28503 21137
rect 28445 21128 28457 21131
rect 28307 21100 28457 21128
rect 28307 21097 28319 21100
rect 28261 21091 28319 21097
rect 28445 21097 28457 21100
rect 28491 21097 28503 21131
rect 28445 21091 28503 21097
rect 30190 21088 30196 21140
rect 30248 21128 30254 21140
rect 30929 21131 30987 21137
rect 30929 21128 30941 21131
rect 30248 21100 30941 21128
rect 30248 21088 30254 21100
rect 30929 21097 30941 21100
rect 30975 21097 30987 21131
rect 30929 21091 30987 21097
rect 27706 21020 27712 21072
rect 27764 21020 27770 21072
rect 27724 20992 27752 21020
rect 27453 20964 27568 20992
rect 27724 20964 27844 20992
rect 27341 20955 27399 20961
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 26418 20884 26424 20936
rect 26476 20884 26482 20936
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20924 26571 20927
rect 26878 20924 26884 20936
rect 26559 20896 26884 20924
rect 26559 20893 26571 20896
rect 26513 20887 26571 20893
rect 26878 20884 26884 20896
rect 26936 20884 26942 20936
rect 24728 20828 25820 20856
rect 25869 20859 25927 20865
rect 24728 20816 24734 20828
rect 25869 20825 25881 20859
rect 25915 20856 25927 20859
rect 27249 20859 27307 20865
rect 27249 20856 27261 20859
rect 25915 20828 27261 20856
rect 25915 20825 25927 20828
rect 25869 20819 25927 20825
rect 27249 20825 27261 20828
rect 27295 20825 27307 20859
rect 27362 20856 27390 20955
rect 27540 20933 27568 20964
rect 27816 20933 27844 20964
rect 27525 20927 27583 20933
rect 27525 20893 27537 20927
rect 27571 20893 27583 20927
rect 27525 20887 27583 20893
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20893 27859 20927
rect 27801 20887 27859 20893
rect 27985 20927 28043 20933
rect 27985 20893 27997 20927
rect 28031 20893 28043 20927
rect 27985 20887 28043 20893
rect 28077 20927 28135 20933
rect 28077 20893 28089 20927
rect 28123 20893 28135 20927
rect 28184 20924 28212 21088
rect 28353 20927 28411 20933
rect 28353 20924 28365 20927
rect 28184 20896 28365 20924
rect 28077 20887 28135 20893
rect 28353 20893 28365 20896
rect 28399 20893 28411 20927
rect 28353 20887 28411 20893
rect 28000 20856 28028 20887
rect 27362 20828 28028 20856
rect 28092 20856 28120 20887
rect 28626 20884 28632 20936
rect 28684 20884 28690 20936
rect 28721 20927 28779 20933
rect 28721 20893 28733 20927
rect 28767 20924 28779 20927
rect 28810 20924 28816 20936
rect 28767 20896 28816 20924
rect 28767 20893 28779 20896
rect 28721 20887 28779 20893
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 28902 20884 28908 20936
rect 28960 20924 28966 20936
rect 29454 20924 29460 20936
rect 28960 20896 29460 20924
rect 28960 20884 28966 20896
rect 29454 20884 29460 20896
rect 29512 20924 29518 20936
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 29512 20896 29561 20924
rect 29512 20884 29518 20896
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 28644 20856 28672 20884
rect 29794 20859 29852 20865
rect 29794 20856 29806 20859
rect 28092 20828 28672 20856
rect 28920 20828 29806 20856
rect 27249 20819 27307 20825
rect 24544 20760 24624 20788
rect 25041 20791 25099 20797
rect 24544 20748 24550 20760
rect 25041 20757 25053 20791
rect 25087 20788 25099 20791
rect 25498 20788 25504 20800
rect 25087 20760 25504 20788
rect 25087 20757 25099 20760
rect 25041 20751 25099 20757
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 25590 20748 25596 20800
rect 25648 20748 25654 20800
rect 26234 20748 26240 20800
rect 26292 20788 26298 20800
rect 26881 20791 26939 20797
rect 26881 20788 26893 20791
rect 26292 20760 26893 20788
rect 26292 20748 26298 20760
rect 26881 20757 26893 20760
rect 26927 20788 26939 20791
rect 27338 20788 27344 20800
rect 26927 20760 27344 20788
rect 26927 20757 26939 20760
rect 26881 20751 26939 20757
rect 27338 20748 27344 20760
rect 27396 20748 27402 20800
rect 27430 20748 27436 20800
rect 27488 20788 27494 20800
rect 27709 20791 27767 20797
rect 27709 20788 27721 20791
rect 27488 20760 27721 20788
rect 27488 20748 27494 20760
rect 27709 20757 27721 20760
rect 27755 20757 27767 20791
rect 28000 20788 28028 20828
rect 28626 20788 28632 20800
rect 28000 20760 28632 20788
rect 27709 20751 27767 20757
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 28920 20797 28948 20828
rect 29794 20825 29806 20828
rect 29840 20825 29852 20859
rect 29794 20819 29852 20825
rect 28905 20791 28963 20797
rect 28905 20757 28917 20791
rect 28951 20757 28963 20791
rect 28905 20751 28963 20757
rect 1104 20698 43884 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 43884 20698
rect 1104 20624 43884 20646
rect 1673 20587 1731 20593
rect 1673 20553 1685 20587
rect 1719 20584 1731 20587
rect 5258 20584 5264 20596
rect 1719 20556 5264 20584
rect 1719 20553 1731 20556
rect 1673 20547 1731 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 5408 20556 5780 20584
rect 5408 20544 5414 20556
rect 3418 20516 3424 20528
rect 1504 20488 3424 20516
rect 1504 20457 1532 20488
rect 3418 20476 3424 20488
rect 3476 20476 3482 20528
rect 3694 20476 3700 20528
rect 3752 20476 3758 20528
rect 3878 20476 3884 20528
rect 3936 20516 3942 20528
rect 5068 20519 5126 20525
rect 3936 20488 5028 20516
rect 3936 20476 3942 20488
rect 1489 20451 1547 20457
rect 1489 20417 1501 20451
rect 1535 20417 1547 20451
rect 1489 20411 1547 20417
rect 1670 20408 1676 20460
rect 1728 20408 1734 20460
rect 1854 20408 1860 20460
rect 1912 20408 1918 20460
rect 2032 20451 2090 20457
rect 2032 20417 2044 20451
rect 2078 20448 2090 20451
rect 2958 20448 2964 20460
rect 2078 20420 2964 20448
rect 2078 20417 2090 20420
rect 2032 20411 2090 20417
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 3602 20408 3608 20460
rect 3660 20408 3666 20460
rect 4154 20408 4160 20460
rect 4212 20408 4218 20460
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20448 4859 20451
rect 4890 20448 4896 20460
rect 4847 20420 4896 20448
rect 4847 20417 4859 20420
rect 4801 20411 4859 20417
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5000 20448 5028 20488
rect 5068 20485 5080 20519
rect 5114 20516 5126 20519
rect 5626 20516 5632 20528
rect 5114 20488 5632 20516
rect 5114 20485 5126 20488
rect 5068 20479 5126 20485
rect 5626 20476 5632 20488
rect 5684 20476 5690 20528
rect 5752 20516 5780 20556
rect 5810 20544 5816 20596
rect 5868 20584 5874 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 5868 20556 6377 20584
rect 5868 20544 5874 20556
rect 6365 20553 6377 20556
rect 6411 20553 6423 20587
rect 6365 20547 6423 20553
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 7282 20584 7288 20596
rect 6512 20556 6894 20584
rect 6512 20544 6518 20556
rect 6866 20525 6894 20556
rect 7024 20556 7288 20584
rect 6851 20519 6909 20525
rect 5752 20488 5948 20516
rect 5534 20448 5540 20460
rect 5000 20420 5540 20448
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 1872 20380 1900 20408
rect 1811 20352 1900 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 3786 20380 3792 20392
rect 2832 20352 3792 20380
rect 2832 20340 2838 20352
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 3145 20315 3203 20321
rect 3145 20281 3157 20315
rect 3191 20312 3203 20315
rect 4172 20312 4200 20408
rect 5920 20380 5948 20488
rect 6851 20485 6863 20519
rect 6897 20485 6909 20519
rect 6851 20479 6909 20485
rect 6270 20408 6276 20460
rect 6328 20448 6334 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6328 20420 6561 20448
rect 6328 20408 6334 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6178 20380 6184 20392
rect 5920 20352 6184 20380
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 3191 20284 4200 20312
rect 3191 20281 3203 20284
rect 3145 20275 3203 20281
rect 5810 20272 5816 20324
rect 5868 20312 5874 20324
rect 6086 20312 6092 20324
rect 5868 20284 6092 20312
rect 5868 20272 5874 20284
rect 6086 20272 6092 20284
rect 6144 20312 6150 20324
rect 6656 20312 6684 20411
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 7024 20457 7052 20556
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 7926 20544 7932 20596
rect 7984 20544 7990 20596
rect 9030 20544 9036 20596
rect 9088 20584 9094 20596
rect 9088 20556 10180 20584
rect 9088 20544 9094 20556
rect 7960 20516 7988 20544
rect 7852 20488 7988 20516
rect 7009 20451 7067 20457
rect 6788 20420 6833 20448
rect 6788 20408 6794 20420
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 7156 20420 7297 20448
rect 7156 20408 7162 20420
rect 7285 20417 7297 20420
rect 7331 20448 7343 20451
rect 7397 20448 7687 20470
rect 7852 20457 7880 20488
rect 8386 20476 8392 20528
rect 8444 20476 8450 20528
rect 9490 20476 9496 20528
rect 9548 20516 9554 20528
rect 10045 20519 10103 20525
rect 10045 20516 10057 20519
rect 9548 20488 10057 20516
rect 9548 20476 9554 20488
rect 7331 20442 7687 20448
rect 7837 20451 7895 20457
rect 7331 20420 7425 20442
rect 7659 20438 7687 20442
rect 7738 20441 7796 20447
rect 7738 20438 7750 20441
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 7659 20410 7750 20438
rect 7738 20407 7750 20410
rect 7784 20407 7796 20441
rect 7837 20417 7849 20451
rect 7883 20417 7895 20451
rect 7837 20411 7895 20417
rect 7948 20451 8006 20457
rect 7948 20417 7960 20451
rect 7994 20417 8006 20451
rect 7948 20411 8006 20417
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8159 20420 8340 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 7738 20401 7796 20407
rect 7374 20380 7380 20392
rect 7300 20352 7380 20380
rect 7101 20315 7159 20321
rect 7101 20312 7113 20315
rect 6144 20284 7113 20312
rect 6144 20272 6150 20284
rect 7101 20281 7113 20284
rect 7147 20281 7159 20315
rect 7101 20275 7159 20281
rect 7300 20256 7328 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 7485 20312 7513 20343
rect 7558 20340 7564 20392
rect 7616 20340 7622 20392
rect 7960 20312 7988 20411
rect 8202 20340 8208 20392
rect 8260 20340 8266 20392
rect 7485 20284 7988 20312
rect 8312 20312 8340 20420
rect 8478 20408 8484 20460
rect 8536 20408 8542 20460
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 8680 20380 8708 20411
rect 8846 20408 8852 20460
rect 8904 20448 8910 20460
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 8904 20420 9045 20448
rect 8904 20408 8910 20420
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 9125 20451 9183 20457
rect 9125 20417 9137 20451
rect 9171 20448 9183 20451
rect 9306 20448 9312 20460
rect 9171 20420 9312 20448
rect 9171 20417 9183 20420
rect 9125 20411 9183 20417
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 9398 20408 9404 20460
rect 9456 20448 9462 20460
rect 9692 20457 9720 20488
rect 10045 20485 10057 20488
rect 10091 20485 10103 20519
rect 10045 20479 10103 20485
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 9456 20420 9597 20448
rect 9456 20408 9462 20420
rect 9585 20417 9597 20420
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 9766 20408 9772 20460
rect 9824 20408 9830 20460
rect 10152 20457 10180 20556
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10468 20556 10609 20584
rect 10468 20544 10474 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 10597 20547 10655 20553
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 11977 20587 12035 20593
rect 11977 20584 11989 20587
rect 11940 20556 11989 20584
rect 11940 20544 11946 20556
rect 11977 20553 11989 20556
rect 12023 20553 12035 20587
rect 11977 20547 12035 20553
rect 12069 20587 12127 20593
rect 12069 20553 12081 20587
rect 12115 20584 12127 20587
rect 13078 20584 13084 20596
rect 12115 20556 13084 20584
rect 12115 20553 12127 20556
rect 12069 20547 12127 20553
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 13725 20587 13783 20593
rect 13725 20553 13737 20587
rect 13771 20584 13783 20587
rect 14274 20584 14280 20596
rect 13771 20556 14280 20584
rect 13771 20553 13783 20556
rect 13725 20547 13783 20553
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 14553 20587 14611 20593
rect 14553 20553 14565 20587
rect 14599 20584 14611 20587
rect 15102 20584 15108 20596
rect 14599 20556 15108 20584
rect 14599 20553 14611 20556
rect 14553 20547 14611 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 15838 20544 15844 20596
rect 15896 20544 15902 20596
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 16448 20556 17049 20584
rect 16448 20544 16454 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 17037 20547 17095 20553
rect 17678 20544 17684 20596
rect 17736 20584 17742 20596
rect 17736 20556 17908 20584
rect 17736 20544 17742 20556
rect 10502 20476 10508 20528
rect 10560 20476 10566 20528
rect 14912 20519 14970 20525
rect 10704 20488 11560 20516
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20417 10195 20451
rect 10137 20411 10195 20417
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20448 10471 20451
rect 10704 20448 10732 20488
rect 11532 20460 11560 20488
rect 12360 20488 14688 20516
rect 10459 20420 10732 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 8444 20352 8708 20380
rect 8444 20340 8450 20352
rect 9214 20340 9220 20392
rect 9272 20380 9278 20392
rect 9493 20383 9551 20389
rect 9493 20380 9505 20383
rect 9272 20352 9505 20380
rect 9272 20340 9278 20352
rect 9493 20349 9505 20352
rect 9539 20349 9551 20383
rect 9968 20380 9996 20411
rect 10778 20408 10784 20460
rect 10836 20408 10842 20460
rect 10870 20408 10876 20460
rect 10928 20457 10934 20460
rect 10928 20448 10937 20457
rect 11057 20451 11115 20457
rect 10928 20420 10973 20448
rect 10928 20411 10937 20420
rect 11057 20417 11069 20451
rect 11103 20417 11115 20451
rect 11057 20411 11115 20417
rect 10928 20408 10934 20411
rect 10594 20380 10600 20392
rect 9493 20343 9551 20349
rect 9591 20352 10600 20380
rect 8754 20312 8760 20324
rect 8312 20284 8760 20312
rect 3234 20204 3240 20256
rect 3292 20204 3298 20256
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 4709 20247 4767 20253
rect 4709 20244 4721 20247
rect 3660 20216 4721 20244
rect 3660 20204 3666 20216
rect 4709 20213 4721 20216
rect 4755 20244 4767 20247
rect 5166 20244 5172 20256
rect 4755 20216 5172 20244
rect 4755 20213 4767 20216
rect 4709 20207 4767 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 6178 20204 6184 20256
rect 6236 20204 6242 20256
rect 7282 20204 7288 20256
rect 7340 20204 7346 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7485 20244 7513 20284
rect 8754 20272 8760 20284
rect 8812 20312 8818 20324
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8812 20284 9321 20312
rect 8812 20272 8818 20284
rect 9309 20281 9321 20284
rect 9355 20281 9367 20315
rect 9309 20275 9367 20281
rect 7432 20216 7513 20244
rect 7432 20204 7438 20216
rect 8018 20204 8024 20256
rect 8076 20204 8082 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9591 20244 9619 20352
rect 10594 20340 10600 20352
rect 10652 20380 10658 20392
rect 10893 20380 10921 20408
rect 10652 20352 10921 20380
rect 10652 20340 10658 20352
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 11072 20380 11100 20411
rect 11514 20408 11520 20460
rect 11572 20408 11578 20460
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20448 11943 20451
rect 12066 20448 12072 20460
rect 11931 20420 12072 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12360 20457 12388 20488
rect 14660 20460 14688 20488
rect 14912 20485 14924 20519
rect 14958 20516 14970 20519
rect 15010 20516 15016 20528
rect 14958 20488 15016 20516
rect 14958 20485 14970 20488
rect 14912 20479 14970 20485
rect 15010 20476 15016 20488
rect 15068 20476 15074 20528
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12612 20451 12670 20457
rect 12612 20417 12624 20451
rect 12658 20448 12670 20451
rect 12894 20448 12900 20460
rect 12658 20420 12900 20448
rect 12658 20417 12670 20420
rect 12612 20411 12670 20417
rect 11020 20352 11100 20380
rect 11020 20340 11026 20352
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 12158 20380 12164 20392
rect 11204 20352 12164 20380
rect 11204 20340 11210 20352
rect 12158 20340 12164 20352
rect 12216 20380 12222 20392
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 12216 20352 12265 20380
rect 12216 20340 12222 20352
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 9766 20272 9772 20324
rect 9824 20312 9830 20324
rect 12360 20312 12388 20411
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 14274 20448 14280 20460
rect 13863 20420 14280 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 14642 20408 14648 20460
rect 14700 20408 14706 20460
rect 15856 20448 15884 20544
rect 16316 20488 17264 20516
rect 14752 20420 15884 20448
rect 14182 20340 14188 20392
rect 14240 20380 14246 20392
rect 14752 20380 14780 20420
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16206 20448 16212 20460
rect 16080 20420 16212 20448
rect 16080 20408 16086 20420
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16316 20457 16344 20488
rect 17236 20460 17264 20488
rect 17586 20476 17592 20528
rect 17644 20516 17650 20528
rect 17880 20516 17908 20556
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18138 20584 18144 20596
rect 18012 20556 18144 20584
rect 18012 20544 18018 20556
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18414 20544 18420 20596
rect 18472 20544 18478 20596
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 19153 20587 19211 20593
rect 19153 20584 19165 20587
rect 18932 20556 19165 20584
rect 18932 20544 18938 20556
rect 19153 20553 19165 20556
rect 19199 20553 19211 20587
rect 19153 20547 19211 20553
rect 19521 20587 19579 20593
rect 19521 20553 19533 20587
rect 19567 20584 19579 20587
rect 21266 20584 21272 20596
rect 19567 20556 21272 20584
rect 19567 20553 19579 20556
rect 19521 20547 19579 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 21692 20556 22201 20584
rect 21692 20544 21698 20556
rect 22189 20553 22201 20556
rect 22235 20584 22247 20587
rect 22235 20556 22692 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 19889 20519 19947 20525
rect 17644 20488 17816 20516
rect 17644 20476 17650 20488
rect 17788 20460 17816 20488
rect 17880 20488 19288 20516
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 16485 20451 16543 20457
rect 16485 20417 16497 20451
rect 16531 20448 16543 20451
rect 16669 20451 16727 20457
rect 16531 20420 16620 20448
rect 16531 20417 16543 20420
rect 16485 20411 16543 20417
rect 14240 20352 14780 20380
rect 14240 20340 14246 20352
rect 9824 20284 12388 20312
rect 16592 20312 16620 20420
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17126 20448 17132 20460
rect 16715 20420 17132 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17310 20408 17316 20460
rect 17368 20408 17374 20460
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 16761 20383 16819 20389
rect 16761 20349 16773 20383
rect 16807 20380 16819 20383
rect 16850 20380 16856 20392
rect 16807 20352 16856 20380
rect 16807 20349 16819 20352
rect 16761 20343 16819 20349
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 17328 20380 17356 20408
rect 16960 20352 17356 20380
rect 17512 20380 17540 20411
rect 17770 20408 17776 20460
rect 17828 20408 17834 20460
rect 17880 20457 17908 20488
rect 19260 20460 19288 20488
rect 19352 20488 19656 20516
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 18138 20408 18144 20460
rect 18196 20448 18202 20460
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 18196 20420 18245 20448
rect 18196 20408 18202 20420
rect 18233 20417 18245 20420
rect 18279 20448 18291 20451
rect 18322 20448 18328 20460
rect 18279 20420 18328 20448
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 18785 20451 18843 20457
rect 18785 20448 18797 20451
rect 18472 20420 18797 20448
rect 18472 20408 18478 20420
rect 18785 20417 18797 20420
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19352 20457 19380 20488
rect 19628 20460 19656 20488
rect 19889 20485 19901 20519
rect 19935 20516 19947 20519
rect 19978 20516 19984 20528
rect 19935 20488 19984 20516
rect 19935 20485 19947 20488
rect 19889 20479 19947 20485
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 20165 20519 20223 20525
rect 20165 20485 20177 20519
rect 20211 20516 20223 20519
rect 21082 20516 21088 20528
rect 20211 20488 21088 20516
rect 20211 20485 20223 20488
rect 20165 20479 20223 20485
rect 21082 20476 21088 20488
rect 21140 20516 21146 20528
rect 22002 20516 22008 20528
rect 21140 20488 22008 20516
rect 21140 20476 21146 20488
rect 22002 20476 22008 20488
rect 22060 20476 22066 20528
rect 22462 20476 22468 20528
rect 22520 20476 22526 20528
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20417 19395 20451
rect 19337 20411 19395 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 19426 20380 19432 20392
rect 17512 20352 19432 20380
rect 16960 20312 16988 20352
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 19536 20380 19564 20411
rect 19610 20408 19616 20460
rect 19668 20408 19674 20460
rect 19702 20408 19708 20460
rect 19760 20448 19766 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19760 20420 20085 20448
rect 19760 20408 19766 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20530 20448 20536 20460
rect 20303 20420 20536 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20448 20683 20451
rect 22480 20448 22508 20476
rect 22664 20457 22692 20556
rect 24486 20544 24492 20596
rect 24544 20544 24550 20596
rect 25406 20584 25412 20596
rect 24928 20556 25412 20584
rect 22848 20488 24256 20516
rect 22848 20457 22876 20488
rect 24228 20460 24256 20488
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 20671 20420 21128 20448
rect 22480 20420 22569 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 21100 20392 21128 20420
rect 22557 20417 22569 20420
rect 22603 20417 22615 20451
rect 22557 20411 22615 20417
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 22922 20408 22928 20460
rect 22980 20408 22986 20460
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 23569 20451 23627 20457
rect 23569 20448 23581 20451
rect 23532 20420 23581 20448
rect 23532 20408 23538 20420
rect 23569 20417 23581 20420
rect 23615 20448 23627 20451
rect 24118 20448 24124 20460
rect 23615 20420 24124 20448
rect 23615 20417 23627 20420
rect 23569 20411 23627 20417
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24210 20408 24216 20460
rect 24268 20408 24274 20460
rect 19794 20380 19800 20392
rect 19536 20352 19800 20380
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 19886 20340 19892 20392
rect 19944 20380 19950 20392
rect 20806 20380 20812 20392
rect 19944 20352 20812 20380
rect 19944 20340 19950 20352
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 21082 20340 21088 20392
rect 21140 20340 21146 20392
rect 22940 20380 22968 20408
rect 23385 20383 23443 20389
rect 23385 20380 23397 20383
rect 22940 20352 23397 20380
rect 23385 20349 23397 20352
rect 23431 20349 23443 20383
rect 23385 20343 23443 20349
rect 24026 20340 24032 20392
rect 24084 20380 24090 20392
rect 24394 20380 24400 20392
rect 24084 20352 24400 20380
rect 24084 20340 24090 20352
rect 24394 20340 24400 20352
rect 24452 20340 24458 20392
rect 16592 20284 16988 20312
rect 9824 20272 9830 20284
rect 17034 20272 17040 20324
rect 17092 20312 17098 20324
rect 20346 20312 20352 20324
rect 17092 20284 20352 20312
rect 17092 20272 17098 20284
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 24504 20312 24532 20544
rect 24578 20476 24584 20528
rect 24636 20476 24642 20528
rect 24596 20380 24624 20476
rect 24762 20408 24768 20460
rect 24820 20408 24826 20460
rect 24928 20457 24956 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25590 20544 25596 20596
rect 25648 20584 25654 20596
rect 26697 20587 26755 20593
rect 25648 20556 26285 20584
rect 25648 20544 25654 20556
rect 25133 20519 25191 20525
rect 25133 20485 25145 20519
rect 25179 20516 25191 20519
rect 25958 20516 25964 20528
rect 25179 20488 25964 20516
rect 25179 20485 25191 20488
rect 25133 20479 25191 20485
rect 25958 20476 25964 20488
rect 26016 20476 26022 20528
rect 26257 20516 26285 20556
rect 26697 20553 26709 20587
rect 26743 20584 26755 20587
rect 26970 20584 26976 20596
rect 26743 20556 26976 20584
rect 26743 20553 26755 20556
rect 26697 20547 26755 20553
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 28258 20584 28264 20596
rect 27081 20556 28264 20584
rect 27081 20516 27109 20556
rect 28258 20544 28264 20556
rect 28316 20584 28322 20596
rect 28629 20587 28687 20593
rect 28629 20584 28641 20587
rect 28316 20556 28641 20584
rect 28316 20544 28322 20556
rect 28629 20553 28641 20556
rect 28675 20553 28687 20587
rect 28629 20547 28687 20553
rect 26257 20488 26372 20516
rect 24913 20451 24971 20457
rect 24913 20417 24925 20451
rect 24959 20417 24971 20451
rect 24913 20411 24971 20417
rect 25041 20451 25099 20457
rect 25041 20417 25053 20451
rect 25087 20417 25099 20451
rect 25041 20411 25099 20417
rect 25230 20451 25288 20457
rect 25230 20417 25242 20451
rect 25276 20417 25288 20451
rect 25230 20411 25288 20417
rect 25056 20380 25084 20411
rect 24596 20352 25084 20380
rect 24780 20324 24808 20352
rect 20916 20284 24532 20312
rect 8352 20216 9619 20244
rect 8352 20204 8358 20216
rect 10226 20204 10232 20256
rect 10284 20244 10290 20256
rect 10505 20247 10563 20253
rect 10505 20244 10517 20247
rect 10284 20216 10517 20244
rect 10284 20204 10290 20216
rect 10505 20213 10517 20216
rect 10551 20213 10563 20247
rect 10505 20207 10563 20213
rect 10870 20204 10876 20256
rect 10928 20244 10934 20256
rect 10965 20247 11023 20253
rect 10965 20244 10977 20247
rect 10928 20216 10977 20244
rect 10928 20204 10934 20216
rect 10965 20213 10977 20216
rect 11011 20213 11023 20247
rect 10965 20207 11023 20213
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11793 20247 11851 20253
rect 11793 20244 11805 20247
rect 11204 20216 11805 20244
rect 11204 20204 11210 20216
rect 11793 20213 11805 20216
rect 11839 20244 11851 20247
rect 12066 20244 12072 20256
rect 11839 20216 12072 20244
rect 11839 20213 11851 20216
rect 11793 20207 11851 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 12161 20247 12219 20253
rect 12161 20213 12173 20247
rect 12207 20244 12219 20247
rect 12526 20244 12532 20256
rect 12207 20216 12532 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13814 20244 13820 20256
rect 13320 20216 13820 20244
rect 13320 20204 13326 20216
rect 13814 20204 13820 20216
rect 13872 20244 13878 20256
rect 14001 20247 14059 20253
rect 14001 20244 14013 20247
rect 13872 20216 14013 20244
rect 13872 20204 13878 20216
rect 14001 20213 14013 20216
rect 14047 20213 14059 20247
rect 14001 20207 14059 20213
rect 16301 20247 16359 20253
rect 16301 20213 16313 20247
rect 16347 20244 16359 20247
rect 16390 20244 16396 20256
rect 16347 20216 16396 20244
rect 16347 20213 16359 20216
rect 16301 20207 16359 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16853 20247 16911 20253
rect 16853 20213 16865 20247
rect 16899 20244 16911 20247
rect 17494 20244 17500 20256
rect 16899 20216 17500 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 17586 20204 17592 20256
rect 17644 20244 17650 20256
rect 20916 20244 20944 20284
rect 24762 20272 24768 20324
rect 24820 20272 24826 20324
rect 17644 20216 20944 20244
rect 17644 20204 17650 20216
rect 21082 20204 21088 20256
rect 21140 20244 21146 20256
rect 21177 20247 21235 20253
rect 21177 20244 21189 20247
rect 21140 20216 21189 20244
rect 21140 20204 21146 20216
rect 21177 20213 21189 20216
rect 21223 20244 21235 20247
rect 21545 20247 21603 20253
rect 21545 20244 21557 20247
rect 21223 20216 21557 20244
rect 21223 20213 21235 20216
rect 21177 20207 21235 20213
rect 21545 20213 21557 20216
rect 21591 20244 21603 20247
rect 22186 20244 22192 20256
rect 21591 20216 22192 20244
rect 21591 20213 21603 20216
rect 21545 20207 21603 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 22373 20247 22431 20253
rect 22373 20213 22385 20247
rect 22419 20244 22431 20247
rect 23290 20244 23296 20256
rect 22419 20216 23296 20244
rect 22419 20213 22431 20216
rect 22373 20207 22431 20213
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 23569 20247 23627 20253
rect 23569 20213 23581 20247
rect 23615 20244 23627 20247
rect 23658 20244 23664 20256
rect 23615 20216 23664 20244
rect 23615 20213 23627 20216
rect 23569 20207 23627 20213
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 23750 20204 23756 20256
rect 23808 20204 23814 20256
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24946 20244 24952 20256
rect 24360 20216 24952 20244
rect 24360 20204 24366 20216
rect 24946 20204 24952 20216
rect 25004 20244 25010 20256
rect 25245 20244 25273 20411
rect 25774 20408 25780 20460
rect 25832 20408 25838 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26234 20448 26240 20460
rect 26099 20420 26240 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 26344 20457 26372 20488
rect 26988 20488 27109 20516
rect 27157 20519 27215 20525
rect 26329 20451 26387 20457
rect 26329 20417 26341 20451
rect 26375 20417 26387 20451
rect 26329 20411 26387 20417
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 25869 20383 25927 20389
rect 25869 20380 25881 20383
rect 25556 20352 25881 20380
rect 25556 20340 25562 20352
rect 25869 20349 25881 20352
rect 25915 20349 25927 20383
rect 26418 20380 26424 20392
rect 25869 20343 25927 20349
rect 25976 20352 26424 20380
rect 25976 20312 26004 20352
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 25332 20284 26004 20312
rect 25332 20256 25360 20284
rect 26234 20272 26240 20324
rect 26292 20272 26298 20324
rect 26988 20312 27016 20488
rect 27157 20485 27169 20519
rect 27203 20516 27215 20519
rect 27890 20516 27896 20528
rect 27203 20488 27896 20516
rect 27203 20485 27215 20488
rect 27157 20479 27215 20485
rect 27890 20476 27896 20488
rect 27948 20476 27954 20528
rect 28000 20488 29132 20516
rect 27062 20408 27068 20460
rect 27120 20408 27126 20460
rect 27338 20408 27344 20460
rect 27396 20448 27402 20460
rect 28000 20457 28028 20488
rect 29104 20460 29132 20488
rect 27433 20451 27491 20457
rect 27433 20448 27445 20451
rect 27396 20420 27445 20448
rect 27396 20408 27402 20420
rect 27433 20417 27445 20420
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 27709 20451 27767 20457
rect 27709 20417 27721 20451
rect 27755 20417 27767 20451
rect 27709 20411 27767 20417
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 27080 20380 27108 20408
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 27080 20352 27261 20380
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27724 20380 27752 20411
rect 28258 20408 28264 20460
rect 28316 20408 28322 20460
rect 28442 20408 28448 20460
rect 28500 20408 28506 20460
rect 28534 20408 28540 20460
rect 28592 20408 28598 20460
rect 29086 20408 29092 20460
rect 29144 20408 29150 20460
rect 27249 20343 27307 20349
rect 27448 20352 27752 20380
rect 27448 20324 27476 20352
rect 27798 20340 27804 20392
rect 27856 20340 27862 20392
rect 28166 20340 28172 20392
rect 28224 20340 28230 20392
rect 26988 20284 27200 20312
rect 25004 20216 25273 20244
rect 25004 20204 25010 20216
rect 25314 20204 25320 20256
rect 25372 20204 25378 20256
rect 25406 20204 25412 20256
rect 25464 20204 25470 20256
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 25777 20247 25835 20253
rect 25777 20244 25789 20247
rect 25740 20216 25789 20244
rect 25740 20204 25746 20216
rect 25777 20213 25789 20216
rect 25823 20213 25835 20247
rect 25777 20207 25835 20213
rect 26513 20247 26571 20253
rect 26513 20213 26525 20247
rect 26559 20244 26571 20247
rect 26786 20244 26792 20256
rect 26559 20216 26792 20244
rect 26559 20213 26571 20216
rect 26513 20207 26571 20213
rect 26786 20204 26792 20216
rect 26844 20204 26850 20256
rect 27172 20253 27200 20284
rect 27338 20272 27344 20324
rect 27396 20272 27402 20324
rect 27430 20272 27436 20324
rect 27488 20272 27494 20324
rect 27617 20315 27675 20321
rect 27617 20281 27629 20315
rect 27663 20312 27675 20315
rect 28184 20312 28212 20340
rect 28552 20312 28580 20408
rect 27663 20284 28212 20312
rect 28276 20284 28580 20312
rect 27663 20281 27675 20284
rect 27617 20275 27675 20281
rect 27157 20247 27215 20253
rect 27157 20213 27169 20247
rect 27203 20213 27215 20247
rect 27356 20244 27384 20272
rect 27798 20244 27804 20256
rect 27356 20216 27804 20244
rect 27157 20207 27215 20213
rect 27798 20204 27804 20216
rect 27856 20204 27862 20256
rect 27985 20247 28043 20253
rect 27985 20213 27997 20247
rect 28031 20244 28043 20247
rect 28074 20244 28080 20256
rect 28031 20216 28080 20244
rect 28031 20213 28043 20216
rect 27985 20207 28043 20213
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 28166 20204 28172 20256
rect 28224 20244 28230 20256
rect 28276 20244 28304 20284
rect 28224 20216 28304 20244
rect 28353 20247 28411 20253
rect 28224 20204 28230 20216
rect 28353 20213 28365 20247
rect 28399 20244 28411 20247
rect 28442 20244 28448 20256
rect 28399 20216 28448 20244
rect 28399 20213 28411 20216
rect 28353 20207 28411 20213
rect 28442 20204 28448 20216
rect 28500 20204 28506 20256
rect 1104 20154 43884 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 43884 20154
rect 1104 20080 43884 20102
rect 2958 20000 2964 20052
rect 3016 20040 3022 20052
rect 3605 20043 3663 20049
rect 3016 20012 3556 20040
rect 3016 20000 3022 20012
rect 3528 19972 3556 20012
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 3786 20040 3792 20052
rect 3651 20012 3792 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 3786 20000 3792 20012
rect 3844 20040 3850 20052
rect 4890 20040 4896 20052
rect 3844 20012 4896 20040
rect 3844 20000 3850 20012
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 5040 20012 5365 20040
rect 5040 20000 5046 20012
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 5994 20040 6000 20052
rect 5684 20012 6000 20040
rect 5684 20000 5690 20012
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6454 20000 6460 20052
rect 6512 20040 6518 20052
rect 8018 20040 8024 20052
rect 6512 20012 8024 20040
rect 6512 20000 6518 20012
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 9030 20000 9036 20052
rect 9088 20040 9094 20052
rect 9585 20043 9643 20049
rect 9585 20040 9597 20043
rect 9088 20012 9597 20040
rect 9088 20000 9094 20012
rect 9585 20009 9597 20012
rect 9631 20009 9643 20043
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 9585 20003 9643 20009
rect 10980 20012 11897 20040
rect 10980 19984 11008 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 12952 20012 13277 20040
rect 12952 20000 12958 20012
rect 13265 20009 13277 20012
rect 13311 20009 13323 20043
rect 13265 20003 13323 20009
rect 13909 20043 13967 20049
rect 13909 20009 13921 20043
rect 13955 20040 13967 20043
rect 15194 20040 15200 20052
rect 13955 20012 15200 20040
rect 13955 20009 13967 20012
rect 13909 20003 13967 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 17678 20000 17684 20052
rect 17736 20040 17742 20052
rect 18598 20040 18604 20052
rect 17736 20012 18604 20040
rect 17736 20000 17742 20012
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19150 20040 19156 20052
rect 18739 20012 19156 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 21082 20000 21088 20052
rect 21140 20040 21146 20052
rect 21453 20043 21511 20049
rect 21453 20040 21465 20043
rect 21140 20012 21465 20040
rect 21140 20000 21146 20012
rect 21453 20009 21465 20012
rect 21499 20009 21511 20043
rect 21453 20003 21511 20009
rect 21634 20000 21640 20052
rect 21692 20040 21698 20052
rect 22097 20043 22155 20049
rect 22097 20040 22109 20043
rect 21692 20012 22109 20040
rect 21692 20000 21698 20012
rect 22097 20009 22109 20012
rect 22143 20040 22155 20043
rect 22738 20040 22744 20052
rect 22143 20012 22744 20040
rect 22143 20009 22155 20012
rect 22097 20003 22155 20009
rect 22738 20000 22744 20012
rect 22796 20000 22802 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 24762 20040 24768 20052
rect 24176 20012 24768 20040
rect 24176 20000 24182 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 25406 20000 25412 20052
rect 25464 20000 25470 20052
rect 25774 20000 25780 20052
rect 25832 20000 25838 20052
rect 26418 20000 26424 20052
rect 26476 20040 26482 20052
rect 26881 20043 26939 20049
rect 26881 20040 26893 20043
rect 26476 20012 26893 20040
rect 26476 20000 26482 20012
rect 26881 20009 26893 20012
rect 26927 20009 26939 20043
rect 27522 20040 27528 20052
rect 26881 20003 26939 20009
rect 27172 20012 27528 20040
rect 5813 19975 5871 19981
rect 5813 19972 5825 19975
rect 3528 19944 5825 19972
rect 5813 19941 5825 19944
rect 5859 19941 5871 19975
rect 5813 19935 5871 19941
rect 6365 19975 6423 19981
rect 6365 19941 6377 19975
rect 6411 19972 6423 19975
rect 7282 19972 7288 19984
rect 6411 19944 7288 19972
rect 6411 19941 6423 19944
rect 6365 19935 6423 19941
rect 7282 19932 7288 19944
rect 7340 19932 7346 19984
rect 8757 19975 8815 19981
rect 8757 19941 8769 19975
rect 8803 19972 8815 19975
rect 8803 19944 9076 19972
rect 8803 19941 8815 19944
rect 8757 19935 8815 19941
rect 1210 19864 1216 19916
rect 1268 19904 1274 19916
rect 1857 19907 1915 19913
rect 1857 19904 1869 19907
rect 1268 19876 1869 19904
rect 1268 19864 1274 19876
rect 1857 19873 1869 19876
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 3050 19864 3056 19916
rect 3108 19864 3114 19916
rect 3234 19864 3240 19916
rect 3292 19904 3298 19916
rect 9048 19913 9076 19944
rect 10962 19932 10968 19984
rect 11020 19932 11026 19984
rect 11149 19975 11207 19981
rect 11149 19941 11161 19975
rect 11195 19972 11207 19975
rect 11195 19944 11284 19972
rect 11195 19941 11207 19944
rect 11149 19935 11207 19941
rect 11256 19916 11284 19944
rect 11974 19932 11980 19984
rect 12032 19972 12038 19984
rect 12032 19944 12480 19972
rect 12032 19932 12038 19944
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3292 19876 4077 19904
rect 3292 19864 3298 19876
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 9033 19907 9091 19913
rect 4755 19876 5672 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19836 1639 19839
rect 3694 19836 3700 19848
rect 1627 19808 3700 19836
rect 1627 19805 1639 19808
rect 1581 19799 1639 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 4798 19796 4804 19848
rect 4856 19796 4862 19848
rect 4982 19796 4988 19848
rect 5040 19796 5046 19848
rect 5074 19796 5080 19848
rect 5132 19796 5138 19848
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 5184 19768 5212 19799
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5644 19845 5672 19876
rect 9033 19873 9045 19907
rect 9079 19904 9091 19907
rect 9122 19904 9128 19916
rect 9079 19876 9128 19904
rect 9079 19873 9091 19876
rect 9033 19867 9091 19873
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 9766 19864 9772 19916
rect 9824 19864 9830 19916
rect 11238 19864 11244 19916
rect 11296 19864 11302 19916
rect 11698 19864 11704 19916
rect 11756 19904 11762 19916
rect 11882 19904 11888 19916
rect 11756 19876 11888 19904
rect 11756 19864 11762 19876
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12342 19864 12348 19916
rect 12400 19864 12406 19916
rect 12452 19904 12480 19944
rect 12986 19932 12992 19984
rect 13044 19972 13050 19984
rect 14185 19975 14243 19981
rect 14185 19972 14197 19975
rect 13044 19944 14197 19972
rect 13044 19932 13050 19944
rect 14185 19941 14197 19944
rect 14231 19941 14243 19975
rect 14185 19935 14243 19941
rect 16206 19932 16212 19984
rect 16264 19932 16270 19984
rect 16758 19972 16764 19984
rect 16316 19944 16764 19972
rect 12452 19876 13032 19904
rect 5445 19839 5503 19845
rect 5445 19836 5457 19839
rect 5316 19808 5457 19836
rect 5316 19796 5322 19808
rect 5445 19805 5457 19808
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 5629 19839 5687 19845
rect 5629 19805 5641 19839
rect 5675 19805 5687 19839
rect 5629 19799 5687 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19836 6331 19839
rect 6362 19836 6368 19848
rect 6319 19808 6368 19836
rect 6319 19805 6331 19808
rect 6273 19799 6331 19805
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 7073 19839 7131 19845
rect 6779 19808 6960 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6181 19771 6239 19777
rect 6181 19768 6193 19771
rect 4028 19740 6193 19768
rect 4028 19728 4034 19740
rect 6181 19737 6193 19740
rect 6227 19768 6239 19771
rect 6822 19768 6828 19780
rect 6227 19740 6828 19768
rect 6227 19737 6239 19740
rect 6181 19731 6239 19737
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 6932 19700 6960 19808
rect 7073 19805 7085 19839
rect 7119 19836 7131 19839
rect 7119 19808 7200 19836
rect 7119 19805 7131 19808
rect 7073 19799 7131 19805
rect 7172 19768 7200 19808
rect 7282 19796 7288 19848
rect 7340 19796 7346 19848
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 7466 19836 7472 19848
rect 7423 19808 7472 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 8202 19836 8208 19848
rect 7576 19808 8208 19836
rect 7576 19768 7604 19808
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 10410 19836 10416 19848
rect 9732 19808 10416 19836
rect 9732 19796 9738 19808
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10778 19796 10784 19848
rect 10836 19796 10842 19848
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11572 19808 12173 19836
rect 11572 19796 11578 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 12437 19839 12495 19845
rect 12299 19808 12388 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 7172 19740 7604 19768
rect 7644 19771 7702 19777
rect 7644 19737 7656 19771
rect 7690 19768 7702 19771
rect 8478 19768 8484 19780
rect 7690 19740 8484 19768
rect 7690 19737 7702 19740
rect 7644 19731 7702 19737
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 8846 19728 8852 19780
rect 8904 19768 8910 19780
rect 9692 19768 9720 19796
rect 8904 19740 9720 19768
rect 10036 19771 10094 19777
rect 8904 19728 8910 19740
rect 10036 19737 10048 19771
rect 10082 19768 10094 19771
rect 10686 19768 10692 19780
rect 10082 19740 10692 19768
rect 10082 19737 10094 19740
rect 10036 19731 10094 19737
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 10796 19768 10824 19796
rect 12360 19780 12388 19808
rect 12437 19805 12449 19839
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 10796 19740 12296 19768
rect 8386 19700 8392 19712
rect 5316 19672 8392 19700
rect 5316 19660 5322 19672
rect 8386 19660 8392 19672
rect 8444 19700 8450 19712
rect 10134 19700 10140 19712
rect 8444 19672 10140 19700
rect 8444 19660 8450 19672
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 10318 19660 10324 19712
rect 10376 19700 10382 19712
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 10376 19672 11989 19700
rect 10376 19660 10382 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 12268 19700 12296 19740
rect 12342 19728 12348 19780
rect 12400 19728 12406 19780
rect 12452 19700 12480 19799
rect 12618 19796 12624 19848
rect 12676 19796 12682 19848
rect 13004 19780 13032 19876
rect 13538 19864 13544 19916
rect 13596 19904 13602 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 13596 19876 14381 19904
rect 13596 19864 13602 19876
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 14476 19876 15332 19904
rect 13078 19796 13084 19848
rect 13136 19836 13142 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13136 19808 14105 19836
rect 13136 19796 13142 19808
rect 14093 19805 14105 19808
rect 14139 19836 14151 19839
rect 14476 19836 14504 19876
rect 15304 19848 15332 19876
rect 16022 19864 16028 19916
rect 16080 19864 16086 19916
rect 14139 19808 14504 19836
rect 14553 19839 14611 19845
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 12986 19728 12992 19780
rect 13044 19768 13050 19780
rect 14458 19768 14464 19780
rect 13044 19740 14464 19768
rect 13044 19728 13050 19740
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 12268 19672 12480 19700
rect 11977 19663 12035 19669
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 13078 19700 13084 19712
rect 12860 19672 13084 19700
rect 12860 19660 12866 19672
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14568 19700 14596 19799
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14826 19836 14832 19848
rect 14700 19808 14832 19836
rect 14700 19796 14706 19808
rect 14826 19796 14832 19808
rect 14884 19836 14890 19848
rect 14921 19839 14979 19845
rect 14921 19836 14933 19839
rect 14884 19808 14933 19836
rect 14884 19796 14890 19808
rect 14921 19805 14933 19808
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15102 19796 15108 19848
rect 15160 19796 15166 19848
rect 15286 19796 15292 19848
rect 15344 19796 15350 19848
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 16316 19845 16344 19944
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 16850 19932 16856 19984
rect 16908 19972 16914 19984
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 16908 19944 17601 19972
rect 16908 19932 16914 19944
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 17589 19935 17647 19941
rect 18966 19932 18972 19984
rect 19024 19972 19030 19984
rect 19024 19944 19840 19972
rect 19024 19932 19030 19944
rect 18141 19907 18199 19913
rect 18141 19904 18153 19907
rect 16408 19876 18153 19904
rect 16301 19839 16359 19845
rect 15436 19808 16160 19836
rect 15436 19796 15442 19808
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15654 19768 15660 19780
rect 15243 19740 15660 19768
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 16132 19768 16160 19808
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16408 19768 16436 19876
rect 18141 19873 18153 19876
rect 18187 19904 18199 19907
rect 18598 19904 18604 19916
rect 18187 19876 18604 19904
rect 18187 19873 18199 19876
rect 18141 19867 18199 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 16132 19740 16436 19768
rect 14240 19672 14596 19700
rect 14240 19660 14246 19672
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 16500 19700 16528 19799
rect 16758 19796 16764 19848
rect 16816 19796 16822 19848
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17586 19836 17592 19848
rect 17092 19808 17592 19836
rect 17092 19796 17098 19808
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17770 19796 17776 19848
rect 17828 19796 17834 19848
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 17310 19728 17316 19780
rect 17368 19768 17374 19780
rect 17880 19768 17908 19799
rect 17368 19740 17908 19768
rect 18248 19768 18276 19799
rect 18322 19796 18328 19848
rect 18380 19836 18386 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18380 19808 18705 19836
rect 18380 19796 18386 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18840 19808 18889 19836
rect 18840 19796 18846 19808
rect 18877 19805 18889 19808
rect 18923 19836 18935 19839
rect 19076 19836 19104 19944
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 19392 19876 19717 19904
rect 19392 19864 19398 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 19812 19904 19840 19944
rect 20162 19932 20168 19984
rect 20220 19972 20226 19984
rect 21726 19972 21732 19984
rect 20220 19944 21732 19972
rect 20220 19932 20226 19944
rect 21726 19932 21732 19944
rect 21784 19932 21790 19984
rect 22186 19932 22192 19984
rect 22244 19972 22250 19984
rect 22462 19972 22468 19984
rect 22244 19944 22468 19972
rect 22244 19932 22250 19944
rect 22462 19932 22468 19944
rect 22520 19972 22526 19984
rect 24026 19972 24032 19984
rect 22520 19944 24032 19972
rect 22520 19932 22526 19944
rect 24026 19932 24032 19944
rect 24084 19932 24090 19984
rect 24210 19932 24216 19984
rect 24268 19972 24274 19984
rect 24854 19972 24860 19984
rect 24268 19944 24860 19972
rect 24268 19932 24274 19944
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 25130 19932 25136 19984
rect 25188 19932 25194 19984
rect 25332 19944 27108 19972
rect 19812 19876 20576 19904
rect 19705 19867 19763 19873
rect 20548 19848 20576 19876
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 20717 19907 20775 19913
rect 20717 19904 20729 19907
rect 20680 19876 20729 19904
rect 20680 19864 20686 19876
rect 20717 19873 20729 19876
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 22094 19904 22100 19916
rect 20864 19876 22100 19904
rect 20864 19864 20870 19876
rect 22094 19864 22100 19876
rect 22152 19864 22158 19916
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 23842 19904 23848 19916
rect 23348 19876 23848 19904
rect 23348 19864 23354 19876
rect 23842 19864 23848 19876
rect 23900 19904 23906 19916
rect 25148 19904 25176 19932
rect 23900 19876 24716 19904
rect 23900 19864 23906 19876
rect 18923 19808 19104 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19150 19796 19156 19848
rect 19208 19796 19214 19848
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19168 19768 19196 19796
rect 18248 19740 19196 19768
rect 19444 19768 19472 19799
rect 19518 19796 19524 19848
rect 19576 19796 19582 19848
rect 19966 19845 20015 19846
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 19935 19839 20015 19845
rect 19935 19805 19947 19839
rect 19981 19836 20015 19839
rect 20070 19836 20076 19848
rect 19981 19808 20076 19836
rect 19981 19805 19993 19808
rect 19935 19799 19993 19805
rect 19812 19768 19840 19799
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20441 19799 20499 19805
rect 19444 19740 19840 19768
rect 17368 19728 17374 19740
rect 15068 19672 16528 19700
rect 17880 19700 17908 19740
rect 19536 19712 19564 19740
rect 20346 19728 20352 19780
rect 20404 19768 20410 19780
rect 20456 19768 20484 19799
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20404 19740 20484 19768
rect 20404 19728 20410 19740
rect 18230 19700 18236 19712
rect 17880 19672 18236 19700
rect 15068 19660 15074 19672
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18874 19700 18880 19712
rect 18472 19672 18880 19700
rect 18472 19660 18478 19672
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 19518 19660 19524 19712
rect 19576 19660 19582 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20640 19700 20668 19864
rect 24688 19848 24716 19876
rect 25056 19876 25176 19904
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 20956 19808 21312 19836
rect 20956 19796 20962 19808
rect 21284 19768 21312 19808
rect 21450 19796 21456 19848
rect 21508 19796 21514 19848
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19836 21695 19839
rect 21910 19836 21916 19848
rect 21683 19808 21916 19836
rect 21683 19805 21695 19808
rect 21637 19799 21695 19805
rect 21910 19796 21916 19808
rect 21968 19796 21974 19848
rect 24394 19836 24400 19848
rect 22066 19808 24400 19836
rect 22066 19768 22094 19808
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 24578 19796 24584 19848
rect 24636 19796 24642 19848
rect 24670 19796 24676 19848
rect 24728 19836 24734 19848
rect 24946 19836 24952 19848
rect 24728 19808 24952 19836
rect 24728 19796 24734 19808
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 21284 19740 22094 19768
rect 22281 19771 22339 19777
rect 22281 19737 22293 19771
rect 22327 19737 22339 19771
rect 22281 19731 22339 19737
rect 20036 19672 20668 19700
rect 20036 19660 20042 19672
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21821 19703 21879 19709
rect 21821 19700 21833 19703
rect 21324 19672 21833 19700
rect 21324 19660 21330 19672
rect 21821 19669 21833 19672
rect 21867 19669 21879 19703
rect 21821 19663 21879 19669
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 22296 19700 22324 19731
rect 22738 19728 22744 19780
rect 22796 19768 22802 19780
rect 23017 19771 23075 19777
rect 23017 19768 23029 19771
rect 22796 19740 23029 19768
rect 22796 19728 22802 19740
rect 23017 19737 23029 19740
rect 23063 19768 23075 19771
rect 24302 19768 24308 19780
rect 23063 19740 24308 19768
rect 23063 19737 23075 19740
rect 23017 19731 23075 19737
rect 24302 19728 24308 19740
rect 24360 19728 24366 19780
rect 24762 19728 24768 19780
rect 24820 19728 24826 19780
rect 24857 19771 24915 19777
rect 24857 19737 24869 19771
rect 24903 19768 24915 19771
rect 25056 19768 25084 19876
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 25332 19845 25360 19944
rect 25406 19864 25412 19916
rect 25464 19864 25470 19916
rect 26142 19864 26148 19916
rect 26200 19904 26206 19916
rect 26200 19876 26280 19904
rect 26200 19864 26206 19876
rect 25317 19839 25375 19845
rect 25317 19836 25329 19839
rect 25188 19808 25329 19836
rect 25188 19796 25194 19808
rect 25317 19805 25329 19808
rect 25363 19805 25375 19839
rect 25317 19799 25375 19805
rect 25593 19839 25651 19845
rect 25593 19805 25605 19839
rect 25639 19836 25651 19839
rect 25774 19836 25780 19848
rect 25639 19808 25780 19836
rect 25639 19805 25651 19808
rect 25593 19799 25651 19805
rect 24903 19740 25084 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 22152 19672 22324 19700
rect 22152 19660 22158 19672
rect 23474 19660 23480 19712
rect 23532 19660 23538 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 25038 19700 25044 19712
rect 23808 19672 25044 19700
rect 23808 19660 23814 19672
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 25608 19700 25636 19799
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 26252 19845 26280 19876
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 26973 19907 27031 19913
rect 26973 19904 26985 19907
rect 26384 19876 26985 19904
rect 26384 19864 26390 19876
rect 26973 19873 26985 19876
rect 27019 19873 27031 19907
rect 26973 19867 27031 19873
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19805 26295 19839
rect 26237 19799 26295 19805
rect 26510 19796 26516 19848
rect 26568 19796 26574 19848
rect 26602 19796 26608 19848
rect 26660 19836 26666 19848
rect 26660 19808 27016 19836
rect 26660 19796 26666 19808
rect 26988 19780 27016 19808
rect 26326 19728 26332 19780
rect 26384 19768 26390 19780
rect 26421 19771 26479 19777
rect 26421 19768 26433 19771
rect 26384 19740 26433 19768
rect 26384 19728 26390 19740
rect 26421 19737 26433 19740
rect 26467 19737 26479 19771
rect 26421 19731 26479 19737
rect 26878 19728 26884 19780
rect 26936 19728 26942 19780
rect 26970 19728 26976 19780
rect 27028 19728 27034 19780
rect 27080 19768 27108 19944
rect 27172 19845 27200 20012
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 27890 20000 27896 20052
rect 27948 20000 27954 20052
rect 28169 20043 28227 20049
rect 28169 20009 28181 20043
rect 28215 20040 28227 20043
rect 28350 20040 28356 20052
rect 28215 20012 28356 20040
rect 28215 20009 28227 20012
rect 28169 20003 28227 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 27246 19932 27252 19984
rect 27304 19972 27310 19984
rect 27341 19975 27399 19981
rect 27341 19972 27353 19975
rect 27304 19944 27353 19972
rect 27304 19932 27310 19944
rect 27341 19941 27353 19944
rect 27387 19941 27399 19975
rect 27341 19935 27399 19941
rect 27430 19864 27436 19916
rect 27488 19904 27494 19916
rect 27525 19907 27583 19913
rect 27525 19904 27537 19907
rect 27488 19876 27537 19904
rect 27488 19864 27494 19876
rect 27525 19873 27537 19876
rect 27571 19904 27583 19907
rect 29178 19904 29184 19916
rect 27571 19876 29184 19904
rect 27571 19873 27583 19876
rect 27525 19867 27583 19873
rect 29178 19864 29184 19876
rect 29236 19864 29242 19916
rect 27157 19839 27215 19845
rect 27157 19805 27169 19839
rect 27203 19805 27215 19839
rect 27709 19839 27767 19845
rect 27709 19836 27721 19839
rect 27157 19799 27215 19805
rect 27264 19808 27721 19836
rect 27264 19768 27292 19808
rect 27709 19805 27721 19808
rect 27755 19805 27767 19839
rect 27973 19839 28031 19845
rect 27973 19836 27985 19839
rect 27709 19799 27767 19805
rect 27908 19808 27985 19836
rect 27080 19740 27292 19768
rect 27430 19728 27436 19780
rect 27488 19728 27494 19780
rect 27908 19768 27936 19808
rect 27973 19805 27985 19808
rect 28019 19805 28031 19839
rect 27973 19799 28031 19805
rect 28074 19796 28080 19848
rect 28132 19796 28138 19848
rect 28258 19796 28264 19848
rect 28316 19836 28322 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28316 19808 28457 19836
rect 28316 19796 28322 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19836 28687 19839
rect 29086 19836 29092 19848
rect 28675 19808 29092 19836
rect 28675 19805 28687 19808
rect 28629 19799 28687 19805
rect 29086 19796 29092 19808
rect 29144 19796 29150 19848
rect 28718 19768 28724 19780
rect 27908 19740 28724 19768
rect 28718 19728 28724 19740
rect 28776 19728 28782 19780
rect 25179 19672 25636 19700
rect 26789 19703 26847 19709
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 26789 19669 26801 19703
rect 26835 19700 26847 19703
rect 27706 19700 27712 19712
rect 26835 19672 27712 19700
rect 26835 19669 26847 19672
rect 26789 19663 26847 19669
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 28350 19660 28356 19712
rect 28408 19660 28414 19712
rect 28810 19660 28816 19712
rect 28868 19660 28874 19712
rect 1104 19610 43884 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 43884 19610
rect 1104 19536 43884 19558
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3237 19499 3295 19505
rect 3237 19496 3249 19499
rect 3108 19468 3249 19496
rect 3108 19456 3114 19468
rect 3237 19465 3249 19468
rect 3283 19465 3295 19499
rect 3237 19459 3295 19465
rect 3326 19456 3332 19508
rect 3384 19456 3390 19508
rect 3697 19499 3755 19505
rect 3697 19465 3709 19499
rect 3743 19496 3755 19499
rect 3786 19496 3792 19508
rect 3743 19468 3792 19496
rect 3743 19465 3755 19468
rect 3697 19459 3755 19465
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 4249 19499 4307 19505
rect 4249 19465 4261 19499
rect 4295 19496 4307 19499
rect 5718 19496 5724 19508
rect 4295 19468 5724 19496
rect 4295 19465 4307 19468
rect 4249 19459 4307 19465
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 6270 19456 6276 19508
rect 6328 19496 6334 19508
rect 6730 19496 6736 19508
rect 6328 19468 6736 19496
rect 6328 19456 6334 19468
rect 6730 19456 6736 19468
rect 6788 19496 6794 19508
rect 6917 19499 6975 19505
rect 6917 19496 6929 19499
rect 6788 19468 6929 19496
rect 6788 19456 6794 19468
rect 1765 19431 1823 19437
rect 1765 19397 1777 19431
rect 1811 19428 1823 19431
rect 2102 19431 2160 19437
rect 2102 19428 2114 19431
rect 1811 19400 2114 19428
rect 1811 19397 1823 19400
rect 1765 19391 1823 19397
rect 2102 19397 2114 19400
rect 2148 19397 2160 19431
rect 3344 19428 3372 19456
rect 3344 19400 4476 19428
rect 2102 19391 2160 19397
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 3510 19360 3516 19372
rect 1627 19332 3516 19360
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4062 19360 4068 19372
rect 3835 19332 4068 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 4448 19369 4476 19400
rect 5350 19388 5356 19440
rect 5408 19388 5414 19440
rect 5736 19428 5764 19456
rect 6638 19428 6644 19440
rect 5552 19400 5764 19428
rect 6564 19400 6644 19428
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 4617 19363 4675 19369
rect 4617 19360 4629 19363
rect 4580 19332 4629 19360
rect 4580 19320 4586 19332
rect 4617 19329 4629 19332
rect 4663 19360 4675 19363
rect 4798 19360 4804 19372
rect 4663 19332 4804 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 4982 19320 4988 19372
rect 5040 19320 5046 19372
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1486 19292 1492 19304
rect 1443 19264 1492 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1486 19252 1492 19264
rect 1544 19252 1550 19304
rect 1762 19252 1768 19304
rect 1820 19292 1826 19304
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1820 19264 1869 19292
rect 1820 19252 1826 19264
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 3878 19252 3884 19304
rect 3936 19252 3942 19304
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19292 4215 19295
rect 4893 19295 4951 19301
rect 4203 19264 4844 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 1504 19156 1532 19252
rect 4246 19224 4252 19236
rect 3252 19196 4252 19224
rect 2866 19156 2872 19168
rect 1504 19128 2872 19156
rect 2866 19116 2872 19128
rect 2924 19156 2930 19168
rect 3252 19156 3280 19196
rect 4246 19184 4252 19196
rect 4304 19184 4310 19236
rect 4816 19224 4844 19264
rect 4893 19261 4905 19295
rect 4939 19292 4951 19295
rect 5166 19292 5172 19304
rect 4939 19264 5172 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5258 19252 5264 19304
rect 5316 19252 5322 19304
rect 5276 19224 5304 19252
rect 4816 19196 5304 19224
rect 5368 19224 5396 19388
rect 5442 19320 5448 19372
rect 5500 19320 5506 19372
rect 5552 19301 5580 19400
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19360 5779 19363
rect 5810 19360 5816 19372
rect 5767 19332 5816 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 6089 19363 6147 19369
rect 6089 19360 6101 19363
rect 6052 19332 6101 19360
rect 6052 19320 6058 19332
rect 6089 19329 6101 19332
rect 6135 19329 6147 19363
rect 6089 19323 6147 19329
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6564 19369 6592 19400
rect 6638 19388 6644 19400
rect 6696 19388 6702 19440
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19261 5595 19295
rect 5537 19255 5595 19261
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 5644 19224 5672 19255
rect 5368 19196 5672 19224
rect 6380 19224 6408 19323
rect 6840 19292 6868 19468
rect 6917 19465 6929 19468
rect 6963 19465 6975 19499
rect 6917 19459 6975 19465
rect 7285 19499 7343 19505
rect 7285 19465 7297 19499
rect 7331 19496 7343 19499
rect 7374 19496 7380 19508
rect 7331 19468 7380 19496
rect 7331 19465 7343 19468
rect 7285 19459 7343 19465
rect 7374 19456 7380 19468
rect 7432 19456 7438 19508
rect 8294 19456 8300 19508
rect 8352 19456 8358 19508
rect 8478 19456 8484 19508
rect 8536 19456 8542 19508
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 8864 19468 9260 19496
rect 8312 19428 8340 19456
rect 7116 19400 8340 19428
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7116 19369 7144 19400
rect 7101 19363 7159 19369
rect 7101 19360 7113 19363
rect 6972 19332 7113 19360
rect 6972 19320 6978 19332
rect 7101 19329 7113 19332
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7190 19320 7196 19372
rect 7248 19360 7254 19372
rect 8772 19369 8800 19456
rect 8864 19437 8892 19468
rect 8849 19431 8907 19437
rect 8849 19397 8861 19431
rect 8895 19397 8907 19431
rect 9232 19428 9260 19468
rect 9398 19456 9404 19508
rect 9456 19456 9462 19508
rect 9490 19456 9496 19508
rect 9548 19456 9554 19508
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19465 9643 19499
rect 9585 19459 9643 19465
rect 9600 19428 9628 19459
rect 10502 19456 10508 19508
rect 10560 19456 10566 19508
rect 10686 19456 10692 19508
rect 10744 19456 10750 19508
rect 11330 19456 11336 19508
rect 11388 19456 11394 19508
rect 12342 19496 12348 19508
rect 11624 19468 12348 19496
rect 9232 19400 9628 19428
rect 8849 19391 8907 19397
rect 10134 19388 10140 19440
rect 10192 19428 10198 19440
rect 10520 19428 10548 19456
rect 11624 19437 11652 19468
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 12526 19456 12532 19508
rect 12584 19456 12590 19508
rect 12618 19456 12624 19508
rect 12676 19456 12682 19508
rect 12710 19456 12716 19508
rect 12768 19496 12774 19508
rect 15102 19496 15108 19508
rect 12768 19468 12940 19496
rect 12768 19456 12774 19468
rect 11609 19431 11667 19437
rect 11609 19428 11621 19431
rect 10192 19400 10456 19428
rect 10520 19400 11621 19428
rect 10192 19388 10198 19400
rect 9122 19369 9128 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 7248 19332 7297 19360
rect 7248 19320 7254 19332
rect 7285 19329 7297 19332
rect 7331 19329 7343 19363
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 7285 19323 7343 19329
rect 7944 19332 8585 19360
rect 7944 19301 7972 19332
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 9079 19363 9128 19369
rect 9079 19329 9091 19363
rect 9125 19329 9128 19363
rect 9079 19323 9128 19329
rect 7929 19295 7987 19301
rect 6840 19264 7880 19292
rect 6546 19224 6552 19236
rect 6380 19196 6552 19224
rect 6546 19184 6552 19196
rect 6604 19184 6610 19236
rect 7282 19184 7288 19236
rect 7340 19224 7346 19236
rect 7650 19224 7656 19236
rect 7340 19196 7656 19224
rect 7340 19184 7346 19196
rect 7650 19184 7656 19196
rect 7708 19184 7714 19236
rect 7852 19224 7880 19264
rect 7929 19261 7941 19295
rect 7975 19261 7987 19295
rect 7929 19255 7987 19261
rect 8754 19224 8760 19236
rect 7852 19196 8760 19224
rect 8754 19184 8760 19196
rect 8812 19224 8818 19236
rect 8956 19224 8984 19323
rect 9122 19320 9128 19323
rect 9180 19320 9186 19372
rect 9306 19320 9312 19372
rect 9364 19320 9370 19372
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 10318 19360 10324 19372
rect 9723 19332 10324 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10428 19360 10456 19400
rect 11609 19397 11621 19400
rect 11655 19397 11667 19431
rect 11609 19391 11667 19397
rect 12066 19388 12072 19440
rect 12124 19388 12130 19440
rect 12158 19388 12164 19440
rect 12216 19428 12222 19440
rect 12544 19428 12572 19456
rect 12912 19437 12940 19468
rect 13372 19468 15108 19496
rect 12897 19431 12955 19437
rect 12216 19400 12480 19428
rect 12544 19400 12848 19428
rect 12216 19388 12222 19400
rect 11698 19360 11704 19372
rect 10428 19332 11704 19360
rect 11698 19320 11704 19332
rect 11756 19360 11762 19372
rect 11974 19360 11980 19372
rect 11756 19332 11980 19360
rect 11756 19320 11762 19332
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12084 19334 12112 19388
rect 12084 19306 12204 19334
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12345 19363 12403 19369
rect 12345 19360 12357 19363
rect 12308 19332 12357 19360
rect 12308 19320 12314 19332
rect 12345 19329 12357 19332
rect 12391 19329 12403 19363
rect 12452 19360 12480 19400
rect 12820 19369 12848 19400
rect 12897 19397 12909 19431
rect 12943 19397 12955 19431
rect 12897 19391 12955 19397
rect 12986 19388 12992 19440
rect 13044 19388 13050 19440
rect 12529 19363 12587 19369
rect 12529 19360 12541 19363
rect 12452 19332 12541 19360
rect 12345 19323 12403 19329
rect 12529 19329 12541 19332
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 13107 19363 13165 19369
rect 13107 19329 13119 19363
rect 13153 19329 13165 19363
rect 13107 19323 13165 19329
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 9048 19264 9229 19292
rect 9048 19236 9076 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 10042 19252 10048 19304
rect 10100 19252 10106 19304
rect 10134 19252 10140 19304
rect 10192 19292 10198 19304
rect 11514 19292 11520 19304
rect 10192 19264 11520 19292
rect 10192 19252 10198 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 11885 19295 11943 19301
rect 11885 19261 11897 19295
rect 11931 19261 11943 19295
rect 11885 19255 11943 19261
rect 8812 19196 8984 19224
rect 8812 19184 8818 19196
rect 9030 19184 9036 19236
rect 9088 19184 9094 19236
rect 9122 19184 9128 19236
rect 9180 19224 9186 19236
rect 10502 19224 10508 19236
rect 9180 19196 10508 19224
rect 9180 19184 9186 19196
rect 10502 19184 10508 19196
rect 10560 19184 10566 19236
rect 11900 19224 11928 19255
rect 12176 19224 12204 19306
rect 11900 19196 12204 19224
rect 2924 19128 3280 19156
rect 2924 19116 2930 19128
rect 3326 19116 3332 19168
rect 3384 19116 3390 19168
rect 5261 19159 5319 19165
rect 5261 19125 5273 19159
rect 5307 19156 5319 19159
rect 5534 19156 5540 19168
rect 5307 19128 5540 19156
rect 5307 19125 5319 19128
rect 5261 19119 5319 19125
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 5905 19159 5963 19165
rect 5905 19156 5917 19159
rect 5868 19128 5917 19156
rect 5868 19116 5874 19128
rect 5905 19125 5917 19128
rect 5951 19125 5963 19159
rect 5905 19119 5963 19125
rect 6454 19116 6460 19168
rect 6512 19116 6518 19168
rect 7745 19159 7803 19165
rect 7745 19125 7757 19159
rect 7791 19156 7803 19159
rect 8846 19156 8852 19168
rect 7791 19128 8852 19156
rect 7791 19125 7803 19128
rect 7745 19119 7803 19125
rect 8846 19116 8852 19128
rect 8904 19156 8910 19168
rect 12268 19156 12296 19320
rect 12544 19224 12572 19323
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 13122 19292 13150 19323
rect 13262 19320 13268 19372
rect 13320 19320 13326 19372
rect 12676 19264 13150 19292
rect 12676 19252 12682 19264
rect 12710 19224 12716 19236
rect 12544 19196 12716 19224
rect 12710 19184 12716 19196
rect 12768 19224 12774 19236
rect 13372 19224 13400 19468
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 15746 19496 15752 19508
rect 15580 19468 15752 19496
rect 14090 19388 14096 19440
rect 14148 19388 14154 19440
rect 15378 19428 15384 19440
rect 15304 19400 15384 19428
rect 13633 19363 13691 19369
rect 13633 19329 13645 19363
rect 13679 19360 13691 19363
rect 13817 19363 13875 19369
rect 13679 19332 13768 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 13740 19236 13768 19332
rect 13817 19329 13829 19363
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 12768 19196 13400 19224
rect 12768 19184 12774 19196
rect 13446 19184 13452 19236
rect 13504 19224 13510 19236
rect 13722 19224 13728 19236
rect 13504 19196 13728 19224
rect 13504 19184 13510 19196
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 13832 19168 13860 19323
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 15304 19369 15332 19400
rect 15378 19388 15384 19400
rect 15436 19388 15442 19440
rect 15580 19437 15608 19468
rect 15746 19456 15752 19468
rect 15804 19496 15810 19508
rect 16666 19496 16672 19508
rect 15804 19468 16672 19496
rect 15804 19456 15810 19468
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 16758 19456 16764 19508
rect 16816 19456 16822 19508
rect 18782 19496 18788 19508
rect 17696 19468 18788 19496
rect 15565 19431 15623 19437
rect 15565 19397 15577 19431
rect 15611 19397 15623 19431
rect 15565 19391 15623 19397
rect 15856 19400 17172 19428
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14516 19332 14841 19360
rect 14516 19320 14522 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 15856 19360 15884 19400
rect 17144 19372 17172 19400
rect 15519 19332 15884 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15988 19332 16681 19360
rect 15988 19320 15994 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 17126 19320 17132 19372
rect 17184 19320 17190 19372
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17696 19369 17724 19468
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19242 19496 19248 19508
rect 18892 19468 19248 19496
rect 17770 19388 17776 19440
rect 17828 19428 17834 19440
rect 18892 19428 18920 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 19392 19468 21680 19496
rect 19392 19456 19398 19468
rect 19150 19428 19156 19440
rect 17828 19400 18920 19428
rect 18984 19400 19156 19428
rect 17828 19388 17834 19400
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 17276 19332 17325 19360
rect 17276 19320 17282 19332
rect 17313 19329 17325 19332
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 18322 19360 18328 19372
rect 17681 19323 17739 19329
rect 17880 19332 18328 19360
rect 14918 19292 14924 19304
rect 14016 19264 14924 19292
rect 13909 19227 13967 19233
rect 13909 19193 13921 19227
rect 13955 19224 13967 19227
rect 14016 19224 14044 19264
rect 14918 19252 14924 19264
rect 14976 19252 14982 19304
rect 15378 19252 15384 19304
rect 15436 19252 15442 19304
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19292 16359 19295
rect 17034 19292 17040 19304
rect 16347 19264 17040 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 16316 19224 16344 19255
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 13955 19196 14044 19224
rect 15396 19196 16344 19224
rect 17420 19224 17448 19323
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 17880 19292 17908 19332
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18708 19369 18736 19400
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 18984 19369 19012 19400
rect 19150 19388 19156 19400
rect 19208 19428 19214 19440
rect 19208 19400 19840 19428
rect 19208 19388 19214 19400
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18840 19332 18981 19360
rect 18840 19320 18846 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19392 19332 19717 19360
rect 19392 19320 19398 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19812 19360 19840 19400
rect 19886 19388 19892 19440
rect 19944 19428 19950 19440
rect 20622 19428 20628 19440
rect 19944 19400 20116 19428
rect 19944 19388 19950 19400
rect 19978 19360 19984 19372
rect 19812 19332 19984 19360
rect 19705 19323 19763 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 18230 19292 18236 19304
rect 17635 19264 17908 19292
rect 17972 19264 18236 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 17494 19224 17500 19236
rect 17420 19196 17500 19224
rect 13955 19193 13967 19196
rect 13909 19187 13967 19193
rect 15396 19168 15424 19196
rect 17494 19184 17500 19196
rect 17552 19224 17558 19236
rect 17972 19224 18000 19264
rect 18230 19252 18236 19264
rect 18288 19292 18294 19304
rect 18414 19292 18420 19304
rect 18288 19264 18420 19292
rect 18288 19252 18294 19264
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18874 19252 18880 19304
rect 18932 19292 18938 19304
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 18932 19264 19257 19292
rect 18932 19252 18938 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19292 19671 19295
rect 20088 19292 20116 19400
rect 20180 19400 20628 19428
rect 20180 19369 20208 19400
rect 20622 19388 20628 19400
rect 20680 19428 20686 19440
rect 20680 19400 20760 19428
rect 20680 19388 20686 19400
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 20530 19320 20536 19372
rect 20588 19320 20594 19372
rect 20732 19369 20760 19400
rect 20806 19388 20812 19440
rect 20864 19388 20870 19440
rect 21269 19431 21327 19437
rect 21269 19397 21281 19431
rect 21315 19428 21327 19431
rect 21542 19428 21548 19440
rect 21315 19400 21548 19428
rect 21315 19397 21327 19400
rect 21269 19391 21327 19397
rect 21542 19388 21548 19400
rect 21600 19388 21606 19440
rect 21652 19428 21680 19468
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 22646 19496 22652 19508
rect 21968 19468 22652 19496
rect 21968 19456 21974 19468
rect 22646 19456 22652 19468
rect 22704 19456 22710 19508
rect 23106 19456 23112 19508
rect 23164 19456 23170 19508
rect 23400 19468 24256 19496
rect 23400 19437 23428 19468
rect 23385 19431 23443 19437
rect 23385 19428 23397 19431
rect 21652 19400 23397 19428
rect 23385 19397 23397 19400
rect 23431 19397 23443 19431
rect 23385 19391 23443 19397
rect 23566 19388 23572 19440
rect 23624 19428 23630 19440
rect 23624 19400 23888 19428
rect 23624 19388 23630 19400
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 21082 19320 21088 19372
rect 21140 19320 21146 19372
rect 21726 19320 21732 19372
rect 21784 19360 21790 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21784 19332 21833 19360
rect 21784 19320 21790 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21821 19323 21879 19329
rect 21928 19332 22569 19360
rect 20257 19295 20315 19301
rect 20257 19292 20269 19295
rect 19659 19264 20030 19292
rect 20088 19264 20269 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 17552 19196 18000 19224
rect 17552 19184 17558 19196
rect 18138 19184 18144 19236
rect 18196 19184 18202 19236
rect 8904 19128 12296 19156
rect 8904 19116 8910 19128
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13814 19156 13820 19168
rect 12860 19128 13820 19156
rect 12860 19116 12866 19128
rect 13814 19116 13820 19128
rect 13872 19156 13878 19168
rect 14642 19156 14648 19168
rect 13872 19128 14648 19156
rect 13872 19116 13878 19128
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 15378 19116 15384 19168
rect 15436 19116 15442 19168
rect 17129 19159 17187 19165
rect 17129 19125 17141 19159
rect 17175 19156 17187 19159
rect 18892 19156 18920 19252
rect 19150 19184 19156 19236
rect 19208 19224 19214 19236
rect 19702 19224 19708 19236
rect 19208 19196 19708 19224
rect 19208 19184 19214 19196
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 20002 19224 20030 19264
rect 20257 19261 20269 19264
rect 20303 19261 20315 19295
rect 20548 19292 20576 19320
rect 21928 19292 21956 19332
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 23676 19369 23704 19400
rect 23477 19363 23535 19369
rect 23477 19329 23489 19363
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 23661 19363 23719 19369
rect 23661 19329 23673 19363
rect 23707 19329 23719 19363
rect 23661 19323 23719 19329
rect 22094 19292 22100 19304
rect 20548 19264 21956 19292
rect 22024 19264 22100 19292
rect 20257 19255 20315 19261
rect 20002 19196 20116 19224
rect 20088 19168 20116 19196
rect 17175 19128 18920 19156
rect 17175 19125 17187 19128
rect 17129 19119 17187 19125
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19889 19159 19947 19165
rect 19889 19156 19901 19159
rect 19024 19128 19901 19156
rect 19024 19116 19030 19128
rect 19889 19125 19901 19128
rect 19935 19125 19947 19159
rect 19889 19119 19947 19125
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 20272 19156 20300 19255
rect 20806 19184 20812 19236
rect 20864 19224 20870 19236
rect 21450 19224 21456 19236
rect 20864 19196 21456 19224
rect 20864 19184 20870 19196
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 22024 19224 22052 19264
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 22278 19252 22284 19304
rect 22336 19292 22342 19304
rect 23492 19292 23520 19323
rect 23750 19320 23756 19372
rect 23808 19320 23814 19372
rect 23860 19369 23888 19400
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 24228 19437 24256 19468
rect 24394 19456 24400 19508
rect 24452 19456 24458 19508
rect 24489 19499 24547 19505
rect 24489 19465 24501 19499
rect 24535 19496 24547 19499
rect 25314 19496 25320 19508
rect 24535 19468 25320 19496
rect 24535 19465 24547 19468
rect 24489 19459 24547 19465
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 25409 19499 25467 19505
rect 25409 19465 25421 19499
rect 25455 19496 25467 19499
rect 25590 19496 25596 19508
rect 25455 19468 25596 19496
rect 25455 19465 25467 19468
rect 25409 19459 25467 19465
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 25682 19456 25688 19508
rect 25740 19496 25746 19508
rect 25740 19468 28212 19496
rect 25740 19456 25746 19468
rect 24213 19431 24271 19437
rect 24213 19397 24225 19431
rect 24259 19397 24271 19431
rect 24412 19428 24440 19456
rect 25041 19431 25099 19437
rect 25041 19428 25053 19431
rect 24412 19400 25053 19428
rect 24213 19391 24271 19397
rect 25041 19397 25053 19400
rect 25087 19428 25099 19431
rect 27249 19431 27307 19437
rect 27249 19428 27261 19431
rect 25087 19400 27261 19428
rect 25087 19397 25099 19400
rect 25041 19391 25099 19397
rect 27249 19397 27261 19400
rect 27295 19397 27307 19431
rect 27249 19391 27307 19397
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 23934 19320 23940 19372
rect 23992 19360 23998 19372
rect 23992 19332 24037 19360
rect 23992 19320 23998 19332
rect 22336 19264 24164 19292
rect 22336 19252 22342 19264
rect 22646 19224 22652 19236
rect 21836 19196 22052 19224
rect 22103 19196 22652 19224
rect 21836 19156 21864 19196
rect 20272 19128 21864 19156
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22103 19156 22131 19196
rect 22646 19184 22652 19196
rect 22704 19224 22710 19236
rect 23474 19224 23480 19236
rect 22704 19196 23480 19224
rect 22704 19184 22710 19196
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 21968 19128 22131 19156
rect 24136 19156 24164 19264
rect 24228 19224 24256 19391
rect 27338 19388 27344 19440
rect 27396 19388 27402 19440
rect 27614 19388 27620 19440
rect 27672 19428 27678 19440
rect 27709 19431 27767 19437
rect 27709 19428 27721 19431
rect 27672 19400 27721 19428
rect 27672 19388 27678 19400
rect 27709 19397 27721 19400
rect 27755 19397 27767 19431
rect 27709 19391 27767 19397
rect 24349 19363 24407 19369
rect 24349 19329 24361 19363
rect 24395 19360 24407 19363
rect 24670 19360 24676 19372
rect 24395 19332 24676 19360
rect 24395 19329 24407 19332
rect 24349 19323 24407 19329
rect 24670 19320 24676 19332
rect 24728 19360 24734 19372
rect 24857 19363 24915 19369
rect 24857 19360 24869 19363
rect 24728 19332 24869 19360
rect 24728 19320 24734 19332
rect 24857 19329 24869 19332
rect 24903 19329 24915 19363
rect 24857 19323 24915 19329
rect 24946 19320 24952 19372
rect 25004 19360 25010 19372
rect 25133 19363 25191 19369
rect 25133 19360 25145 19363
rect 25004 19332 25145 19360
rect 25004 19320 25010 19332
rect 25133 19329 25145 19332
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 24946 19224 24952 19236
rect 24228 19196 24952 19224
rect 24946 19184 24952 19196
rect 25004 19184 25010 19236
rect 25240 19224 25268 19323
rect 25314 19320 25320 19372
rect 25372 19360 25378 19372
rect 26513 19363 26571 19369
rect 26513 19360 26525 19363
rect 25372 19332 26525 19360
rect 25372 19320 25378 19332
rect 26513 19329 26525 19332
rect 26559 19329 26571 19363
rect 26513 19323 26571 19329
rect 26602 19320 26608 19372
rect 26660 19320 26666 19372
rect 26962 19363 27020 19369
rect 26962 19360 26974 19363
rect 26804 19332 26974 19360
rect 25958 19252 25964 19304
rect 26016 19252 26022 19304
rect 26620 19292 26648 19320
rect 26804 19292 26832 19332
rect 26962 19329 26974 19332
rect 27008 19329 27020 19363
rect 26962 19323 27020 19329
rect 27066 19363 27124 19369
rect 27066 19329 27078 19363
rect 27112 19329 27124 19363
rect 27066 19323 27124 19329
rect 27438 19363 27496 19369
rect 27438 19329 27450 19363
rect 27484 19329 27496 19363
rect 27985 19363 28043 19369
rect 27985 19360 27997 19363
rect 27438 19323 27496 19329
rect 27632 19332 27997 19360
rect 27080 19306 27109 19323
rect 27080 19292 27108 19306
rect 26620 19264 26832 19292
rect 26988 19264 27108 19292
rect 26142 19224 26148 19236
rect 25240 19196 26148 19224
rect 26142 19184 26148 19196
rect 26200 19184 26206 19236
rect 24578 19156 24584 19168
rect 24136 19128 24584 19156
rect 21968 19116 21974 19128
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 26160 19156 26188 19184
rect 26988 19156 27016 19264
rect 27246 19252 27252 19304
rect 27304 19292 27310 19304
rect 27453 19292 27481 19323
rect 27304 19264 27481 19292
rect 27304 19252 27310 19264
rect 27632 19233 27660 19332
rect 27908 19329 27997 19332
rect 28031 19329 28043 19363
rect 28184 19360 28212 19468
rect 28442 19456 28448 19508
rect 28500 19456 28506 19508
rect 28626 19456 28632 19508
rect 28684 19456 28690 19508
rect 28460 19428 28488 19456
rect 28368 19400 28488 19428
rect 28261 19363 28319 19369
rect 28261 19360 28273 19363
rect 28184 19332 28273 19360
rect 27908 19323 28043 19329
rect 28261 19329 28273 19332
rect 28307 19329 28319 19363
rect 28261 19323 28319 19329
rect 27908 19306 28028 19323
rect 27798 19252 27804 19304
rect 27856 19252 27862 19304
rect 28000 19292 28028 19306
rect 28368 19292 28396 19400
rect 28445 19363 28503 19369
rect 28445 19329 28457 19363
rect 28491 19329 28503 19363
rect 28445 19323 28503 19329
rect 28000 19264 28396 19292
rect 27617 19227 27675 19233
rect 27617 19193 27629 19227
rect 27663 19193 27675 19227
rect 28460 19224 28488 19323
rect 27617 19187 27675 19193
rect 27724 19196 28488 19224
rect 27724 19168 27752 19196
rect 27246 19156 27252 19168
rect 26160 19128 27252 19156
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 27706 19116 27712 19168
rect 27764 19116 27770 19168
rect 28166 19116 28172 19168
rect 28224 19116 28230 19168
rect 1104 19066 43884 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 43884 19066
rect 1104 18992 43884 19014
rect 3510 18912 3516 18964
rect 3568 18912 3574 18964
rect 4062 18952 4068 18964
rect 3804 18924 4068 18952
rect 3804 18884 3832 18924
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 5224 18924 5365 18952
rect 5224 18912 5230 18924
rect 5353 18921 5365 18924
rect 5399 18921 5411 18955
rect 5353 18915 5411 18921
rect 5902 18912 5908 18964
rect 5960 18952 5966 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 5960 18924 6745 18952
rect 5960 18912 5966 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 6733 18915 6791 18921
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 8386 18952 8392 18964
rect 7892 18924 8392 18952
rect 7892 18912 7898 18924
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 9493 18955 9551 18961
rect 9493 18952 9505 18955
rect 8812 18924 9505 18952
rect 8812 18912 8818 18924
rect 9493 18921 9505 18924
rect 9539 18921 9551 18955
rect 9493 18915 9551 18921
rect 6086 18884 6092 18896
rect 1596 18856 3832 18884
rect 5920 18856 6092 18884
rect 1596 18757 1624 18856
rect 1854 18776 1860 18828
rect 1912 18816 1918 18828
rect 3789 18819 3847 18825
rect 3789 18816 3801 18819
rect 1912 18788 3801 18816
rect 1912 18776 1918 18788
rect 3789 18785 3801 18788
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 5920 18825 5948 18856
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 6178 18844 6184 18896
rect 6236 18884 6242 18896
rect 8294 18884 8300 18896
rect 6236 18856 6868 18884
rect 6236 18844 6242 18856
rect 5905 18819 5963 18825
rect 5316 18788 5764 18816
rect 5316 18776 5322 18788
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18717 1639 18751
rect 1581 18711 1639 18717
rect 2682 18708 2688 18760
rect 2740 18708 2746 18760
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3326 18748 3332 18760
rect 3007 18720 3332 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 5626 18708 5632 18760
rect 5684 18708 5690 18760
rect 5736 18748 5764 18788
rect 5905 18785 5917 18819
rect 5951 18785 5963 18819
rect 6362 18816 6368 18828
rect 5905 18779 5963 18785
rect 6104 18788 6368 18816
rect 6104 18757 6132 18788
rect 6362 18776 6368 18788
rect 6420 18816 6426 18828
rect 6840 18816 6868 18856
rect 8266 18844 8300 18884
rect 8352 18844 8358 18896
rect 8266 18816 8294 18844
rect 6420 18788 6776 18816
rect 6420 18776 6426 18788
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 5736 18720 6101 18748
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 6178 18708 6184 18760
rect 6236 18708 6242 18760
rect 6457 18751 6515 18757
rect 6457 18748 6469 18751
rect 6288 18720 6469 18748
rect 1210 18640 1216 18692
rect 1268 18680 1274 18692
rect 2317 18683 2375 18689
rect 2317 18680 2329 18683
rect 1268 18652 2329 18680
rect 1268 18640 1274 18652
rect 2317 18649 2329 18652
rect 2363 18649 2375 18683
rect 2317 18643 2375 18649
rect 2700 18612 2728 18708
rect 6288 18692 6316 18720
rect 6457 18717 6469 18720
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 6546 18708 6552 18760
rect 6604 18757 6610 18760
rect 6604 18748 6612 18757
rect 6604 18720 6649 18748
rect 6604 18711 6612 18720
rect 6604 18708 6610 18711
rect 4056 18683 4114 18689
rect 4056 18649 4068 18683
rect 4102 18680 4114 18683
rect 4890 18680 4896 18692
rect 4102 18652 4896 18680
rect 4102 18649 4114 18652
rect 4056 18643 4114 18649
rect 4890 18640 4896 18652
rect 4948 18640 4954 18692
rect 5994 18640 6000 18692
rect 6052 18640 6058 18692
rect 6270 18640 6276 18692
rect 6328 18640 6334 18692
rect 6365 18683 6423 18689
rect 6365 18649 6377 18683
rect 6411 18649 6423 18683
rect 6569 18680 6597 18708
rect 6748 18680 6776 18788
rect 6840 18788 8294 18816
rect 6840 18757 6868 18788
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7006 18708 7012 18760
rect 7064 18708 7070 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 9398 18748 9404 18760
rect 8260 18720 9404 18748
rect 8260 18708 8266 18720
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 7926 18680 7932 18692
rect 6569 18652 6684 18680
rect 6748 18652 7932 18680
rect 6365 18643 6423 18649
rect 5074 18612 5080 18624
rect 2700 18584 5080 18612
rect 5074 18572 5080 18584
rect 5132 18612 5138 18624
rect 5169 18615 5227 18621
rect 5169 18612 5181 18615
rect 5132 18584 5181 18612
rect 5132 18572 5138 18584
rect 5169 18581 5181 18584
rect 5215 18581 5227 18615
rect 5169 18575 5227 18581
rect 5813 18615 5871 18621
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 6012 18612 6040 18640
rect 5859 18584 6040 18612
rect 6380 18612 6408 18643
rect 6546 18612 6552 18624
rect 6380 18584 6552 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 6656 18612 6684 18652
rect 7926 18640 7932 18652
rect 7984 18680 7990 18692
rect 8757 18683 8815 18689
rect 7984 18652 8708 18680
rect 7984 18640 7990 18652
rect 6730 18612 6736 18624
rect 6656 18584 6736 18612
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 6914 18572 6920 18624
rect 6972 18572 6978 18624
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 7558 18612 7564 18624
rect 7432 18584 7564 18612
rect 7432 18572 7438 18584
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 7650 18572 7656 18624
rect 7708 18572 7714 18624
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8386 18612 8392 18624
rect 8260 18584 8392 18612
rect 8260 18572 8266 18584
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 8680 18612 8708 18652
rect 8757 18649 8769 18683
rect 8803 18680 8815 18683
rect 8846 18680 8852 18692
rect 8803 18652 8852 18680
rect 8803 18649 8815 18652
rect 8757 18643 8815 18649
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9508 18680 9536 18915
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 11609 18955 11667 18961
rect 11609 18921 11621 18955
rect 11655 18952 11667 18955
rect 11698 18952 11704 18964
rect 11655 18924 11704 18952
rect 11655 18921 11667 18924
rect 11609 18915 11667 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 15010 18952 15016 18964
rect 12216 18924 15016 18952
rect 12216 18912 12222 18924
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 15473 18955 15531 18961
rect 15473 18921 15485 18955
rect 15519 18952 15531 18955
rect 15838 18952 15844 18964
rect 15519 18924 15844 18952
rect 15519 18921 15531 18924
rect 15473 18915 15531 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 15930 18912 15936 18964
rect 15988 18912 15994 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16172 18924 17632 18952
rect 16172 18912 16178 18924
rect 11514 18844 11520 18896
rect 11572 18884 11578 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 11572 18856 12725 18884
rect 11572 18844 11578 18856
rect 12713 18853 12725 18856
rect 12759 18884 12771 18887
rect 13078 18884 13084 18896
rect 12759 18856 13084 18884
rect 12759 18853 12771 18856
rect 12713 18847 12771 18853
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 13170 18844 13176 18896
rect 13228 18844 13234 18896
rect 13280 18856 14228 18884
rect 10689 18819 10747 18825
rect 10689 18785 10701 18819
rect 10735 18816 10747 18819
rect 10962 18816 10968 18828
rect 10735 18788 10968 18816
rect 10735 18785 10747 18788
rect 10689 18779 10747 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18816 11299 18819
rect 13280 18816 13308 18856
rect 14200 18816 14228 18856
rect 14274 18844 14280 18896
rect 14332 18884 14338 18896
rect 14369 18887 14427 18893
rect 14369 18884 14381 18887
rect 14332 18856 14381 18884
rect 14332 18844 14338 18856
rect 14369 18853 14381 18856
rect 14415 18853 14427 18887
rect 14369 18847 14427 18853
rect 14550 18844 14556 18896
rect 14608 18884 14614 18896
rect 14608 18856 16344 18884
rect 14608 18844 14614 18856
rect 15838 18816 15844 18828
rect 11287 18788 13308 18816
rect 13372 18788 14044 18816
rect 14200 18788 15844 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 10226 18708 10232 18760
rect 10284 18708 10290 18760
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 10928 18720 11529 18748
rect 10928 18708 10934 18720
rect 11517 18717 11529 18720
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12158 18748 12164 18760
rect 11756 18720 12164 18748
rect 11756 18708 11762 18720
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12308 18720 12357 18748
rect 12308 18708 12314 18720
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 13372 18757 13400 18788
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12768 18720 12817 18748
rect 12768 18708 12774 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 13814 18748 13820 18760
rect 13771 18720 13820 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18717 13967 18751
rect 14016 18748 14044 18788
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 16316 18760 16344 18856
rect 17310 18844 17316 18896
rect 17368 18884 17374 18896
rect 17497 18887 17555 18893
rect 17497 18884 17509 18887
rect 17368 18856 17509 18884
rect 17368 18844 17374 18856
rect 17497 18853 17509 18856
rect 17543 18853 17555 18887
rect 17604 18884 17632 18924
rect 17862 18912 17868 18964
rect 17920 18952 17926 18964
rect 19978 18952 19984 18964
rect 17920 18924 19984 18952
rect 17920 18912 17926 18924
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20254 18912 20260 18964
rect 20312 18952 20318 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 20312 18924 21005 18952
rect 20312 18912 20318 18924
rect 20993 18921 21005 18924
rect 21039 18921 21051 18955
rect 20993 18915 21051 18921
rect 21085 18955 21143 18961
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21821 18955 21879 18961
rect 21131 18924 21772 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21744 18896 21772 18924
rect 21821 18921 21833 18955
rect 21867 18952 21879 18955
rect 22189 18955 22247 18961
rect 21867 18924 22048 18952
rect 21867 18921 21879 18924
rect 21821 18915 21879 18921
rect 22020 18896 22048 18924
rect 22189 18921 22201 18955
rect 22235 18952 22247 18955
rect 22922 18952 22928 18964
rect 22235 18924 22928 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 23109 18955 23167 18961
rect 23109 18921 23121 18955
rect 23155 18952 23167 18955
rect 23382 18952 23388 18964
rect 23155 18924 23388 18952
rect 23155 18921 23167 18924
rect 23109 18915 23167 18921
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 24029 18955 24087 18961
rect 24029 18921 24041 18955
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 19705 18887 19763 18893
rect 17604 18856 19012 18884
rect 17497 18847 17555 18853
rect 17328 18816 17356 18844
rect 16408 18788 17356 18816
rect 17512 18788 18368 18816
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 14016 18720 14197 18748
rect 13909 18711 13967 18717
rect 14185 18717 14197 18720
rect 14231 18748 14243 18751
rect 14274 18748 14280 18760
rect 14231 18720 14280 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 10410 18680 10416 18692
rect 9508 18652 10416 18680
rect 10410 18640 10416 18652
rect 10468 18640 10474 18692
rect 10502 18640 10508 18692
rect 10560 18689 10566 18692
rect 10560 18683 10589 18689
rect 10577 18649 10589 18683
rect 10560 18643 10589 18649
rect 10560 18640 10566 18643
rect 11146 18640 11152 18692
rect 11204 18680 11210 18692
rect 11333 18683 11391 18689
rect 11333 18680 11345 18683
rect 11204 18652 11345 18680
rect 11204 18640 11210 18652
rect 11333 18649 11345 18652
rect 11379 18680 11391 18683
rect 13262 18680 13268 18692
rect 11379 18652 13268 18680
rect 11379 18649 11391 18652
rect 11333 18643 11391 18649
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 13633 18683 13691 18689
rect 13633 18649 13645 18683
rect 13679 18649 13691 18683
rect 13924 18680 13952 18711
rect 14274 18708 14280 18720
rect 14332 18748 14338 18760
rect 14332 18720 14964 18748
rect 14332 18708 14338 18720
rect 14550 18680 14556 18692
rect 13924 18652 14556 18680
rect 13633 18643 13691 18649
rect 9030 18612 9036 18624
rect 8680 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18612 9094 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 9088 18584 9137 18612
rect 9088 18572 9094 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9953 18615 10011 18621
rect 9953 18581 9965 18615
rect 9999 18612 10011 18615
rect 10962 18612 10968 18624
rect 9999 18584 10968 18612
rect 9999 18581 10011 18584
rect 9953 18575 10011 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 12158 18612 12164 18624
rect 11848 18584 12164 18612
rect 11848 18572 11854 18584
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12526 18612 12532 18624
rect 12391 18584 12532 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12897 18615 12955 18621
rect 12897 18581 12909 18615
rect 12943 18612 12955 18615
rect 13538 18612 13544 18624
rect 12943 18584 13544 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13648 18612 13676 18643
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 14936 18680 14964 18720
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 15746 18708 15752 18760
rect 15804 18708 15810 18760
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16114 18748 16120 18760
rect 16071 18720 16120 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16298 18708 16304 18760
rect 16356 18708 16362 18760
rect 16408 18757 16436 18788
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 16758 18748 16764 18760
rect 16684 18720 16764 18748
rect 16500 18680 16528 18708
rect 14936 18652 16528 18680
rect 13722 18612 13728 18624
rect 13648 18584 13728 18612
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 13814 18572 13820 18624
rect 13872 18572 13878 18624
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 14056 18584 15577 18612
rect 14056 18572 14062 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 16684 18612 16712 18720
rect 16758 18708 16764 18720
rect 16816 18748 16822 18760
rect 17512 18757 17540 18788
rect 18340 18760 18368 18788
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 18874 18816 18880 18828
rect 18656 18788 18880 18816
rect 18656 18776 18662 18788
rect 18874 18776 18880 18788
rect 18932 18776 18938 18828
rect 18984 18825 19012 18856
rect 19705 18853 19717 18887
rect 19751 18884 19763 18887
rect 21358 18884 21364 18896
rect 19751 18856 21364 18884
rect 19751 18853 19763 18856
rect 19705 18847 19763 18853
rect 21358 18844 21364 18856
rect 21416 18844 21422 18896
rect 21726 18844 21732 18896
rect 21784 18844 21790 18896
rect 22002 18844 22008 18896
rect 22060 18844 22066 18896
rect 22281 18887 22339 18893
rect 22281 18853 22293 18887
rect 22327 18884 22339 18887
rect 22462 18884 22468 18896
rect 22327 18856 22468 18884
rect 22327 18853 22339 18856
rect 22281 18847 22339 18853
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 23017 18887 23075 18893
rect 22572 18856 22876 18884
rect 18969 18819 19027 18825
rect 18969 18785 18981 18819
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 19300 18788 19748 18816
rect 19300 18776 19306 18788
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16816 18720 16865 18748
rect 16816 18708 16822 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17497 18751 17555 18757
rect 17359 18720 17448 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 15896 18584 16712 18612
rect 15896 18572 15902 18584
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17420 18612 17448 18720
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 17880 18680 17908 18711
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 18012 18720 18153 18748
rect 18012 18708 18018 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18380 18720 18521 18748
rect 18380 18708 18386 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 18782 18748 18788 18760
rect 18739 18720 18788 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 18248 18680 18276 18708
rect 17880 18652 18276 18680
rect 18414 18640 18420 18692
rect 18472 18640 18478 18692
rect 18708 18612 18736 18711
rect 18782 18708 18788 18720
rect 18840 18748 18846 18760
rect 19720 18757 19748 18788
rect 20254 18776 20260 18828
rect 20312 18776 20318 18828
rect 22186 18816 22192 18828
rect 21376 18788 22192 18816
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 18840 18720 19441 18748
rect 18840 18708 18846 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 19751 18720 20300 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 19889 18683 19947 18689
rect 19889 18680 19901 18683
rect 19576 18652 19901 18680
rect 19576 18640 19582 18652
rect 19889 18649 19901 18652
rect 19935 18649 19947 18683
rect 19889 18643 19947 18649
rect 17184 18584 18736 18612
rect 19904 18612 19932 18643
rect 20070 18640 20076 18692
rect 20128 18640 20134 18692
rect 20162 18612 20168 18624
rect 19904 18584 20168 18612
rect 17184 18572 17190 18584
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 20272 18612 20300 18720
rect 20346 18708 20352 18760
rect 20404 18708 20410 18760
rect 21376 18757 21404 18788
rect 22186 18776 22192 18788
rect 22244 18776 22250 18828
rect 22572 18816 22600 18856
rect 22480 18788 22600 18816
rect 22649 18819 22707 18825
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 20438 18612 20444 18624
rect 20272 18584 20444 18612
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 21284 18612 21312 18711
rect 21450 18708 21456 18760
rect 21508 18708 21514 18760
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 21910 18748 21916 18760
rect 21775 18720 21916 18748
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 21591 18683 21649 18689
rect 21591 18649 21603 18683
rect 21637 18680 21649 18683
rect 22480 18680 22508 18788
rect 22649 18785 22661 18819
rect 22695 18816 22707 18819
rect 22738 18816 22744 18828
rect 22695 18788 22744 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 22848 18757 22876 18856
rect 23017 18853 23029 18887
rect 23063 18884 23075 18887
rect 23474 18884 23480 18896
rect 23063 18856 23480 18884
rect 23063 18853 23075 18856
rect 23017 18847 23075 18853
rect 23474 18844 23480 18856
rect 23532 18844 23538 18896
rect 24044 18884 24072 18915
rect 24210 18912 24216 18964
rect 24268 18912 24274 18964
rect 24486 18912 24492 18964
rect 24544 18912 24550 18964
rect 24578 18912 24584 18964
rect 24636 18912 24642 18964
rect 25038 18912 25044 18964
rect 25096 18952 25102 18964
rect 25133 18955 25191 18961
rect 25133 18952 25145 18955
rect 25096 18924 25145 18952
rect 25096 18912 25102 18924
rect 25133 18921 25145 18924
rect 25179 18952 25191 18955
rect 25682 18952 25688 18964
rect 25179 18924 25688 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 25682 18912 25688 18924
rect 25740 18912 25746 18964
rect 26513 18955 26571 18961
rect 25977 18924 26464 18952
rect 24504 18884 24532 18912
rect 24044 18856 24532 18884
rect 24118 18816 24124 18828
rect 23308 18788 24124 18816
rect 23308 18757 23336 18788
rect 24118 18776 24124 18788
rect 24176 18816 24182 18828
rect 24596 18816 24624 18912
rect 24670 18844 24676 18896
rect 24728 18884 24734 18896
rect 24728 18856 25641 18884
rect 24728 18844 24734 18856
rect 25613 18816 25641 18856
rect 25977 18816 26005 18924
rect 26142 18844 26148 18896
rect 26200 18844 26206 18896
rect 26436 18884 26464 18924
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 26878 18952 26884 18964
rect 26559 18924 26884 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 26878 18912 26884 18924
rect 26936 18912 26942 18964
rect 29086 18912 29092 18964
rect 29144 18912 29150 18964
rect 26436 18856 26741 18884
rect 24176 18788 24532 18816
rect 24596 18788 25544 18816
rect 24176 18776 24182 18788
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18750 22615 18751
rect 22833 18751 22891 18757
rect 22603 18722 22692 18750
rect 22603 18717 22615 18722
rect 22557 18711 22615 18717
rect 21637 18652 22508 18680
rect 22664 18680 22692 18722
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 22879 18720 23305 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 23474 18708 23480 18760
rect 23532 18708 23538 18760
rect 23658 18757 23664 18760
rect 23615 18751 23664 18757
rect 23615 18717 23627 18751
rect 23661 18717 23664 18751
rect 23615 18711 23664 18717
rect 23658 18708 23664 18711
rect 23716 18708 23722 18760
rect 23750 18708 23756 18760
rect 23808 18708 23814 18760
rect 24026 18708 24032 18760
rect 24084 18748 24090 18760
rect 24302 18748 24308 18760
rect 24084 18720 24308 18748
rect 24084 18708 24090 18720
rect 23385 18683 23443 18689
rect 23385 18680 23397 18683
rect 22664 18652 23397 18680
rect 21637 18649 21649 18652
rect 21591 18643 21649 18649
rect 23124 18624 23152 18652
rect 23385 18649 23397 18652
rect 23431 18649 23443 18683
rect 23385 18643 23443 18649
rect 23842 18640 23848 18692
rect 23900 18640 23906 18692
rect 22186 18612 22192 18624
rect 21284 18584 22192 18612
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 22462 18572 22468 18624
rect 22520 18572 22526 18624
rect 23106 18572 23112 18624
rect 23164 18572 23170 18624
rect 23934 18572 23940 18624
rect 23992 18612 23998 18624
rect 24045 18615 24103 18621
rect 24045 18612 24057 18615
rect 23992 18584 24057 18612
rect 23992 18572 23998 18584
rect 24045 18581 24057 18584
rect 24091 18581 24103 18615
rect 24136 18612 24164 18720
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 24394 18708 24400 18760
rect 24452 18708 24458 18760
rect 24504 18748 24532 18788
rect 25516 18757 25544 18788
rect 25613 18788 26005 18816
rect 26160 18816 26188 18844
rect 26160 18788 26377 18816
rect 25613 18757 25641 18788
rect 25977 18757 26005 18788
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 24504 18720 25329 18748
rect 25317 18717 25329 18720
rect 25363 18717 25375 18751
rect 25317 18711 25375 18717
rect 25501 18751 25559 18757
rect 25501 18717 25513 18751
rect 25547 18717 25559 18751
rect 25613 18751 25677 18757
rect 25613 18720 25631 18751
rect 25501 18711 25559 18717
rect 25619 18717 25631 18720
rect 25665 18717 25677 18751
rect 25619 18711 25677 18717
rect 25777 18751 25835 18757
rect 25777 18717 25789 18751
rect 25823 18717 25835 18751
rect 25777 18711 25835 18717
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 25962 18751 26020 18757
rect 25962 18717 25974 18751
rect 26008 18717 26020 18751
rect 25962 18711 26020 18717
rect 24946 18640 24952 18692
rect 25004 18680 25010 18692
rect 25409 18683 25467 18689
rect 25409 18680 25421 18683
rect 25004 18652 25421 18680
rect 25004 18640 25010 18652
rect 25409 18649 25421 18652
rect 25455 18649 25467 18683
rect 25409 18643 25467 18649
rect 24857 18615 24915 18621
rect 24857 18612 24869 18615
rect 24136 18584 24869 18612
rect 24045 18575 24103 18581
rect 24857 18581 24869 18584
rect 24903 18581 24915 18615
rect 24857 18575 24915 18581
rect 25038 18572 25044 18624
rect 25096 18612 25102 18624
rect 25792 18612 25820 18711
rect 25884 18680 25912 18711
rect 26234 18708 26240 18760
rect 26292 18708 26298 18760
rect 26349 18757 26377 18788
rect 26713 18757 26741 18856
rect 26970 18844 26976 18896
rect 27028 18844 27034 18896
rect 26334 18751 26392 18757
rect 26334 18717 26346 18751
rect 26380 18717 26392 18751
rect 26605 18751 26663 18757
rect 26605 18742 26617 18751
rect 26334 18711 26392 18717
rect 26528 18717 26617 18742
rect 26651 18717 26663 18751
rect 26528 18714 26663 18717
rect 25884 18652 26004 18680
rect 25976 18624 26004 18652
rect 26142 18640 26148 18692
rect 26200 18640 26206 18692
rect 25096 18584 25820 18612
rect 25096 18572 25102 18584
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26050 18572 26056 18624
rect 26108 18612 26114 18624
rect 26528 18612 26556 18714
rect 26605 18711 26663 18714
rect 26698 18751 26756 18757
rect 26698 18717 26710 18751
rect 26744 18717 26756 18751
rect 26988 18748 27016 18844
rect 26698 18711 26756 18717
rect 26896 18720 27016 18748
rect 27070 18751 27128 18757
rect 26896 18689 26924 18720
rect 27070 18717 27082 18751
rect 27116 18748 27128 18751
rect 27246 18748 27252 18760
rect 27116 18720 27252 18748
rect 27116 18717 27128 18720
rect 27070 18711 27128 18717
rect 27246 18708 27252 18720
rect 27304 18708 27310 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 27982 18757 27988 18760
rect 27709 18751 27767 18757
rect 27709 18748 27721 18751
rect 27672 18720 27721 18748
rect 27672 18708 27678 18720
rect 27709 18717 27721 18720
rect 27755 18717 27767 18751
rect 27709 18711 27767 18717
rect 27976 18711 27988 18757
rect 26881 18683 26939 18689
rect 26881 18649 26893 18683
rect 26927 18649 26939 18683
rect 26881 18643 26939 18649
rect 26973 18683 27031 18689
rect 26973 18649 26985 18683
rect 27019 18649 27031 18683
rect 27724 18680 27752 18711
rect 27982 18708 27988 18711
rect 28040 18708 28046 18760
rect 28902 18680 28908 18692
rect 27724 18652 28908 18680
rect 26973 18643 27031 18649
rect 26108 18584 26556 18612
rect 26108 18572 26114 18584
rect 26694 18572 26700 18624
rect 26752 18612 26758 18624
rect 26988 18612 27016 18643
rect 28902 18640 28908 18652
rect 28960 18640 28966 18692
rect 26752 18584 27016 18612
rect 26752 18572 26758 18584
rect 27246 18572 27252 18624
rect 27304 18572 27310 18624
rect 1104 18522 43884 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 43884 18522
rect 1104 18448 43884 18470
rect 3050 18368 3056 18420
rect 3108 18368 3114 18420
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 4890 18368 4896 18420
rect 4948 18368 4954 18420
rect 5074 18368 5080 18420
rect 5132 18368 5138 18420
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 5721 18411 5779 18417
rect 5721 18408 5733 18411
rect 5684 18380 5733 18408
rect 5684 18368 5690 18380
rect 5721 18377 5733 18380
rect 5767 18408 5779 18411
rect 5994 18408 6000 18420
rect 5767 18380 6000 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 7107 18411 7165 18417
rect 6380 18380 7052 18408
rect 2590 18300 2596 18352
rect 2648 18340 2654 18352
rect 4798 18340 4804 18352
rect 2648 18312 4804 18340
rect 2648 18300 2654 18312
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1762 18272 1768 18284
rect 1719 18244 1768 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 1940 18275 1998 18281
rect 1940 18241 1952 18275
rect 1986 18272 1998 18275
rect 3234 18272 3240 18284
rect 1986 18244 3240 18272
rect 1986 18241 1998 18244
rect 1940 18235 1998 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 5092 18281 5120 18368
rect 6380 18352 6408 18380
rect 5902 18300 5908 18352
rect 5960 18340 5966 18352
rect 6362 18340 6368 18352
rect 5960 18312 6368 18340
rect 5960 18300 5966 18312
rect 6362 18300 6368 18312
rect 6420 18300 6426 18352
rect 6914 18300 6920 18352
rect 6972 18300 6978 18352
rect 7024 18349 7052 18380
rect 7107 18377 7119 18411
rect 7153 18408 7165 18411
rect 7374 18408 7380 18420
rect 7153 18380 7380 18408
rect 7153 18377 7165 18380
rect 7107 18371 7165 18377
rect 7374 18368 7380 18380
rect 7432 18408 7438 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 7432 18380 7849 18408
rect 7432 18368 7438 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 7926 18368 7932 18420
rect 7984 18368 7990 18420
rect 8478 18368 8484 18420
rect 8536 18368 8542 18420
rect 8573 18411 8631 18417
rect 8573 18377 8585 18411
rect 8619 18408 8631 18411
rect 9030 18408 9036 18420
rect 8619 18380 8800 18408
rect 8619 18377 8631 18380
rect 8573 18371 8631 18377
rect 7009 18343 7067 18349
rect 7009 18309 7021 18343
rect 7055 18309 7067 18343
rect 7009 18303 7067 18309
rect 7193 18343 7251 18349
rect 7193 18309 7205 18343
rect 7239 18309 7251 18343
rect 8202 18340 8208 18352
rect 7193 18303 7251 18309
rect 7392 18312 8208 18340
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5810 18272 5816 18284
rect 5077 18235 5135 18241
rect 5276 18244 5816 18272
rect 3694 18164 3700 18216
rect 3752 18204 3758 18216
rect 3789 18207 3847 18213
rect 3789 18204 3801 18207
rect 3752 18176 3801 18204
rect 3752 18164 3758 18176
rect 3789 18173 3801 18176
rect 3835 18204 3847 18207
rect 3878 18204 3884 18216
rect 3835 18176 3884 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18204 4399 18207
rect 4614 18204 4620 18216
rect 4387 18176 4620 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 5276 18136 5304 18244
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 6012 18204 6040 18235
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6144 18244 6745 18272
rect 6144 18232 6150 18244
rect 6733 18241 6745 18244
rect 6779 18272 6791 18275
rect 6932 18272 6960 18300
rect 6779 18244 6960 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5500 18176 6377 18204
rect 5500 18164 5506 18176
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 6454 18164 6460 18216
rect 6512 18204 6518 18216
rect 6549 18207 6607 18213
rect 6549 18204 6561 18207
rect 6512 18176 6561 18204
rect 6512 18164 6518 18176
rect 6549 18173 6561 18176
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 3896 18108 5304 18136
rect 3896 18080 3924 18108
rect 5902 18096 5908 18148
rect 5960 18136 5966 18148
rect 6656 18136 6684 18167
rect 6822 18164 6828 18216
rect 6880 18164 6886 18216
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7208 18204 7236 18303
rect 7282 18232 7288 18284
rect 7340 18232 7346 18284
rect 7392 18281 7420 18312
rect 8202 18300 8208 18312
rect 8260 18300 8266 18352
rect 8496 18340 8524 18368
rect 8496 18312 8616 18340
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 6972 18176 7236 18204
rect 6972 18164 6978 18176
rect 5960 18108 6684 18136
rect 5960 18096 5966 18108
rect 6730 18096 6736 18148
rect 6788 18136 6794 18148
rect 7392 18136 7420 18235
rect 7558 18232 7564 18284
rect 7616 18232 7622 18284
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 8386 18272 8392 18284
rect 8444 18281 8450 18284
rect 8351 18244 8392 18272
rect 7745 18235 7803 18241
rect 7760 18204 7788 18235
rect 8386 18232 8392 18244
rect 8444 18235 8451 18281
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8444 18232 8450 18235
rect 6788 18108 7420 18136
rect 7576 18176 7788 18204
rect 6788 18096 6794 18108
rect 3142 18028 3148 18080
rect 3200 18028 3206 18080
rect 3878 18028 3884 18080
rect 3936 18028 3942 18080
rect 4706 18028 4712 18080
rect 4764 18068 4770 18080
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 4764 18040 6193 18068
rect 4764 18028 4770 18040
rect 6181 18037 6193 18040
rect 6227 18068 6239 18071
rect 7190 18068 7196 18080
rect 6227 18040 7196 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7469 18071 7527 18077
rect 7469 18068 7481 18071
rect 7340 18040 7481 18068
rect 7340 18028 7346 18040
rect 7469 18037 7481 18040
rect 7515 18068 7527 18071
rect 7576 18068 7604 18176
rect 8110 18164 8116 18216
rect 8168 18164 8174 18216
rect 8496 18136 8524 18235
rect 8588 18204 8616 18312
rect 8772 18272 8800 18380
rect 8864 18380 9036 18408
rect 8864 18349 8892 18380
rect 9030 18368 9036 18380
rect 9088 18408 9094 18420
rect 9950 18408 9956 18420
rect 9088 18380 9956 18408
rect 9088 18368 9094 18380
rect 9784 18349 9812 18380
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10060 18380 10732 18408
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18309 8907 18343
rect 9769 18343 9827 18349
rect 8849 18303 8907 18309
rect 9140 18312 9674 18340
rect 9140 18281 9168 18312
rect 9646 18284 9674 18312
rect 9769 18309 9781 18343
rect 9815 18309 9827 18343
rect 10060 18340 10088 18380
rect 10594 18340 10600 18352
rect 9769 18303 9827 18309
rect 9876 18312 10088 18340
rect 9033 18275 9091 18281
rect 8772 18244 8984 18272
rect 8588 18176 8708 18204
rect 8680 18145 8708 18176
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 8665 18139 8723 18145
rect 8496 18108 8616 18136
rect 7515 18040 7604 18068
rect 7515 18037 7527 18040
rect 7469 18031 7527 18037
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7800 18040 7849 18068
rect 7800 18028 7806 18040
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 8588 18068 8616 18108
rect 8665 18105 8677 18139
rect 8711 18105 8723 18139
rect 8846 18136 8852 18148
rect 8665 18099 8723 18105
rect 8772 18108 8852 18136
rect 8772 18068 8800 18108
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 8588 18040 8800 18068
rect 8956 18068 8984 18244
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18241 9183 18275
rect 9125 18235 9183 18241
rect 9048 18136 9076 18235
rect 9214 18232 9220 18284
rect 9272 18232 9278 18284
rect 9398 18232 9404 18284
rect 9456 18232 9462 18284
rect 9582 18232 9588 18284
rect 9640 18272 9674 18284
rect 9876 18272 9904 18312
rect 9640 18244 9904 18272
rect 9640 18232 9646 18244
rect 9950 18232 9956 18284
rect 10008 18232 10014 18284
rect 10060 18281 10088 18312
rect 10336 18312 10600 18340
rect 10336 18281 10364 18312
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 10704 18340 10732 18380
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11333 18411 11391 18417
rect 11333 18408 11345 18411
rect 11020 18380 11345 18408
rect 11020 18368 11026 18380
rect 11333 18377 11345 18380
rect 11379 18408 11391 18411
rect 12802 18408 12808 18420
rect 11379 18380 12808 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13173 18411 13231 18417
rect 13173 18408 13185 18411
rect 13044 18380 13185 18408
rect 13044 18368 13050 18380
rect 13173 18377 13185 18380
rect 13219 18377 13231 18411
rect 13173 18371 13231 18377
rect 13538 18368 13544 18420
rect 13596 18368 13602 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 13814 18408 13820 18420
rect 13771 18380 13820 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 14550 18368 14556 18420
rect 14608 18368 14614 18420
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 15930 18408 15936 18420
rect 14792 18380 15936 18408
rect 14792 18368 14798 18380
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16482 18368 16488 18420
rect 16540 18368 16546 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 16724 18380 16957 18408
rect 16724 18368 16730 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 17954 18408 17960 18420
rect 16945 18371 17003 18377
rect 17052 18380 17960 18408
rect 11146 18340 11152 18352
rect 10704 18312 11152 18340
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 11974 18340 11980 18352
rect 11256 18312 11980 18340
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 9232 18204 9260 18232
rect 10152 18204 10180 18235
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 11256 18272 11284 18312
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 12115 18343 12173 18349
rect 12115 18309 12127 18343
rect 12161 18340 12173 18343
rect 12618 18340 12624 18352
rect 12161 18312 12624 18340
rect 12161 18309 12173 18312
rect 12115 18303 12173 18309
rect 12618 18300 12624 18312
rect 12676 18300 12682 18352
rect 13556 18340 13584 18368
rect 14568 18340 14596 18368
rect 16574 18340 16580 18352
rect 13004 18312 13400 18340
rect 13556 18312 14228 18340
rect 10468 18244 11284 18272
rect 10468 18232 10474 18244
rect 11790 18232 11796 18284
rect 11848 18232 11854 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 11931 18244 12388 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 11698 18204 11704 18216
rect 9232 18176 11704 18204
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 9214 18136 9220 18148
rect 9048 18108 9220 18136
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 10410 18136 10416 18148
rect 9815 18108 10416 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10410 18096 10416 18108
rect 10468 18096 10474 18148
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 11514 18136 11520 18148
rect 10928 18108 11520 18136
rect 10928 18096 10934 18108
rect 11514 18096 11520 18108
rect 11572 18136 11578 18148
rect 11900 18136 11928 18235
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 12360 18213 12388 18244
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 13004 18281 13032 18312
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18173 12679 18207
rect 12621 18167 12679 18173
rect 11572 18108 11928 18136
rect 12636 18136 12664 18167
rect 12710 18164 12716 18216
rect 12768 18164 12774 18216
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 13170 18204 13176 18216
rect 12851 18176 13176 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13280 18136 13308 18232
rect 13372 18204 13400 18312
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 13504 18244 13553 18272
rect 13504 18232 13510 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18272 13875 18275
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13863 18244 13921 18272
rect 13863 18241 13875 18244
rect 13817 18235 13875 18241
rect 13909 18241 13921 18244
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 14200 18281 14228 18312
rect 14384 18312 14596 18340
rect 15580 18312 16580 18340
rect 14384 18281 14412 18312
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18272 14611 18275
rect 14642 18272 14648 18284
rect 14599 18244 14648 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 14016 18204 14044 18232
rect 13372 18176 14044 18204
rect 13446 18136 13452 18148
rect 12636 18108 13032 18136
rect 13280 18108 13452 18136
rect 11572 18096 11578 18108
rect 9030 18068 9036 18080
rect 8956 18040 9036 18068
rect 7837 18031 7895 18037
rect 9030 18028 9036 18040
rect 9088 18028 9094 18080
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 9180 18040 9321 18068
rect 9180 18028 9186 18040
rect 9309 18037 9321 18040
rect 9355 18037 9367 18071
rect 9309 18031 9367 18037
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 11606 18028 11612 18080
rect 11664 18028 11670 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12894 18068 12900 18080
rect 12032 18040 12900 18068
rect 12032 18028 12038 18040
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13004 18077 13032 18108
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 13722 18096 13728 18148
rect 13780 18136 13786 18148
rect 14108 18136 14136 18235
rect 14274 18164 14280 18216
rect 14332 18204 14338 18216
rect 14476 18204 14504 18235
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 14332 18176 14504 18204
rect 14332 18164 14338 18176
rect 13780 18108 14136 18136
rect 13780 18096 13786 18108
rect 14016 18080 14044 18108
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 14752 18136 14780 18235
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15010 18272 15016 18284
rect 14967 18244 15016 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 15286 18232 15292 18284
rect 15344 18232 15350 18284
rect 15580 18281 15608 18312
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 17052 18340 17080 18380
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18693 18411 18751 18417
rect 18693 18408 18705 18411
rect 18380 18380 18705 18408
rect 18380 18368 18386 18380
rect 18693 18377 18705 18380
rect 18739 18377 18751 18411
rect 18693 18371 18751 18377
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 18840 18380 19840 18408
rect 18840 18368 18846 18380
rect 18340 18340 18368 18368
rect 19426 18340 19432 18352
rect 16960 18312 17080 18340
rect 17604 18312 18368 18340
rect 18892 18312 19432 18340
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16960 18281 16988 18312
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 15896 18244 16129 18272
rect 15896 18232 15902 18244
rect 16117 18241 16129 18244
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 16301 18275 16359 18281
rect 16301 18241 16313 18275
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16945 18275 17003 18281
rect 16945 18241 16957 18275
rect 16991 18241 17003 18275
rect 16945 18235 17003 18241
rect 15028 18204 15056 18232
rect 15470 18204 15476 18216
rect 15028 18176 15476 18204
rect 15470 18164 15476 18176
rect 15528 18204 15534 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 15528 18176 15761 18204
rect 15528 18164 15534 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16316 18204 16344 18235
rect 17126 18232 17132 18284
rect 17184 18232 17190 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17494 18272 17500 18284
rect 17359 18244 17500 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17604 18281 17632 18312
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18241 17647 18275
rect 17589 18235 17647 18241
rect 17678 18232 17684 18284
rect 17736 18272 17742 18284
rect 17865 18275 17923 18281
rect 17865 18272 17877 18275
rect 17736 18244 17877 18272
rect 17736 18232 17742 18244
rect 17865 18241 17877 18244
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18272 18015 18275
rect 18046 18272 18052 18284
rect 18003 18244 18052 18272
rect 18003 18241 18015 18244
rect 17957 18235 18015 18241
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 18892 18281 18920 18312
rect 19426 18300 19432 18312
rect 19484 18340 19490 18352
rect 19702 18340 19708 18352
rect 19484 18312 19708 18340
rect 19484 18300 19490 18312
rect 19702 18300 19708 18312
rect 19760 18300 19766 18352
rect 19812 18340 19840 18380
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 20438 18408 20444 18420
rect 19944 18380 20444 18408
rect 19944 18368 19950 18380
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 20898 18368 20904 18420
rect 20956 18368 20962 18420
rect 21085 18411 21143 18417
rect 21085 18377 21097 18411
rect 21131 18408 21143 18411
rect 21174 18408 21180 18420
rect 21131 18380 21180 18408
rect 21131 18377 21143 18380
rect 21085 18371 21143 18377
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 21358 18368 21364 18420
rect 21416 18368 21422 18420
rect 23845 18411 23903 18417
rect 23845 18408 23857 18411
rect 21652 18380 23857 18408
rect 21376 18340 21404 18368
rect 19812 18312 21404 18340
rect 18877 18275 18935 18281
rect 18248 18244 18552 18272
rect 18248 18238 18276 18244
rect 16080 18176 16344 18204
rect 16080 18164 16086 18176
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 18156 18210 18276 18238
rect 18156 18204 18184 18210
rect 17460 18176 18184 18204
rect 18417 18207 18475 18213
rect 17460 18164 17466 18176
rect 18417 18173 18429 18207
rect 18463 18173 18475 18207
rect 18524 18204 18552 18244
rect 18877 18241 18889 18275
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 19150 18232 19156 18284
rect 19208 18232 19214 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 19978 18272 19984 18284
rect 19935 18244 19984 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20680 18244 20821 18272
rect 20680 18232 20686 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20956 18244 21005 18272
rect 20956 18232 20962 18244
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21361 18275 21419 18281
rect 21361 18241 21373 18275
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 18524 18176 19349 18204
rect 18417 18167 18475 18173
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 14918 18136 14924 18148
rect 14700 18108 14924 18136
rect 14700 18096 14706 18108
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 15381 18139 15439 18145
rect 15381 18136 15393 18139
rect 15344 18108 15393 18136
rect 15344 18096 15350 18108
rect 15381 18105 15393 18108
rect 15427 18105 15439 18139
rect 17034 18136 17040 18148
rect 15381 18099 15439 18105
rect 16408 18108 17040 18136
rect 12989 18071 13047 18077
rect 12989 18037 13001 18071
rect 13035 18068 13047 18071
rect 13078 18068 13084 18080
rect 13035 18040 13084 18068
rect 13035 18037 13047 18040
rect 12989 18031 13047 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13357 18071 13415 18077
rect 13357 18037 13369 18071
rect 13403 18068 13415 18071
rect 13538 18068 13544 18080
rect 13403 18040 13544 18068
rect 13403 18037 13415 18040
rect 13357 18031 13415 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13998 18028 14004 18080
rect 14056 18028 14062 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14550 18068 14556 18080
rect 14424 18040 14556 18068
rect 14424 18028 14430 18040
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 16408 18068 16436 18108
rect 17034 18096 17040 18108
rect 17092 18096 17098 18148
rect 17586 18096 17592 18148
rect 17644 18096 17650 18148
rect 18046 18096 18052 18148
rect 18104 18136 18110 18148
rect 18432 18136 18460 18167
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 20916 18204 20944 18232
rect 20496 18176 20944 18204
rect 20496 18164 20502 18176
rect 18598 18136 18604 18148
rect 18104 18108 18604 18136
rect 18104 18096 18110 18108
rect 18598 18096 18604 18108
rect 18656 18096 18662 18148
rect 18969 18139 19027 18145
rect 18969 18105 18981 18139
rect 19015 18136 19027 18139
rect 20162 18136 20168 18148
rect 19015 18108 20168 18136
rect 19015 18105 19027 18108
rect 18969 18099 19027 18105
rect 20162 18096 20168 18108
rect 20220 18136 20226 18148
rect 20714 18136 20720 18148
rect 20220 18108 20720 18136
rect 20220 18096 20226 18108
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 21284 18136 21312 18235
rect 21376 18204 21404 18235
rect 21542 18232 21548 18284
rect 21600 18232 21606 18284
rect 21652 18281 21680 18380
rect 23845 18377 23857 18380
rect 23891 18377 23903 18411
rect 23845 18371 23903 18377
rect 24118 18368 24124 18420
rect 24176 18408 24182 18420
rect 24673 18411 24731 18417
rect 24176 18380 24348 18408
rect 24176 18368 24182 18380
rect 22097 18343 22155 18349
rect 22097 18340 22109 18343
rect 21836 18312 22109 18340
rect 21836 18284 21864 18312
rect 22097 18309 22109 18312
rect 22143 18309 22155 18343
rect 22097 18303 22155 18309
rect 22646 18300 22652 18352
rect 22704 18300 22710 18352
rect 23290 18300 23296 18352
rect 23348 18340 23354 18352
rect 24320 18349 24348 18380
rect 24673 18377 24685 18411
rect 24719 18408 24731 18411
rect 25222 18408 25228 18420
rect 24719 18380 25228 18408
rect 24719 18377 24731 18380
rect 24673 18371 24731 18377
rect 25222 18368 25228 18380
rect 25280 18368 25286 18420
rect 25317 18411 25375 18417
rect 25317 18377 25329 18411
rect 25363 18408 25375 18411
rect 25406 18408 25412 18420
rect 25363 18380 25412 18408
rect 25363 18377 25375 18380
rect 25317 18371 25375 18377
rect 25406 18368 25412 18380
rect 25464 18408 25470 18420
rect 26050 18408 26056 18420
rect 25464 18380 26056 18408
rect 25464 18368 25470 18380
rect 26050 18368 26056 18380
rect 26108 18368 26114 18420
rect 26329 18411 26387 18417
rect 26329 18377 26341 18411
rect 26375 18408 26387 18411
rect 26418 18408 26424 18420
rect 26375 18380 26424 18408
rect 26375 18377 26387 18380
rect 26329 18371 26387 18377
rect 26418 18368 26424 18380
rect 26476 18368 26482 18420
rect 28074 18408 28080 18420
rect 27172 18380 28080 18408
rect 23385 18343 23443 18349
rect 23385 18340 23397 18343
rect 23348 18312 23397 18340
rect 23348 18300 23354 18312
rect 23385 18309 23397 18312
rect 23431 18309 23443 18343
rect 23385 18303 23443 18309
rect 24305 18343 24363 18349
rect 24305 18309 24317 18343
rect 24351 18309 24363 18343
rect 27172 18340 27200 18380
rect 28074 18368 28080 18380
rect 28132 18368 28138 18420
rect 24305 18303 24363 18309
rect 24412 18312 24808 18340
rect 21637 18275 21695 18281
rect 21637 18241 21649 18275
rect 21683 18241 21695 18275
rect 21637 18235 21695 18241
rect 21818 18232 21824 18284
rect 21876 18232 21882 18284
rect 21910 18232 21916 18284
rect 21968 18232 21974 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22020 18244 22201 18272
rect 21928 18204 21956 18232
rect 21376 18176 21956 18204
rect 21726 18136 21732 18148
rect 21284 18108 21732 18136
rect 21726 18096 21732 18108
rect 21784 18136 21790 18148
rect 22020 18136 22048 18244
rect 22189 18241 22201 18244
rect 22235 18272 22247 18275
rect 22833 18275 22891 18281
rect 22833 18272 22845 18275
rect 22235 18244 22845 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22833 18241 22845 18244
rect 22879 18272 22891 18275
rect 23934 18272 23940 18284
rect 22879 18244 23940 18272
rect 22879 18241 22891 18244
rect 22833 18235 22891 18241
rect 23934 18232 23940 18244
rect 23992 18232 23998 18284
rect 24118 18232 24124 18284
rect 24176 18232 24182 18284
rect 22462 18164 22468 18216
rect 22520 18204 22526 18216
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22520 18176 22753 18204
rect 22520 18164 22526 18176
rect 22741 18173 22753 18176
rect 22787 18204 22799 18207
rect 22922 18204 22928 18216
rect 22787 18176 22928 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23293 18207 23351 18213
rect 23293 18204 23305 18207
rect 23072 18176 23305 18204
rect 23072 18164 23078 18176
rect 23293 18173 23305 18176
rect 23339 18204 23351 18207
rect 24320 18204 24348 18303
rect 24412 18284 24440 18312
rect 24394 18232 24400 18284
rect 24452 18232 24458 18284
rect 24489 18275 24547 18281
rect 24489 18241 24501 18275
rect 24535 18272 24547 18275
rect 24670 18272 24676 18284
rect 24535 18244 24676 18272
rect 24535 18241 24547 18244
rect 24489 18235 24547 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 24780 18281 24808 18312
rect 25056 18312 25452 18340
rect 25056 18281 25084 18312
rect 25424 18284 25452 18312
rect 25516 18312 27200 18340
rect 27240 18343 27298 18349
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18241 24823 18275
rect 24765 18235 24823 18241
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18241 25007 18275
rect 24949 18235 25007 18241
rect 25041 18275 25099 18281
rect 25041 18241 25053 18275
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 24578 18204 24584 18216
rect 23339 18176 24072 18204
rect 24320 18176 24584 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 21784 18108 22048 18136
rect 23753 18139 23811 18145
rect 21784 18096 21790 18108
rect 23753 18105 23765 18139
rect 23799 18105 23811 18139
rect 24044 18136 24072 18176
rect 24578 18164 24584 18176
rect 24636 18204 24642 18216
rect 24964 18204 24992 18235
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 25406 18232 25412 18284
rect 25464 18232 25470 18284
rect 25516 18281 25544 18312
rect 27240 18309 27252 18343
rect 27286 18340 27298 18343
rect 28166 18340 28172 18352
rect 27286 18312 28172 18340
rect 27286 18309 27298 18312
rect 27240 18303 27298 18309
rect 28166 18300 28172 18312
rect 28224 18300 28230 18352
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 26513 18275 26571 18281
rect 26513 18272 26525 18275
rect 25648 18244 26525 18272
rect 25648 18232 25654 18244
rect 26513 18241 26525 18244
rect 26559 18241 26571 18275
rect 27614 18272 27620 18284
rect 26513 18235 26571 18241
rect 26988 18244 27620 18272
rect 24636 18176 24992 18204
rect 24636 18164 24642 18176
rect 25682 18164 25688 18216
rect 25740 18204 25746 18216
rect 26789 18207 26847 18213
rect 26789 18204 26801 18207
rect 25740 18176 26801 18204
rect 25740 18164 25746 18176
rect 26789 18173 26801 18176
rect 26835 18173 26847 18207
rect 26789 18167 26847 18173
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 26988 18213 27016 18244
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26936 18176 26985 18204
rect 26936 18164 26942 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 24044 18108 24440 18136
rect 23753 18099 23811 18105
rect 15151 18040 16436 18068
rect 18325 18071 18383 18077
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 18325 18037 18337 18071
rect 18371 18068 18383 18071
rect 18506 18068 18512 18080
rect 18371 18040 18512 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 19794 18068 19800 18080
rect 18748 18040 19800 18068
rect 18748 18028 18754 18040
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18068 21971 18071
rect 22002 18068 22008 18080
rect 21959 18040 22008 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 23768 18068 23796 18099
rect 24026 18068 24032 18080
rect 23768 18040 24032 18068
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 24412 18068 24440 18108
rect 24486 18096 24492 18148
rect 24544 18136 24550 18148
rect 24544 18108 26234 18136
rect 24544 18096 24550 18108
rect 25038 18068 25044 18080
rect 24412 18040 25044 18068
rect 25038 18028 25044 18040
rect 25096 18028 25102 18080
rect 26050 18028 26056 18080
rect 26108 18028 26114 18080
rect 26206 18068 26234 18108
rect 26694 18096 26700 18148
rect 26752 18096 26758 18148
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 26206 18040 28365 18068
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 28353 18031 28411 18037
rect 1104 17978 43884 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 43884 17978
rect 1104 17904 43884 17926
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 3605 17867 3663 17873
rect 3605 17864 3617 17867
rect 3568 17836 3617 17864
rect 3568 17824 3574 17836
rect 3605 17833 3617 17836
rect 3651 17833 3663 17867
rect 3605 17827 3663 17833
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4614 17864 4620 17876
rect 4387 17836 4620 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5534 17864 5540 17876
rect 4816 17836 5540 17864
rect 4816 17796 4844 17836
rect 5534 17824 5540 17836
rect 5592 17864 5598 17876
rect 5592 17836 6684 17864
rect 5592 17824 5598 17836
rect 6656 17808 6684 17836
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6880 17836 7113 17864
rect 6880 17824 6886 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7926 17864 7932 17876
rect 7101 17827 7159 17833
rect 7484 17836 7932 17864
rect 2746 17768 4844 17796
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 1857 17731 1915 17737
rect 1857 17728 1869 17731
rect 1268 17700 1869 17728
rect 1268 17688 1274 17700
rect 1857 17697 1869 17700
rect 1903 17697 1915 17731
rect 1857 17691 1915 17697
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 1596 17592 1624 17623
rect 1670 17620 1676 17672
rect 1728 17660 1734 17672
rect 2746 17660 2774 17768
rect 2958 17688 2964 17740
rect 3016 17688 3022 17740
rect 3602 17728 3608 17740
rect 3068 17700 3608 17728
rect 1728 17632 2774 17660
rect 1728 17620 1734 17632
rect 3068 17592 3096 17700
rect 3602 17688 3608 17700
rect 3660 17688 3666 17740
rect 4614 17688 4620 17740
rect 4672 17688 4678 17740
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3936 17632 4077 17660
rect 3936 17620 3942 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4430 17660 4436 17672
rect 4295 17632 4436 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 4525 17663 4583 17669
rect 4525 17629 4537 17663
rect 4571 17660 4583 17663
rect 4632 17660 4660 17688
rect 4724 17669 4752 17768
rect 5810 17756 5816 17808
rect 5868 17796 5874 17808
rect 6454 17796 6460 17808
rect 5868 17768 6460 17796
rect 5868 17756 5874 17768
rect 6454 17756 6460 17768
rect 6512 17756 6518 17808
rect 6638 17756 6644 17808
rect 6696 17756 6702 17808
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 5077 17731 5135 17737
rect 5077 17728 5089 17731
rect 4856 17700 5089 17728
rect 4856 17688 4862 17700
rect 5077 17697 5089 17700
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 5626 17688 5632 17740
rect 5684 17688 5690 17740
rect 6181 17731 6239 17737
rect 6181 17697 6193 17731
rect 6227 17728 6239 17731
rect 6840 17728 6868 17824
rect 6227 17700 6868 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 7374 17688 7380 17740
rect 7432 17688 7438 17740
rect 7484 17737 7512 17836
rect 7926 17824 7932 17836
rect 7984 17864 7990 17876
rect 8665 17867 8723 17873
rect 8665 17864 8677 17867
rect 7984 17836 8677 17864
rect 7984 17824 7990 17836
rect 8665 17833 8677 17836
rect 8711 17833 8723 17867
rect 8665 17827 8723 17833
rect 8754 17824 8760 17876
rect 8812 17864 8818 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 8812 17836 9444 17864
rect 8812 17824 8818 17836
rect 8110 17796 8116 17808
rect 7576 17768 8116 17796
rect 7576 17737 7604 17768
rect 8110 17756 8116 17768
rect 8168 17796 8174 17808
rect 8941 17799 8999 17805
rect 8941 17796 8953 17799
rect 8168 17768 8953 17796
rect 8168 17756 8174 17768
rect 8941 17765 8953 17768
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 9030 17756 9036 17808
rect 9088 17796 9094 17808
rect 9088 17768 9352 17796
rect 9088 17756 9094 17768
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17697 7527 17731
rect 7469 17691 7527 17697
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8352 17700 8616 17728
rect 8352 17688 8358 17700
rect 4571 17632 4660 17660
rect 4709 17663 4767 17669
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5644 17660 5672 17688
rect 5031 17632 5672 17660
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 5902 17620 5908 17672
rect 5960 17620 5966 17672
rect 6086 17660 6092 17672
rect 6012 17632 6092 17660
rect 1596 17564 3096 17592
rect 3436 17524 3464 17620
rect 4157 17595 4215 17601
rect 4157 17561 4169 17595
rect 4203 17592 4215 17595
rect 4617 17595 4675 17601
rect 4617 17592 4629 17595
rect 4203 17564 4629 17592
rect 4203 17561 4215 17564
rect 4157 17555 4215 17561
rect 4617 17561 4629 17564
rect 4663 17561 4675 17595
rect 4617 17555 4675 17561
rect 4827 17595 4885 17601
rect 4827 17561 4839 17595
rect 4873 17561 4885 17595
rect 4827 17555 4885 17561
rect 4842 17524 4870 17555
rect 5718 17552 5724 17604
rect 5776 17552 5782 17604
rect 5626 17524 5632 17536
rect 3436 17496 5632 17524
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 6012 17533 6040 17632
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 7834 17620 7840 17672
rect 7892 17620 7898 17672
rect 8588 17669 8616 17700
rect 8846 17688 8852 17740
rect 8904 17728 8910 17740
rect 9324 17737 9352 17768
rect 9416 17737 9444 17836
rect 9876 17836 11069 17864
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 8904 17700 9229 17728
rect 8904 17688 8910 17700
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 9309 17731 9367 17737
rect 9309 17697 9321 17731
rect 9355 17697 9367 17731
rect 9309 17691 9367 17697
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 6638 17552 6644 17604
rect 6696 17592 6702 17604
rect 6696 17564 7696 17592
rect 6696 17552 6702 17564
rect 5997 17527 6055 17533
rect 5997 17493 6009 17527
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6086 17484 6092 17536
rect 6144 17484 6150 17536
rect 6546 17484 6552 17536
rect 6604 17524 6610 17536
rect 6917 17527 6975 17533
rect 6917 17524 6929 17527
rect 6604 17496 6929 17524
rect 6604 17484 6610 17496
rect 6917 17493 6929 17496
rect 6963 17493 6975 17527
rect 7668 17524 7696 17564
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 8772 17592 8800 17623
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 7800 17564 8800 17592
rect 9416 17592 9444 17691
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17659 9827 17663
rect 9876 17659 9904 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13504 17836 13921 17864
rect 13504 17824 13510 17836
rect 13909 17833 13921 17836
rect 13955 17833 13967 17867
rect 13909 17827 13967 17833
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14274 17864 14280 17876
rect 14231 17836 14280 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14384 17836 16988 17864
rect 10226 17756 10232 17808
rect 10284 17796 10290 17808
rect 10284 17768 11192 17796
rect 10284 17756 10290 17768
rect 10520 17737 10548 17768
rect 10505 17731 10563 17737
rect 9968 17700 10364 17728
rect 9968 17669 9996 17700
rect 10336 17672 10364 17700
rect 10505 17697 10517 17731
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 10870 17688 10876 17740
rect 10928 17688 10934 17740
rect 9815 17631 9904 17659
rect 9953 17663 10011 17669
rect 9815 17629 9827 17631
rect 9769 17623 9827 17629
rect 9953 17629 9965 17663
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10226 17620 10232 17672
rect 10284 17620 10290 17672
rect 10318 17620 10324 17672
rect 10376 17620 10382 17672
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10468 17632 10609 17660
rect 10468 17620 10474 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 10888 17660 10916 17688
rect 10827 17632 10916 17660
rect 10965 17663 11023 17669
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 10965 17629 10977 17663
rect 11011 17659 11023 17663
rect 11164 17660 11192 17768
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 14384 17796 14412 17836
rect 16960 17808 16988 17836
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 17092 17836 17233 17864
rect 17092 17824 17098 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17221 17827 17279 17833
rect 17954 17824 17960 17876
rect 18012 17824 18018 17876
rect 18506 17824 18512 17876
rect 18564 17824 18570 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 19116 17836 20637 17864
rect 19116 17824 19122 17836
rect 20625 17833 20637 17836
rect 20671 17833 20683 17867
rect 20625 17827 20683 17833
rect 21174 17824 21180 17876
rect 21232 17824 21238 17876
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 22554 17864 22560 17876
rect 21600 17836 22560 17864
rect 21600 17824 21606 17836
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 23198 17864 23204 17876
rect 23155 17836 23204 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 23308 17836 23520 17864
rect 15286 17796 15292 17808
rect 13596 17768 14412 17796
rect 14568 17768 15292 17796
rect 13596 17756 13602 17768
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11514 17728 11520 17740
rect 11379 17700 11520 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 11664 17700 11713 17728
rect 11664 17688 11670 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13354 17728 13360 17740
rect 12860 17700 13360 17728
rect 12860 17688 12866 17700
rect 13354 17688 13360 17700
rect 13412 17728 13418 17740
rect 13412 17700 14142 17728
rect 13412 17688 13418 17700
rect 11072 17659 11192 17660
rect 11011 17632 11192 17659
rect 11011 17631 11100 17632
rect 11011 17629 11023 17631
rect 10965 17623 11023 17629
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9416 17564 9873 17592
rect 7800 17552 7806 17564
rect 9861 17561 9873 17564
rect 9907 17561 9919 17595
rect 9861 17555 9919 17561
rect 10091 17595 10149 17601
rect 10091 17561 10103 17595
rect 10137 17592 10149 17595
rect 10502 17592 10508 17604
rect 10137 17564 10508 17592
rect 10137 17561 10149 17564
rect 10091 17555 10149 17561
rect 7926 17524 7932 17536
rect 7668 17496 7932 17524
rect 6917 17487 6975 17493
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8444 17496 8493 17524
rect 8444 17484 8450 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 8481 17487 8539 17493
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 9398 17524 9404 17536
rect 8628 17496 9404 17524
rect 8628 17484 8634 17496
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9585 17527 9643 17533
rect 9585 17493 9597 17527
rect 9631 17524 9643 17527
rect 9766 17524 9772 17536
rect 9631 17496 9772 17524
rect 9631 17493 9643 17496
rect 9585 17487 9643 17493
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 9876 17524 9904 17555
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 9876 17496 10333 17524
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10612 17524 10640 17623
rect 10704 17592 10732 17623
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12713 17663 12771 17669
rect 12713 17660 12725 17663
rect 11940 17632 12725 17660
rect 11940 17620 11946 17632
rect 12713 17629 12725 17632
rect 12759 17660 12771 17663
rect 12894 17660 12900 17672
rect 12759 17632 12900 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 14114 17669 14142 17700
rect 14568 17669 14596 17768
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 15672 17768 16436 17796
rect 14642 17688 14648 17740
rect 14700 17688 14706 17740
rect 15672 17728 15700 17768
rect 14890 17700 15700 17728
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14660 17660 14688 17688
rect 14890 17672 14918 17700
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 16408 17737 16436 17768
rect 16942 17756 16948 17808
rect 17000 17756 17006 17808
rect 17586 17756 17592 17808
rect 17644 17756 17650 17808
rect 17972 17796 18000 17824
rect 23308 17808 23336 17836
rect 18690 17796 18696 17808
rect 17972 17768 18696 17796
rect 18690 17756 18696 17768
rect 18748 17756 18754 17808
rect 21637 17799 21695 17805
rect 21637 17796 21649 17799
rect 18800 17768 21649 17796
rect 16025 17731 16083 17737
rect 16025 17728 16037 17731
rect 15804 17700 16037 17728
rect 15804 17688 15810 17700
rect 16025 17697 16037 17700
rect 16071 17697 16083 17731
rect 16025 17691 16083 17697
rect 16393 17731 16451 17737
rect 16393 17697 16405 17731
rect 16439 17697 16451 17731
rect 16393 17691 16451 17697
rect 18046 17688 18052 17740
rect 18104 17688 18110 17740
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 18601 17731 18659 17737
rect 18601 17728 18613 17731
rect 18472 17700 18613 17728
rect 18472 17688 18478 17700
rect 18601 17697 18613 17700
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 14660 17632 14780 17660
rect 14553 17623 14611 17629
rect 10870 17592 10876 17604
rect 10704 17564 10876 17592
rect 10870 17552 10876 17564
rect 10928 17592 10934 17604
rect 13357 17595 13415 17601
rect 10928 17564 11192 17592
rect 10928 17552 10934 17564
rect 11164 17533 11192 17564
rect 13357 17561 13369 17595
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10612 17496 11069 17524
rect 10321 17487 10379 17493
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 12342 17484 12348 17536
rect 12400 17484 12406 17536
rect 13262 17484 13268 17536
rect 13320 17484 13326 17536
rect 13372 17524 13400 17555
rect 13630 17552 13636 17604
rect 13688 17552 13694 17604
rect 13725 17595 13783 17601
rect 13725 17561 13737 17595
rect 13771 17592 13783 17595
rect 14274 17592 14280 17604
rect 13771 17564 14280 17592
rect 13771 17561 13783 17564
rect 13725 17555 13783 17561
rect 14274 17552 14280 17564
rect 14332 17552 14338 17604
rect 14366 17552 14372 17604
rect 14424 17552 14430 17604
rect 14752 17601 14780 17632
rect 14826 17620 14832 17672
rect 14884 17669 14918 17672
rect 14884 17663 14933 17669
rect 14884 17629 14887 17663
rect 14921 17629 14933 17663
rect 14884 17623 14933 17629
rect 14884 17620 14890 17623
rect 15010 17620 15016 17672
rect 15068 17620 15074 17672
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15151 17632 15332 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 14645 17595 14703 17601
rect 14645 17561 14657 17595
rect 14691 17561 14703 17595
rect 14645 17555 14703 17561
rect 14737 17595 14795 17601
rect 14737 17561 14749 17595
rect 14783 17561 14795 17595
rect 15304 17592 15332 17632
rect 15378 17620 15384 17672
rect 15436 17620 15442 17672
rect 15470 17620 15476 17672
rect 15528 17660 15534 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 15528 17632 15577 17660
rect 15528 17620 15534 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 15856 17592 15884 17620
rect 15304 17564 15884 17592
rect 14737 17555 14795 17561
rect 14660 17524 14688 17555
rect 14918 17524 14924 17536
rect 13372 17496 14924 17524
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 15197 17527 15255 17533
rect 15197 17524 15209 17527
rect 15160 17496 15209 17524
rect 15160 17484 15166 17496
rect 15197 17493 15209 17496
rect 15243 17493 15255 17527
rect 15197 17487 15255 17493
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 15841 17527 15899 17533
rect 15841 17524 15853 17527
rect 15344 17496 15853 17524
rect 15344 17484 15350 17496
rect 15841 17493 15853 17496
rect 15887 17493 15899 17527
rect 16132 17524 16160 17623
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16761 17663 16819 17669
rect 16761 17660 16773 17663
rect 16632 17632 16773 17660
rect 16632 17620 16638 17632
rect 16761 17629 16773 17632
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17629 17095 17663
rect 17037 17623 17095 17629
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 16482 17552 16488 17604
rect 16540 17552 16546 17604
rect 16206 17524 16212 17536
rect 16132 17496 16212 17524
rect 15841 17487 15899 17493
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16356 17496 16589 17524
rect 16356 17484 16362 17496
rect 16577 17493 16589 17496
rect 16623 17493 16635 17527
rect 17052 17524 17080 17623
rect 17236 17592 17264 17623
rect 17310 17620 17316 17672
rect 17368 17620 17374 17672
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 17736 17632 18153 17660
rect 17736 17620 17742 17632
rect 18141 17629 18153 17632
rect 18187 17629 18199 17663
rect 18141 17623 18199 17629
rect 17586 17592 17592 17604
rect 17236 17564 17592 17592
rect 17586 17552 17592 17564
rect 17644 17592 17650 17604
rect 17644 17564 18092 17592
rect 17644 17552 17650 17564
rect 17494 17524 17500 17536
rect 17052 17496 17500 17524
rect 16577 17487 16635 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18064 17524 18092 17564
rect 18800 17524 18828 17768
rect 21637 17765 21649 17768
rect 21683 17765 21695 17799
rect 21637 17759 21695 17765
rect 21910 17756 21916 17808
rect 21968 17756 21974 17808
rect 22002 17756 22008 17808
rect 22060 17796 22066 17808
rect 22097 17799 22155 17805
rect 22097 17796 22109 17799
rect 22060 17768 22109 17796
rect 22060 17756 22066 17768
rect 22097 17765 22109 17768
rect 22143 17765 22155 17799
rect 22097 17759 22155 17765
rect 23290 17756 23296 17808
rect 23348 17756 23354 17808
rect 23492 17805 23520 17836
rect 24670 17824 24676 17876
rect 24728 17864 24734 17876
rect 25130 17864 25136 17876
rect 24728 17836 25136 17864
rect 24728 17824 24734 17836
rect 23477 17799 23535 17805
rect 23477 17765 23489 17799
rect 23523 17765 23535 17799
rect 23477 17759 23535 17765
rect 24029 17799 24087 17805
rect 24029 17765 24041 17799
rect 24075 17796 24087 17799
rect 24075 17768 24992 17796
rect 24075 17765 24087 17768
rect 24029 17759 24087 17765
rect 19245 17731 19303 17737
rect 19245 17697 19257 17731
rect 19291 17728 19303 17731
rect 19291 17700 20852 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 19518 17620 19524 17672
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19628 17592 19656 17623
rect 19702 17620 19708 17672
rect 19760 17620 19766 17672
rect 19794 17620 19800 17672
rect 19852 17660 19858 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19852 17632 19901 17660
rect 19852 17620 19858 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 19978 17620 19984 17672
rect 20036 17620 20042 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20824 17669 20852 17700
rect 21008 17700 21312 17728
rect 21008 17672 21036 17700
rect 20533 17663 20591 17669
rect 20128 17632 20392 17660
rect 20128 17620 20134 17632
rect 19484 17564 19656 17592
rect 19996 17592 20024 17620
rect 20257 17595 20315 17601
rect 20257 17592 20269 17595
rect 19996 17564 20269 17592
rect 19484 17552 19490 17564
rect 20257 17561 20269 17564
rect 20303 17561 20315 17595
rect 20257 17555 20315 17561
rect 18064 17496 18828 17524
rect 20364 17524 20392 17632
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 20548 17592 20576 17623
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 20714 17592 20720 17604
rect 20548 17564 20720 17592
rect 20714 17552 20720 17564
rect 20772 17592 20778 17604
rect 21100 17592 21128 17623
rect 21174 17620 21180 17672
rect 21232 17620 21238 17672
rect 21284 17660 21312 17700
rect 21358 17688 21364 17740
rect 21416 17688 21422 17740
rect 24044 17728 24072 17759
rect 21836 17700 24072 17728
rect 21450 17660 21456 17672
rect 21284 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 21836 17669 21864 17700
rect 24762 17688 24768 17740
rect 24820 17688 24826 17740
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 21968 17632 22293 17660
rect 21968 17620 21974 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 23106 17660 23112 17672
rect 22428 17632 23112 17660
rect 22428 17620 22434 17632
rect 23106 17620 23112 17632
rect 23164 17660 23170 17672
rect 23293 17663 23351 17669
rect 23293 17660 23305 17663
rect 23164 17632 23305 17660
rect 23164 17620 23170 17632
rect 23293 17629 23305 17632
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23474 17620 23480 17672
rect 23532 17657 23538 17672
rect 23569 17663 23627 17669
rect 23569 17657 23581 17663
rect 23532 17629 23581 17657
rect 23615 17629 23627 17663
rect 23532 17620 23538 17629
rect 23569 17623 23627 17629
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 24780 17660 24808 17688
rect 24964 17660 24992 17768
rect 25056 17737 25084 17836
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 25406 17824 25412 17876
rect 25464 17824 25470 17876
rect 25590 17824 25596 17876
rect 25648 17824 25654 17876
rect 25869 17867 25927 17873
rect 25869 17833 25881 17867
rect 25915 17864 25927 17867
rect 26142 17864 26148 17876
rect 25915 17836 26148 17864
rect 25915 17833 25927 17836
rect 25869 17827 25927 17833
rect 26142 17824 26148 17836
rect 26200 17824 26206 17876
rect 26786 17824 26792 17876
rect 26844 17824 26850 17876
rect 25608 17796 25636 17824
rect 25424 17768 25636 17796
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17728 25099 17731
rect 25424 17728 25452 17768
rect 26326 17728 26332 17740
rect 25087 17700 25452 17728
rect 25516 17700 26332 17728
rect 25087 17697 25099 17700
rect 25041 17691 25099 17697
rect 25314 17660 25320 17672
rect 24780 17632 24926 17660
rect 24964 17632 25320 17660
rect 21358 17592 21364 17604
rect 20772 17564 21364 17592
rect 20772 17552 20778 17564
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 22922 17552 22928 17604
rect 22980 17592 22986 17604
rect 22980 17564 23612 17592
rect 22980 17552 22986 17564
rect 20993 17527 21051 17533
rect 20993 17524 21005 17527
rect 20364 17496 21005 17524
rect 20993 17493 21005 17496
rect 21039 17524 21051 17527
rect 23382 17524 23388 17536
rect 21039 17496 23388 17524
rect 21039 17493 21051 17496
rect 20993 17487 21051 17493
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 23584 17524 23612 17564
rect 23658 17552 23664 17604
rect 23716 17592 23722 17604
rect 24486 17592 24492 17604
rect 23716 17564 24492 17592
rect 23716 17552 23722 17564
rect 24486 17552 24492 17564
rect 24544 17552 24550 17604
rect 24670 17552 24676 17604
rect 24728 17552 24734 17604
rect 24762 17552 24768 17604
rect 24820 17552 24826 17604
rect 24898 17601 24926 17632
rect 25314 17620 25320 17632
rect 25372 17620 25378 17672
rect 25516 17604 25544 17700
rect 26326 17688 26332 17700
rect 26384 17728 26390 17740
rect 26970 17728 26976 17740
rect 26384 17700 26976 17728
rect 26384 17688 26390 17700
rect 26970 17688 26976 17700
rect 27028 17688 27034 17740
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 26145 17663 26203 17669
rect 26145 17660 26157 17663
rect 25832 17632 26157 17660
rect 25832 17620 25838 17632
rect 26145 17629 26157 17632
rect 26191 17629 26203 17663
rect 26145 17623 26203 17629
rect 26421 17663 26479 17669
rect 26421 17629 26433 17663
rect 26467 17660 26479 17663
rect 27246 17660 27252 17672
rect 26467 17632 27252 17660
rect 26467 17629 26479 17632
rect 26421 17623 26479 17629
rect 27246 17620 27252 17632
rect 27304 17620 27310 17672
rect 27430 17620 27436 17672
rect 27488 17620 27494 17672
rect 24883 17595 24941 17601
rect 24883 17561 24895 17595
rect 24929 17561 24941 17595
rect 24883 17555 24941 17561
rect 25240 17564 25452 17592
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 23532 17496 24133 17524
rect 23532 17484 23538 17496
rect 24121 17493 24133 17496
rect 24167 17493 24179 17527
rect 24121 17487 24179 17493
rect 24397 17527 24455 17533
rect 24397 17493 24409 17527
rect 24443 17524 24455 17527
rect 25240 17524 25268 17564
rect 24443 17496 25268 17524
rect 25424 17524 25452 17564
rect 25498 17552 25504 17604
rect 25556 17552 25562 17604
rect 25590 17552 25596 17604
rect 25648 17592 25654 17604
rect 25685 17595 25743 17601
rect 25685 17592 25697 17595
rect 25648 17564 25697 17592
rect 25648 17552 25654 17564
rect 25685 17561 25697 17564
rect 25731 17592 25743 17595
rect 25866 17592 25872 17604
rect 25731 17564 25872 17592
rect 25731 17561 25743 17564
rect 25685 17555 25743 17561
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 25958 17552 25964 17604
rect 26016 17552 26022 17604
rect 26329 17595 26387 17601
rect 26329 17561 26341 17595
rect 26375 17592 26387 17595
rect 26605 17595 26663 17601
rect 26605 17592 26617 17595
rect 26375 17564 26617 17592
rect 26375 17561 26387 17564
rect 26329 17555 26387 17561
rect 26605 17561 26617 17564
rect 26651 17592 26663 17595
rect 27448 17592 27476 17620
rect 26651 17564 27476 17592
rect 26651 17561 26663 17564
rect 26605 17555 26663 17561
rect 25976 17524 26004 17552
rect 25424 17496 26004 17524
rect 24443 17493 24455 17496
rect 24397 17487 24455 17493
rect 1104 17434 43884 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 43884 17434
rect 1104 17360 43884 17382
rect 1670 17280 1676 17332
rect 1728 17280 1734 17332
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 3292 17292 3617 17320
rect 3292 17280 3298 17292
rect 3605 17289 3617 17292
rect 3651 17289 3663 17323
rect 3605 17283 3663 17289
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 4856 17292 5089 17320
rect 4856 17280 4862 17292
rect 5077 17289 5089 17292
rect 5123 17289 5135 17323
rect 6086 17320 6092 17332
rect 5077 17283 5135 17289
rect 5368 17292 6092 17320
rect 3712 17224 5304 17252
rect 2032 17187 2090 17193
rect 2032 17153 2044 17187
rect 2078 17184 2090 17187
rect 3326 17184 3332 17196
rect 2078 17156 3332 17184
rect 2078 17153 2090 17156
rect 2032 17147 2090 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 3712 17193 3740 17224
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 3964 17187 4022 17193
rect 3964 17153 3976 17187
rect 4010 17184 4022 17187
rect 4890 17184 4896 17196
rect 4010 17156 4896 17184
rect 4010 17153 4022 17156
rect 3964 17147 4022 17153
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 1762 17076 1768 17128
rect 1820 17076 1826 17128
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 2924 17088 3249 17116
rect 2924 17076 2930 17088
rect 3237 17085 3249 17088
rect 3283 17116 3295 17119
rect 3804 17116 3832 17144
rect 3283 17088 3832 17116
rect 5276 17116 5304 17224
rect 5368 17193 5396 17292
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6362 17280 6368 17332
rect 6420 17280 6426 17332
rect 6822 17320 6828 17332
rect 6564 17292 6828 17320
rect 5442 17212 5448 17264
rect 5500 17212 5506 17264
rect 5534 17212 5540 17264
rect 5592 17212 5598 17264
rect 5626 17212 5632 17264
rect 5684 17261 5690 17264
rect 5684 17255 5713 17261
rect 5701 17252 5713 17255
rect 5905 17255 5963 17261
rect 5701 17224 5856 17252
rect 5701 17221 5713 17224
rect 5684 17215 5713 17221
rect 5684 17212 5690 17215
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5828 17184 5856 17224
rect 5905 17221 5917 17255
rect 5951 17252 5963 17255
rect 5994 17252 6000 17264
rect 5951 17224 6000 17252
rect 5951 17221 5963 17224
rect 5905 17215 5963 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 5828 17156 6040 17184
rect 5353 17147 5411 17153
rect 5626 17116 5632 17128
rect 5276 17088 5632 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5736 17088 5825 17116
rect 5736 17060 5764 17088
rect 5813 17085 5825 17088
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 5902 17076 5908 17128
rect 5960 17076 5966 17128
rect 6012 17116 6040 17156
rect 6086 17144 6092 17196
rect 6144 17144 6150 17196
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 6454 17184 6460 17196
rect 6227 17156 6460 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 6564 17193 6592 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 8478 17320 8484 17332
rect 8036 17292 8484 17320
rect 6641 17255 6699 17261
rect 6641 17221 6653 17255
rect 6687 17252 6699 17255
rect 7098 17252 7104 17264
rect 6687 17224 7104 17252
rect 6687 17221 6699 17224
rect 6641 17215 6699 17221
rect 7098 17212 7104 17224
rect 7156 17212 7162 17264
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6730 17144 6736 17196
rect 6788 17144 6794 17196
rect 6851 17187 6909 17193
rect 6851 17153 6863 17187
rect 6897 17153 6909 17187
rect 6851 17147 6909 17153
rect 6866 17116 6894 17147
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 6012 17088 6894 17116
rect 5442 17048 5448 17060
rect 4632 17020 5448 17048
rect 3145 16983 3203 16989
rect 3145 16949 3157 16983
rect 3191 16980 3203 16983
rect 3234 16980 3240 16992
rect 3191 16952 3240 16980
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 3234 16940 3240 16952
rect 3292 16980 3298 16992
rect 4062 16980 4068 16992
rect 3292 16952 4068 16980
rect 3292 16940 3298 16952
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4430 16940 4436 16992
rect 4488 16980 4494 16992
rect 4632 16980 4660 17020
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 5718 17008 5724 17060
rect 5776 17008 5782 17060
rect 4488 16952 4660 16980
rect 4488 16940 4494 16952
rect 5166 16940 5172 16992
rect 5224 16940 5230 16992
rect 5920 16989 5948 17076
rect 6866 17048 6894 17088
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7558 17116 7564 17128
rect 7055 17088 7564 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7558 17076 7564 17088
rect 7616 17116 7622 17128
rect 7760 17116 7788 17280
rect 7926 17212 7932 17264
rect 7984 17212 7990 17264
rect 7616 17088 7788 17116
rect 7944 17116 7972 17212
rect 8036 17193 8064 17292
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10502 17320 10508 17332
rect 9600 17292 10508 17320
rect 8110 17212 8116 17264
rect 8168 17212 8174 17264
rect 9600 17252 9628 17292
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 11330 17280 11336 17332
rect 11388 17280 11394 17332
rect 11698 17320 11704 17332
rect 11440 17292 11704 17320
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 8496 17224 9628 17252
rect 9692 17224 9965 17252
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 8021 17147 8079 17153
rect 8128 17156 8217 17184
rect 8128 17116 8156 17156
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8323 17187 8381 17193
rect 8323 17184 8335 17187
rect 8205 17147 8263 17153
rect 8312 17153 8335 17184
rect 8369 17184 8381 17187
rect 8496 17184 8524 17224
rect 9692 17196 9720 17224
rect 9953 17221 9965 17224
rect 9999 17252 10011 17255
rect 10226 17252 10232 17264
rect 9999 17224 10232 17252
rect 9999 17221 10011 17224
rect 9953 17215 10011 17221
rect 10226 17212 10232 17224
rect 10284 17252 10290 17264
rect 11348 17252 11376 17280
rect 10284 17224 11008 17252
rect 10284 17212 10290 17224
rect 8369 17156 8524 17184
rect 8369 17153 8381 17156
rect 8312 17147 8381 17153
rect 8312 17116 8340 17147
rect 8662 17144 8668 17196
rect 8720 17144 8726 17196
rect 9398 17144 9404 17196
rect 9456 17144 9462 17196
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 9824 17156 10057 17184
rect 9824 17144 9830 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10778 17184 10784 17196
rect 10045 17147 10103 17153
rect 10152 17156 10784 17184
rect 7944 17088 8156 17116
rect 8220 17088 8340 17116
rect 7616 17076 7622 17088
rect 8220 17048 8248 17088
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8536 17088 9229 17116
rect 8536 17076 8542 17088
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 10152 17116 10180 17156
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 10980 17193 11008 17224
rect 11072 17224 11376 17252
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 9217 17079 9275 17085
rect 9646 17088 10180 17116
rect 6866 17020 8248 17048
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 9646 17048 9674 17088
rect 11072 17048 11100 17224
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11440 17184 11468 17292
rect 11698 17280 11704 17292
rect 11756 17320 11762 17332
rect 12066 17320 12072 17332
rect 11756 17292 12072 17320
rect 11756 17280 11762 17292
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12342 17280 12348 17332
rect 12400 17280 12406 17332
rect 12710 17280 12716 17332
rect 12768 17280 12774 17332
rect 12894 17280 12900 17332
rect 12952 17280 12958 17332
rect 13078 17280 13084 17332
rect 13136 17280 13142 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17289 13231 17323
rect 13173 17283 13231 17289
rect 11784 17255 11842 17261
rect 11784 17221 11796 17255
rect 11830 17252 11842 17255
rect 12360 17252 12388 17280
rect 11830 17224 12388 17252
rect 12728 17252 12756 17280
rect 13188 17252 13216 17283
rect 13446 17280 13452 17332
rect 13504 17280 13510 17332
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 14918 17280 14924 17332
rect 14976 17320 14982 17332
rect 17494 17320 17500 17332
rect 14976 17292 17500 17320
rect 14976 17280 14982 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 20272 17292 20484 17320
rect 13262 17252 13268 17264
rect 12728 17224 13268 17252
rect 11830 17221 11842 17224
rect 11784 17215 11842 17221
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 14568 17252 14596 17280
rect 14568 17224 15516 17252
rect 11379 17156 11468 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12584 17156 13001 17184
rect 12584 17144 12590 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 13228 17156 13369 17184
rect 13228 17144 13234 17156
rect 13357 17153 13369 17156
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 13909 17187 13967 17193
rect 13679 17156 13860 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 11514 17076 11520 17128
rect 11572 17076 11578 17128
rect 8352 17020 9674 17048
rect 9784 17020 11100 17048
rect 13832 17048 13860 17156
rect 13909 17153 13921 17187
rect 13955 17184 13967 17187
rect 13998 17184 14004 17196
rect 13955 17156 14004 17184
rect 13955 17153 13967 17156
rect 13909 17147 13967 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17184 14243 17187
rect 14366 17184 14372 17196
rect 14231 17156 14372 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 15304 17116 15332 17144
rect 14967 17088 15332 17116
rect 15488 17116 15516 17224
rect 15672 17224 15884 17252
rect 15672 17206 15700 17224
rect 15586 17193 15700 17206
rect 15565 17187 15700 17193
rect 15565 17153 15577 17187
rect 15611 17178 15700 17187
rect 15749 17187 15807 17193
rect 15611 17153 15623 17178
rect 15565 17147 15623 17153
rect 15749 17153 15761 17187
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15764 17116 15792 17147
rect 15488 17088 15792 17116
rect 15856 17116 15884 17224
rect 15930 17212 15936 17264
rect 15988 17212 15994 17264
rect 16298 17212 16304 17264
rect 16356 17212 16362 17264
rect 18892 17252 18920 17280
rect 19705 17255 19763 17261
rect 17052 17224 18552 17252
rect 18892 17224 19656 17252
rect 15948 17184 15976 17212
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15948 17156 16037 17184
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16316 17116 16344 17212
rect 17052 17193 17080 17224
rect 18524 17196 18552 17224
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 15856 17088 16344 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 13998 17048 14004 17060
rect 13832 17020 14004 17048
rect 8352 17008 8358 17020
rect 5905 16983 5963 16989
rect 5905 16949 5917 16983
rect 5951 16949 5963 16983
rect 5905 16943 5963 16949
rect 7006 16940 7012 16992
rect 7064 16980 7070 16992
rect 9784 16980 9812 17020
rect 13998 17008 14004 17020
rect 14056 17048 14062 17060
rect 15010 17048 15016 17060
rect 14056 17020 15016 17048
rect 14056 17008 14062 17020
rect 15010 17008 15016 17020
rect 15068 17048 15074 17060
rect 16209 17051 16267 17057
rect 16209 17048 16221 17051
rect 15068 17020 16221 17048
rect 15068 17008 15074 17020
rect 16209 17017 16221 17020
rect 16255 17017 16267 17051
rect 16209 17011 16267 17017
rect 16298 17008 16304 17060
rect 16356 17008 16362 17060
rect 17144 17048 17172 17147
rect 17218 17076 17224 17128
rect 17276 17076 17282 17128
rect 17512 17116 17540 17147
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17736 17156 17785 17184
rect 17736 17144 17742 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18322 17184 18328 17196
rect 17911 17156 18328 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 17880 17116 17908 17147
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 17512 17088 17908 17116
rect 18432 17116 18460 17147
rect 18506 17144 18512 17196
rect 18564 17184 18570 17196
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 18564 17156 19073 17184
rect 18564 17144 18570 17156
rect 19061 17153 19073 17156
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 18598 17116 18604 17128
rect 18432 17088 18604 17116
rect 18432 17048 18460 17088
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19076 17116 19104 17147
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 19628 17193 19656 17224
rect 19705 17221 19717 17255
rect 19751 17252 19763 17255
rect 20272 17252 20300 17292
rect 19751 17224 20300 17252
rect 20456 17252 20484 17292
rect 20622 17280 20628 17332
rect 20680 17280 20686 17332
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 20956 17292 21281 17320
rect 20956 17280 20962 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 21269 17283 21327 17289
rect 21637 17323 21695 17329
rect 21637 17289 21649 17323
rect 21683 17289 21695 17323
rect 21637 17283 21695 17289
rect 21082 17252 21088 17264
rect 20456 17224 21088 17252
rect 19751 17221 19763 17224
rect 19705 17215 19763 17221
rect 21082 17212 21088 17224
rect 21140 17212 21146 17264
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 19208 17156 19257 17184
rect 19208 17144 19214 17156
rect 19245 17153 19257 17156
rect 19291 17184 19303 17187
rect 19613 17187 19671 17193
rect 19291 17156 19564 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19536 17116 19564 17156
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19794 17144 19800 17196
rect 19852 17144 19858 17196
rect 19886 17144 19892 17196
rect 19944 17184 19950 17196
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19944 17156 19993 17184
rect 19944 17144 19950 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20070 17144 20076 17196
rect 20128 17144 20134 17196
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17184 20499 17187
rect 20993 17187 21051 17193
rect 20993 17184 21005 17187
rect 20487 17156 21005 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 20993 17153 21005 17156
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 20456 17116 20484 17147
rect 19076 17088 19288 17116
rect 19536 17088 20484 17116
rect 19260 17060 19288 17088
rect 17144 17020 18460 17048
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 21008 17048 21036 17147
rect 21284 17048 21312 17283
rect 21358 17212 21364 17264
rect 21416 17212 21422 17264
rect 21652 17184 21680 17283
rect 22462 17280 22468 17332
rect 22520 17280 22526 17332
rect 22830 17280 22836 17332
rect 22888 17280 22894 17332
rect 22922 17280 22928 17332
rect 22980 17280 22986 17332
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 24489 17323 24547 17329
rect 24489 17320 24501 17323
rect 23348 17292 24501 17320
rect 23348 17280 23354 17292
rect 24489 17289 24501 17292
rect 24535 17320 24547 17323
rect 24762 17320 24768 17332
rect 24535 17292 24768 17320
rect 24535 17289 24547 17292
rect 24489 17283 24547 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 43254 17280 43260 17332
rect 43312 17280 43318 17332
rect 22005 17255 22063 17261
rect 22005 17221 22017 17255
rect 22051 17252 22063 17255
rect 22646 17252 22652 17264
rect 22051 17224 22652 17252
rect 22051 17221 22063 17224
rect 22005 17215 22063 17221
rect 22646 17212 22652 17224
rect 22704 17212 22710 17264
rect 22940 17252 22968 17280
rect 22940 17224 23428 17252
rect 21726 17184 21732 17196
rect 21652 17156 21732 17184
rect 21726 17144 21732 17156
rect 21784 17144 21790 17196
rect 22741 17187 22799 17193
rect 22020 17156 22692 17184
rect 21450 17076 21456 17128
rect 21508 17125 21514 17128
rect 21508 17119 21536 17125
rect 21524 17085 21536 17119
rect 21508 17079 21536 17085
rect 21508 17076 21514 17079
rect 22020 17060 22048 17156
rect 22557 17119 22615 17125
rect 22557 17085 22569 17119
rect 22603 17085 22615 17119
rect 22664 17116 22692 17156
rect 22741 17153 22753 17187
rect 22787 17184 22799 17187
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22787 17156 23029 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23106 17144 23112 17196
rect 23164 17144 23170 17196
rect 23400 17193 23428 17224
rect 23474 17212 23480 17264
rect 23532 17252 23538 17264
rect 24029 17255 24087 17261
rect 24029 17252 24041 17255
rect 23532 17224 24041 17252
rect 23532 17212 23538 17224
rect 24029 17221 24041 17224
rect 24075 17252 24087 17255
rect 24302 17252 24308 17264
rect 24075 17224 24308 17252
rect 24075 17221 24087 17224
rect 24029 17215 24087 17221
rect 24302 17212 24308 17224
rect 24360 17212 24366 17264
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23566 17144 23572 17196
rect 23624 17144 23630 17196
rect 43162 17144 43168 17196
rect 43220 17144 43226 17196
rect 23845 17119 23903 17125
rect 23845 17116 23857 17119
rect 22664 17088 23857 17116
rect 22557 17079 22615 17085
rect 23845 17085 23857 17088
rect 23891 17085 23903 17119
rect 24670 17116 24676 17128
rect 23845 17079 23903 17085
rect 24320 17088 24676 17116
rect 22002 17048 22008 17060
rect 19300 17020 20484 17048
rect 21008 17020 21220 17048
rect 21284 17020 22008 17048
rect 19300 17008 19306 17020
rect 7064 16952 9812 16980
rect 7064 16940 7070 16952
rect 10686 16940 10692 16992
rect 10744 16940 10750 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 11848 16952 13093 16980
rect 11848 16940 11854 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13814 16940 13820 16992
rect 13872 16940 13878 16992
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14700 16952 14749 16980
rect 14700 16940 14706 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14737 16943 14795 16949
rect 15470 16940 15476 16992
rect 15528 16940 15534 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 16316 16980 16344 17008
rect 15703 16952 16344 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 19150 16980 19156 16992
rect 17736 16952 19156 16980
rect 17736 16940 17742 16952
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19429 16983 19487 16989
rect 19429 16949 19441 16983
rect 19475 16980 19487 16983
rect 19978 16980 19984 16992
rect 19475 16952 19984 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 19978 16940 19984 16952
rect 20036 16980 20042 16992
rect 20254 16980 20260 16992
rect 20036 16952 20260 16980
rect 20036 16940 20042 16952
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 20456 16989 20484 17020
rect 20441 16983 20499 16989
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 21082 16980 21088 16992
rect 20487 16952 21088 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21192 16980 21220 17020
rect 22002 17008 22008 17020
rect 22060 17008 22066 17060
rect 21910 16980 21916 16992
rect 21192 16952 21916 16980
rect 21910 16940 21916 16952
rect 21968 16980 21974 16992
rect 22572 16980 22600 17079
rect 23106 17008 23112 17060
rect 23164 17048 23170 17060
rect 24320 17048 24348 17088
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 23164 17020 24348 17048
rect 24397 17051 24455 17057
rect 23164 17008 23170 17020
rect 24397 17017 24409 17051
rect 24443 17048 24455 17051
rect 24486 17048 24492 17060
rect 24443 17020 24492 17048
rect 24443 17017 24455 17020
rect 24397 17011 24455 17017
rect 24486 17008 24492 17020
rect 24544 17008 24550 17060
rect 21968 16952 22600 16980
rect 21968 16940 21974 16952
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 1104 16890 43884 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 43884 16890
rect 1104 16816 43884 16838
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 3384 16748 4169 16776
rect 3384 16736 3390 16748
rect 4157 16745 4169 16748
rect 4203 16745 4215 16779
rect 4157 16739 4215 16745
rect 4890 16736 4896 16788
rect 4948 16736 4954 16788
rect 5166 16736 5172 16788
rect 5224 16736 5230 16788
rect 5626 16736 5632 16788
rect 5684 16776 5690 16788
rect 5684 16748 7420 16776
rect 5684 16736 5690 16748
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 2915 16680 4016 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16640 3571 16643
rect 3602 16640 3608 16652
rect 3559 16612 3608 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 3786 16600 3792 16652
rect 3844 16600 3850 16652
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 1627 16544 3004 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 1210 16464 1216 16516
rect 1268 16504 1274 16516
rect 2317 16507 2375 16513
rect 2317 16504 2329 16507
rect 1268 16476 2329 16504
rect 1268 16464 1274 16476
rect 2317 16473 2329 16476
rect 2363 16473 2375 16507
rect 2976 16504 3004 16544
rect 3050 16532 3056 16584
rect 3108 16572 3114 16584
rect 3988 16581 4016 16680
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 5184 16640 5212 16736
rect 5920 16649 5948 16748
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 7248 16680 7297 16708
rect 7248 16668 7254 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 4387 16612 5212 16640
rect 5905 16643 5963 16649
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 5905 16609 5917 16643
rect 5951 16609 5963 16643
rect 5905 16603 5963 16609
rect 7006 16600 7012 16652
rect 7064 16600 7070 16652
rect 3237 16575 3295 16581
rect 3237 16572 3249 16575
rect 3108 16544 3249 16572
rect 3108 16532 3114 16544
rect 3237 16541 3249 16544
rect 3283 16541 3295 16575
rect 3237 16535 3295 16541
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16541 3387 16575
rect 3329 16535 3387 16541
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 3344 16504 3372 16535
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 6172 16575 6230 16581
rect 6172 16541 6184 16575
rect 6218 16572 6230 16575
rect 6546 16572 6552 16584
rect 6218 16544 6552 16572
rect 6218 16541 6230 16544
rect 6172 16535 6230 16541
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 7024 16504 7052 16600
rect 7392 16581 7420 16748
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8720 16748 8769 16776
rect 8720 16736 8726 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 11514 16776 11520 16788
rect 9324 16748 11520 16776
rect 9324 16649 9352 16748
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 12250 16736 12256 16788
rect 12308 16736 12314 16788
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13814 16776 13820 16788
rect 13127 16748 13820 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 14185 16779 14243 16785
rect 14185 16745 14197 16779
rect 14231 16776 14243 16779
rect 14274 16776 14280 16788
rect 14231 16748 14280 16776
rect 14231 16745 14243 16748
rect 14185 16739 14243 16745
rect 14274 16736 14280 16748
rect 14332 16776 14338 16788
rect 15010 16776 15016 16788
rect 14332 16748 15016 16776
rect 14332 16736 14338 16748
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15712 16748 16313 16776
rect 15712 16736 15718 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 16758 16736 16764 16788
rect 16816 16736 16822 16788
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 17092 16748 17417 16776
rect 17092 16736 17098 16748
rect 17405 16745 17417 16748
rect 17451 16745 17463 16779
rect 17405 16739 17463 16745
rect 17494 16736 17500 16788
rect 17552 16736 17558 16788
rect 17586 16736 17592 16788
rect 17644 16736 17650 16788
rect 18509 16779 18567 16785
rect 18509 16745 18521 16779
rect 18555 16776 18567 16779
rect 18598 16776 18604 16788
rect 18555 16748 18604 16776
rect 18555 16745 18567 16748
rect 18509 16739 18567 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 18874 16736 18880 16788
rect 18932 16736 18938 16788
rect 19613 16779 19671 16785
rect 19613 16745 19625 16779
rect 19659 16776 19671 16779
rect 19886 16776 19892 16788
rect 19659 16748 19892 16776
rect 19659 16745 19671 16748
rect 19613 16739 19671 16745
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 10778 16708 10784 16720
rect 10376 16680 10784 16708
rect 10376 16668 10382 16680
rect 10778 16668 10784 16680
rect 10836 16708 10842 16720
rect 10965 16711 11023 16717
rect 10965 16708 10977 16711
rect 10836 16680 10977 16708
rect 10836 16668 10842 16680
rect 10965 16677 10977 16680
rect 11011 16677 11023 16711
rect 12268 16708 12296 16736
rect 13354 16708 13360 16720
rect 10965 16671 11023 16677
rect 11532 16680 13360 16708
rect 9309 16643 9367 16649
rect 8496 16612 9168 16640
rect 8496 16584 8524 16612
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 7466 16572 7472 16584
rect 7423 16544 7472 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7644 16575 7702 16581
rect 7644 16541 7656 16575
rect 7690 16572 7702 16575
rect 8386 16572 8392 16584
rect 7690 16544 8392 16572
rect 7690 16541 7702 16544
rect 7644 16535 7702 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 9140 16581 9168 16612
rect 9309 16609 9321 16643
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 2976 16476 7052 16504
rect 2317 16467 2375 16473
rect 8294 16464 8300 16516
rect 8352 16504 8358 16516
rect 8956 16504 8984 16535
rect 9398 16532 9404 16584
rect 9456 16532 9462 16584
rect 9576 16575 9634 16581
rect 9576 16541 9588 16575
rect 9622 16572 9634 16575
rect 10686 16572 10692 16584
rect 9622 16544 10692 16572
rect 9622 16541 9634 16544
rect 9576 16535 9634 16541
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11422 16572 11428 16584
rect 11379 16544 11428 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 11532 16581 11560 16680
rect 11974 16640 11980 16652
rect 11624 16612 11980 16640
rect 11624 16584 11652 16612
rect 11974 16600 11980 16612
rect 12032 16640 12038 16652
rect 12345 16643 12403 16649
rect 12032 16612 12204 16640
rect 12032 16600 12038 16612
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11606 16532 11612 16584
rect 11664 16532 11670 16584
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 12066 16572 12072 16584
rect 11931 16544 12072 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12176 16581 12204 16612
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12802 16640 12808 16652
rect 12391 16612 12808 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13280 16649 13308 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13556 16680 14320 16708
rect 13265 16643 13323 16649
rect 12912 16612 13216 16640
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 8352 16476 8984 16504
rect 8352 16464 8358 16476
rect 5626 16396 5632 16448
rect 5684 16396 5690 16448
rect 9416 16436 9444 16532
rect 12912 16504 12940 16612
rect 13188 16572 13216 16612
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13556 16572 13584 16680
rect 13906 16640 13912 16652
rect 13648 16612 13912 16640
rect 13648 16581 13676 16612
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 13998 16600 14004 16652
rect 14056 16600 14062 16652
rect 13008 16553 13066 16559
rect 13008 16550 13020 16553
rect 12084 16476 12940 16504
rect 13004 16519 13020 16550
rect 13054 16519 13066 16553
rect 13188 16544 13584 16572
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 13817 16575 13875 16581
rect 13817 16541 13829 16575
rect 13863 16572 13875 16575
rect 14016 16572 14044 16600
rect 14292 16581 14320 16680
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 15749 16711 15807 16717
rect 15436 16680 15516 16708
rect 15436 16668 15442 16680
rect 15488 16640 15516 16680
rect 15749 16677 15761 16711
rect 15795 16708 15807 16711
rect 15930 16708 15936 16720
rect 15795 16680 15936 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 16776 16708 16804 16736
rect 17129 16711 17187 16717
rect 17129 16708 17141 16711
rect 16776 16680 17141 16708
rect 17129 16677 17141 16680
rect 17175 16677 17187 16711
rect 17129 16671 17187 16677
rect 17310 16668 17316 16720
rect 17368 16668 17374 16720
rect 16298 16640 16304 16652
rect 15488 16612 16304 16640
rect 16298 16600 16304 16612
rect 16356 16640 16362 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16356 16612 16681 16640
rect 16356 16600 16362 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 13863 16544 14044 16572
rect 14093 16575 14151 16581
rect 13863 16541 13875 16544
rect 13817 16535 13875 16541
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 14458 16572 14464 16584
rect 14415 16544 14464 16572
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 13004 16513 13066 16519
rect 10689 16439 10747 16445
rect 10689 16436 10701 16439
rect 9416 16408 10701 16436
rect 10689 16405 10701 16408
rect 10735 16405 10747 16439
rect 10689 16399 10747 16405
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 11112 16408 11161 16436
rect 11112 16396 11118 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11974 16436 11980 16448
rect 11747 16408 11980 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12084 16445 12112 16476
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16405 12127 16439
rect 12069 16399 12127 16405
rect 12894 16396 12900 16448
rect 12952 16396 12958 16448
rect 13004 16436 13032 16513
rect 13262 16464 13268 16516
rect 13320 16464 13326 16516
rect 13354 16464 13360 16516
rect 13412 16504 13418 16516
rect 13449 16507 13507 16513
rect 13449 16504 13461 16507
rect 13412 16476 13461 16504
rect 13412 16464 13418 16476
rect 13449 16473 13461 16476
rect 13495 16473 13507 16507
rect 13449 16467 13507 16473
rect 13909 16507 13967 16513
rect 13909 16473 13921 16507
rect 13955 16504 13967 16507
rect 13998 16504 14004 16516
rect 13955 16476 14004 16504
rect 13955 16473 13967 16476
rect 13909 16467 13967 16473
rect 13998 16464 14004 16476
rect 14056 16464 14062 16516
rect 13630 16436 13636 16448
rect 13004 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16436 13694 16448
rect 14108 16436 14136 16535
rect 13688 16408 14136 16436
rect 14292 16436 14320 16535
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 14642 16581 14648 16584
rect 14636 16572 14648 16581
rect 14603 16544 14648 16572
rect 14636 16535 14648 16544
rect 14642 16532 14648 16535
rect 14700 16532 14706 16584
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15838 16572 15844 16584
rect 15436 16544 15844 16572
rect 15436 16532 15442 16544
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 17328 16581 17356 16668
rect 17604 16649 17632 16736
rect 18616 16708 18644 16736
rect 19628 16708 19656 16739
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 19981 16779 20039 16785
rect 19981 16745 19993 16779
rect 20027 16776 20039 16779
rect 25498 16776 25504 16788
rect 20027 16748 25504 16776
rect 20027 16745 20039 16748
rect 19981 16739 20039 16745
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 18616 16680 19656 16708
rect 19794 16668 19800 16720
rect 19852 16708 19858 16720
rect 19852 16680 20208 16708
rect 19852 16668 19858 16680
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 18601 16643 18659 16649
rect 18601 16640 18613 16643
rect 18380 16612 18613 16640
rect 18380 16600 18386 16612
rect 18601 16609 18613 16612
rect 18647 16640 18659 16643
rect 19058 16640 19064 16652
rect 18647 16612 19064 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 19058 16600 19064 16612
rect 19116 16640 19122 16652
rect 20180 16640 20208 16680
rect 20438 16668 20444 16720
rect 20496 16668 20502 16720
rect 24394 16708 24400 16720
rect 20548 16680 24400 16708
rect 20456 16640 20484 16668
rect 20548 16649 20576 16680
rect 24394 16668 24400 16680
rect 24452 16668 24458 16720
rect 19116 16612 19840 16640
rect 19116 16600 19122 16612
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16541 17371 16575
rect 17313 16535 17371 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 19150 16572 19156 16584
rect 18187 16544 19156 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18064 16504 18092 16535
rect 19150 16532 19156 16544
rect 19208 16572 19214 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 19208 16544 19257 16572
rect 19208 16532 19214 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16572 19671 16575
rect 19812 16572 19840 16612
rect 19904 16612 20116 16640
rect 19904 16581 19932 16612
rect 19659 16544 19840 16572
rect 19889 16575 19947 16581
rect 19659 16541 19671 16544
rect 19613 16535 19671 16541
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 19996 16504 20024 16535
rect 18064 16476 19288 16504
rect 19260 16448 19288 16476
rect 19444 16476 20024 16504
rect 20088 16504 20116 16612
rect 20180 16612 20484 16640
rect 20533 16643 20591 16649
rect 20180 16581 20208 16612
rect 20533 16609 20545 16643
rect 20579 16609 20591 16643
rect 20806 16640 20812 16652
rect 20533 16603 20591 16609
rect 20732 16612 20812 16640
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20441 16575 20499 16581
rect 20441 16572 20453 16575
rect 20312 16544 20453 16572
rect 20312 16532 20318 16544
rect 20441 16541 20453 16544
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 20622 16532 20628 16584
rect 20680 16532 20686 16584
rect 20732 16581 20760 16612
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 21542 16600 21548 16652
rect 21600 16600 21606 16652
rect 21913 16643 21971 16649
rect 21913 16609 21925 16643
rect 21959 16640 21971 16643
rect 22370 16640 22376 16652
rect 21959 16612 22376 16640
rect 21959 16609 21971 16612
rect 21913 16603 21971 16609
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 21082 16532 21088 16584
rect 21140 16572 21146 16584
rect 21450 16572 21456 16584
rect 21140 16544 21456 16572
rect 21140 16532 21146 16544
rect 21450 16532 21456 16544
rect 21508 16572 21514 16584
rect 21928 16572 21956 16603
rect 22370 16600 22376 16612
rect 22428 16640 22434 16652
rect 22649 16643 22707 16649
rect 22649 16640 22661 16643
rect 22428 16612 22661 16640
rect 22428 16600 22434 16612
rect 22649 16609 22661 16612
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 21508 16544 21956 16572
rect 21508 16532 21514 16544
rect 22094 16532 22100 16584
rect 22152 16532 22158 16584
rect 22462 16532 22468 16584
rect 22520 16532 22526 16584
rect 22554 16532 22560 16584
rect 22612 16572 22618 16584
rect 23014 16572 23020 16584
rect 22612 16544 23020 16572
rect 22612 16532 22618 16544
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 21100 16504 21128 16532
rect 20088 16476 21128 16504
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 14292 16408 16037 16436
rect 13688 16396 13694 16408
rect 16025 16405 16037 16408
rect 16071 16436 16083 16439
rect 16482 16436 16488 16448
rect 16071 16408 16488 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 19242 16396 19248 16448
rect 19300 16396 19306 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19444 16445 19472 16476
rect 21358 16464 21364 16516
rect 21416 16504 21422 16516
rect 21637 16507 21695 16513
rect 21637 16504 21649 16507
rect 21416 16476 21649 16504
rect 21416 16464 21422 16476
rect 21637 16473 21649 16476
rect 21683 16504 21695 16507
rect 22646 16504 22652 16516
rect 21683 16476 22652 16504
rect 21683 16473 21695 16476
rect 21637 16467 21695 16473
rect 22646 16464 22652 16476
rect 22704 16504 22710 16516
rect 23293 16507 23351 16513
rect 23293 16504 23305 16507
rect 22704 16476 23305 16504
rect 22704 16464 22710 16476
rect 23293 16473 23305 16476
rect 23339 16473 23351 16507
rect 23293 16467 23351 16473
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 19392 16408 19441 16436
rect 19392 16396 19398 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20809 16439 20867 16445
rect 20809 16436 20821 16439
rect 20772 16408 20821 16436
rect 20772 16396 20778 16408
rect 20809 16405 20821 16408
rect 20855 16405 20867 16439
rect 20809 16399 20867 16405
rect 21910 16396 21916 16448
rect 21968 16436 21974 16448
rect 22005 16439 22063 16445
rect 22005 16436 22017 16439
rect 21968 16408 22017 16436
rect 21968 16396 21974 16408
rect 22005 16405 22017 16408
rect 22051 16405 22063 16439
rect 22005 16399 22063 16405
rect 22278 16396 22284 16448
rect 22336 16396 22342 16448
rect 1104 16346 43884 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 43884 16346
rect 1104 16272 43884 16294
rect 2866 16232 2872 16244
rect 1688 16204 2872 16232
rect 1688 16108 1716 16204
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3421 16235 3479 16241
rect 3421 16201 3433 16235
rect 3467 16232 3479 16235
rect 4062 16232 4068 16244
rect 3467 16204 4068 16232
rect 3467 16201 3479 16204
rect 3421 16195 3479 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4617 16235 4675 16241
rect 4617 16201 4629 16235
rect 4663 16232 4675 16235
rect 4982 16232 4988 16244
rect 4663 16204 4988 16232
rect 4663 16201 4675 16204
rect 4617 16195 4675 16201
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 6052 16204 6101 16232
rect 6052 16192 6058 16204
rect 6089 16201 6101 16204
rect 6135 16201 6147 16235
rect 6089 16195 6147 16201
rect 7469 16235 7527 16241
rect 7469 16201 7481 16235
rect 7515 16232 7527 16235
rect 7558 16232 7564 16244
rect 7515 16204 7564 16232
rect 7515 16201 7527 16204
rect 7469 16195 7527 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8205 16235 8263 16241
rect 8205 16201 8217 16235
rect 8251 16232 8263 16235
rect 8478 16232 8484 16244
rect 8251 16204 8484 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 9732 16204 9781 16232
rect 9732 16192 9738 16204
rect 9769 16201 9781 16204
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 9858 16192 9864 16244
rect 9916 16192 9922 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 10100 16204 10149 16232
rect 10100 16192 10106 16204
rect 10137 16201 10149 16204
rect 10183 16201 10195 16235
rect 10137 16195 10195 16201
rect 10778 16192 10784 16244
rect 10836 16192 10842 16244
rect 11606 16192 11612 16244
rect 11664 16192 11670 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 12894 16232 12900 16244
rect 11931 16204 12900 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 15838 16192 15844 16244
rect 15896 16192 15902 16244
rect 16114 16192 16120 16244
rect 16172 16192 16178 16244
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 16816 16204 16865 16232
rect 16816 16192 16822 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 16853 16195 16911 16201
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 19521 16235 19579 16241
rect 19521 16232 19533 16235
rect 19484 16204 19533 16232
rect 19484 16192 19490 16204
rect 19521 16201 19533 16204
rect 19567 16201 19579 16235
rect 19521 16195 19579 16201
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 22462 16232 22468 16244
rect 20404 16204 22468 16232
rect 20404 16192 20410 16204
rect 22462 16192 22468 16204
rect 22520 16192 22526 16244
rect 23014 16192 23020 16244
rect 23072 16232 23078 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23072 16204 23213 16232
rect 23072 16192 23078 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 1949 16167 2007 16173
rect 1949 16133 1961 16167
rect 1995 16164 2007 16167
rect 2286 16167 2344 16173
rect 2286 16164 2298 16167
rect 1995 16136 2298 16164
rect 1995 16133 2007 16136
rect 1949 16127 2007 16133
rect 2286 16133 2298 16136
rect 2332 16133 2344 16167
rect 2286 16127 2344 16133
rect 3881 16167 3939 16173
rect 3881 16133 3893 16167
rect 3927 16164 3939 16167
rect 7009 16167 7067 16173
rect 7009 16164 7021 16167
rect 3927 16136 7021 16164
rect 3927 16133 3939 16136
rect 3881 16127 3939 16133
rect 7009 16133 7021 16136
rect 7055 16133 7067 16167
rect 9876 16164 9904 16192
rect 11624 16164 11652 16192
rect 7009 16127 7067 16133
rect 9600 16136 9904 16164
rect 10888 16136 11652 16164
rect 1670 16056 1676 16108
rect 1728 16056 1734 16108
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 1780 15892 1808 16059
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1912 16068 2053 16096
rect 1912 16056 1918 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 4890 16096 4896 16108
rect 2087 16068 3648 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2774 15892 2780 15904
rect 1780 15864 2780 15892
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 3510 15852 3516 15904
rect 3568 15852 3574 15904
rect 3620 15892 3648 16068
rect 3712 16068 4896 16096
rect 3712 16040 3740 16068
rect 3694 15988 3700 16040
rect 3752 15988 3758 16040
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4080 16037 4108 16068
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5031 16068 5488 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3936 16000 3985 16028
rect 3936 15988 3942 16000
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 15997 4123 16031
rect 4065 15991 4123 15997
rect 3988 15960 4016 15991
rect 4706 15988 4712 16040
rect 4764 16028 4770 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4764 16000 5089 16028
rect 4764 15988 4770 16000
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 5166 15988 5172 16040
rect 5224 15988 5230 16040
rect 5460 16028 5488 16068
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 6086 16096 6092 16108
rect 5592 16068 6092 16096
rect 5592 16056 5598 16068
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6454 16056 6460 16108
rect 6512 16056 6518 16108
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16096 7343 16099
rect 7374 16096 7380 16108
rect 7331 16068 7380 16096
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8202 16096 8208 16108
rect 8067 16068 8208 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 5994 16028 6000 16040
rect 5460 16000 6000 16028
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7576 16028 7604 16059
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9600 16105 9628 16136
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 9585 16099 9643 16105
rect 8343 16068 9536 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 8312 16028 8340 16059
rect 7524 16000 8340 16028
rect 7524 15988 7530 16000
rect 8754 15988 8760 16040
rect 8812 15988 8818 16040
rect 9508 16028 9536 16068
rect 9585 16065 9597 16099
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10888 16096 10916 16136
rect 11698 16124 11704 16176
rect 11756 16164 11762 16176
rect 12621 16167 12679 16173
rect 12621 16164 12633 16167
rect 11756 16136 12633 16164
rect 11756 16124 11762 16136
rect 12621 16133 12633 16136
rect 12667 16133 12679 16167
rect 12621 16127 12679 16133
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 14274 16164 14280 16176
rect 13872 16136 14280 16164
rect 13872 16124 13878 16136
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 14728 16167 14786 16173
rect 14728 16133 14740 16167
rect 14774 16164 14786 16167
rect 15470 16164 15476 16176
rect 14774 16136 15476 16164
rect 14774 16133 14786 16136
rect 14728 16127 14786 16133
rect 15470 16124 15476 16136
rect 15528 16124 15534 16176
rect 21358 16124 21364 16176
rect 21416 16164 21422 16176
rect 26878 16164 26884 16176
rect 21416 16136 26884 16164
rect 21416 16124 21422 16136
rect 9907 16068 10916 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 9876 16028 9904 16059
rect 10962 16056 10968 16108
rect 11020 16056 11026 16108
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 12308 16068 13645 16096
rect 12308 16056 12314 16068
rect 13633 16065 13645 16068
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14516 16068 17172 16096
rect 14516 16056 14522 16068
rect 9508 16000 9904 16028
rect 10980 15960 11008 16056
rect 17144 16040 17172 16068
rect 17402 16056 17408 16108
rect 17460 16056 17466 16108
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 19058 16096 19064 16108
rect 19015 16068 19064 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19208 16068 19257 16096
rect 19208 16056 19214 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 20524 16099 20582 16105
rect 20524 16065 20536 16099
rect 20570 16096 20582 16099
rect 20570 16068 21772 16096
rect 20570 16065 20582 16068
rect 20524 16059 20582 16065
rect 11974 15988 11980 16040
rect 12032 15988 12038 16040
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 3988 15932 11008 15960
rect 11241 15963 11299 15969
rect 11241 15929 11253 15963
rect 11287 15960 11299 15963
rect 12084 15960 12112 15991
rect 12986 15988 12992 16040
rect 13044 15988 13050 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17267 16000 18000 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 11287 15932 12112 15960
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 4062 15892 4068 15904
rect 3620 15864 4068 15892
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 7098 15852 7104 15904
rect 7156 15852 7162 15904
rect 7742 15852 7748 15904
rect 7800 15892 7806 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 7800 15864 7849 15892
rect 7800 15852 7806 15864
rect 7837 15861 7849 15864
rect 7883 15861 7895 15895
rect 7837 15855 7895 15861
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 9309 15895 9367 15901
rect 9309 15892 9321 15895
rect 8536 15864 9321 15892
rect 8536 15852 8542 15864
rect 9309 15861 9321 15864
rect 9355 15861 9367 15895
rect 9309 15855 9367 15861
rect 9398 15852 9404 15904
rect 9456 15852 9462 15904
rect 11330 15852 11336 15904
rect 11388 15892 11394 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11388 15864 11529 15892
rect 11388 15852 11394 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 12084 15892 12112 15932
rect 17972 15904 18000 16000
rect 20254 15988 20260 16040
rect 20312 15988 20318 16040
rect 21634 15920 21640 15972
rect 21692 15920 21698 15972
rect 13170 15892 13176 15904
rect 12084 15864 13176 15892
rect 11517 15855 11575 15861
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 17460 15864 17601 15892
rect 17460 15852 17466 15864
rect 17589 15861 17601 15864
rect 17635 15861 17647 15895
rect 17589 15855 17647 15861
rect 17954 15852 17960 15904
rect 18012 15852 18018 15904
rect 19242 15852 19248 15904
rect 19300 15852 19306 15904
rect 21744 15892 21772 16068
rect 21836 16037 21864 16136
rect 26878 16124 26884 16136
rect 26936 16124 26942 16176
rect 28350 16124 28356 16176
rect 28408 16124 28414 16176
rect 22088 16099 22146 16105
rect 22088 16065 22100 16099
rect 22134 16096 22146 16099
rect 28368 16096 28396 16124
rect 22134 16068 28396 16096
rect 22134 16065 22146 16068
rect 22088 16059 22146 16065
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 28810 15892 28816 15904
rect 21744 15864 28816 15892
rect 28810 15852 28816 15864
rect 28868 15852 28874 15904
rect 1104 15802 43884 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 43884 15802
rect 1104 15728 43884 15750
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 3605 15691 3663 15697
rect 3605 15688 3617 15691
rect 3476 15660 3617 15688
rect 3476 15648 3482 15660
rect 3605 15657 3617 15660
rect 3651 15657 3663 15691
rect 3605 15651 3663 15657
rect 3878 15648 3884 15700
rect 3936 15648 3942 15700
rect 5626 15688 5632 15700
rect 3988 15660 5632 15688
rect 1210 15512 1216 15564
rect 1268 15552 1274 15564
rect 1857 15555 1915 15561
rect 1857 15552 1869 15555
rect 1268 15524 1869 15552
rect 1268 15512 1274 15524
rect 1857 15521 1869 15524
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 3053 15555 3111 15561
rect 3053 15521 3065 15555
rect 3099 15552 3111 15555
rect 3142 15552 3148 15564
rect 3099 15524 3148 15552
rect 3099 15521 3111 15524
rect 3053 15515 3111 15521
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 3896 15552 3924 15648
rect 3804 15524 3924 15552
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 3804 15484 3832 15524
rect 3988 15493 4016 15660
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7469 15691 7527 15697
rect 7469 15688 7481 15691
rect 7340 15660 7481 15688
rect 7340 15648 7346 15660
rect 7469 15657 7481 15660
rect 7515 15657 7527 15691
rect 7469 15651 7527 15657
rect 8018 15648 8024 15700
rect 8076 15688 8082 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8076 15660 8585 15688
rect 8076 15648 8082 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 8754 15648 8760 15700
rect 8812 15688 8818 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8812 15660 8953 15688
rect 8812 15648 8818 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 11330 15688 11336 15700
rect 8941 15651 8999 15657
rect 10796 15660 11336 15688
rect 5258 15580 5264 15632
rect 5316 15620 5322 15632
rect 5316 15592 9536 15620
rect 5316 15580 5322 15592
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 6288 15561 6316 15592
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8110 15552 8116 15564
rect 8067 15524 8116 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8110 15512 8116 15524
rect 8168 15552 8174 15564
rect 9214 15552 9220 15564
rect 8168 15524 9220 15552
rect 8168 15512 8174 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9508 15561 9536 15592
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15552 9551 15555
rect 9766 15552 9772 15564
rect 9539 15524 9772 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 9950 15552 9956 15564
rect 9907 15524 9956 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 1627 15456 3832 15484
rect 3881 15487 3939 15493
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 3881 15453 3893 15487
rect 3927 15453 3939 15487
rect 3881 15447 3939 15453
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 3786 15376 3792 15428
rect 3844 15416 3850 15428
rect 3896 15416 3924 15447
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4120 15456 4261 15484
rect 4120 15444 4126 15456
rect 4249 15453 4261 15456
rect 4295 15484 4307 15487
rect 5258 15484 5264 15496
rect 4295 15456 5264 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5408 15456 5856 15484
rect 5408 15444 5414 15456
rect 3844 15388 3924 15416
rect 4157 15419 4215 15425
rect 3844 15376 3850 15388
rect 4157 15385 4169 15419
rect 4203 15416 4215 15419
rect 4494 15419 4552 15425
rect 4494 15416 4506 15419
rect 4203 15388 4506 15416
rect 4203 15385 4215 15388
rect 4157 15379 4215 15385
rect 4494 15385 4506 15388
rect 4540 15385 4552 15419
rect 4494 15379 4552 15385
rect 4798 15376 4804 15428
rect 4856 15416 4862 15428
rect 4856 15388 5764 15416
rect 4856 15376 4862 15388
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 5736 15357 5764 15388
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5592 15320 5641 15348
rect 5592 15308 5598 15320
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 5629 15311 5687 15317
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15317 5779 15351
rect 5828 15348 5856 15456
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5960 15456 6101 15484
rect 5960 15444 5966 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6196 15484 6224 15512
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 6196 15456 6561 15484
rect 6089 15447 6147 15453
rect 6549 15453 6561 15456
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 6104 15416 6132 15447
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 10796 15493 10824 15660
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 12437 15691 12495 15697
rect 12437 15657 12449 15691
rect 12483 15688 12495 15691
rect 12802 15688 12808 15700
rect 12483 15660 12808 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13722 15648 13728 15700
rect 13780 15648 13786 15700
rect 17126 15648 17132 15700
rect 17184 15688 17190 15700
rect 20254 15688 20260 15700
rect 17184 15660 20260 15688
rect 17184 15648 17190 15660
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 22462 15648 22468 15700
rect 22520 15688 22526 15700
rect 22741 15691 22799 15697
rect 22741 15688 22753 15691
rect 22520 15660 22753 15688
rect 22520 15648 22526 15660
rect 22741 15657 22753 15660
rect 22787 15657 22799 15691
rect 22741 15651 22799 15657
rect 13740 15620 13768 15648
rect 15010 15620 15016 15632
rect 13740 15592 14504 15620
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13906 15552 13912 15564
rect 13403 15524 13912 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 10597 15487 10655 15493
rect 8996 15456 9352 15484
rect 8996 15444 9002 15456
rect 9324 15425 9352 15456
rect 10597 15453 10609 15487
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 10781 15487 10839 15493
rect 10781 15453 10793 15487
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15484 11115 15487
rect 11103 15456 11560 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 7193 15419 7251 15425
rect 7193 15416 7205 15419
rect 6104 15388 7205 15416
rect 7193 15385 7205 15388
rect 7239 15385 7251 15419
rect 7193 15379 7251 15385
rect 9309 15419 9367 15425
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 9355 15388 10425 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10413 15379 10471 15385
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 5828 15320 6193 15348
rect 5721 15311 5779 15317
rect 6181 15317 6193 15320
rect 6227 15317 6239 15351
rect 6181 15311 6239 15317
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 7374 15348 7380 15360
rect 6880 15320 7380 15348
rect 6880 15308 6886 15320
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 9398 15308 9404 15360
rect 9456 15308 9462 15360
rect 10612 15348 10640 15447
rect 11532 15428 11560 15456
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 14476 15493 14504 15592
rect 14660 15592 15016 15620
rect 14660 15561 14688 15592
rect 15010 15580 15016 15592
rect 15068 15620 15074 15632
rect 15562 15620 15568 15632
rect 15068 15592 15568 15620
rect 15068 15580 15074 15592
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 16022 15580 16028 15632
rect 16080 15580 16086 15632
rect 16298 15580 16304 15632
rect 16356 15580 16362 15632
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15521 14703 15555
rect 14645 15515 14703 15521
rect 14734 15512 14740 15564
rect 14792 15552 14798 15564
rect 17144 15561 17172 15648
rect 18506 15580 18512 15632
rect 18564 15580 18570 15632
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14792 15524 14933 15552
rect 14792 15512 14798 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 17402 15493 17408 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12308 15456 12909 15484
rect 12308 15444 12314 15456
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14461 15487 14519 15493
rect 13587 15456 14136 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 10965 15419 11023 15425
rect 10965 15385 10977 15419
rect 11011 15416 11023 15419
rect 11302 15419 11360 15425
rect 11302 15416 11314 15419
rect 11011 15388 11314 15416
rect 11011 15385 11023 15388
rect 10965 15379 11023 15385
rect 11302 15385 11314 15388
rect 11348 15385 11360 15419
rect 11302 15379 11360 15385
rect 11514 15376 11520 15428
rect 11572 15376 11578 15428
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 12406 15388 13001 15416
rect 10870 15348 10876 15360
rect 10612 15320 10876 15348
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 12406 15348 12434 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 12989 15379 13047 15385
rect 11112 15320 12434 15348
rect 11112 15308 11118 15320
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 14108 15357 14136 15456
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 14507 15456 15577 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 17396 15484 17408 15493
rect 17363 15456 17408 15484
rect 15565 15447 15623 15453
rect 17396 15447 17408 15456
rect 17402 15444 17408 15447
rect 17460 15444 17466 15496
rect 21628 15487 21686 15493
rect 21628 15453 21640 15487
rect 21674 15484 21686 15487
rect 26050 15484 26056 15496
rect 21674 15456 26056 15484
rect 21674 15453 21686 15456
rect 21628 15447 21686 15453
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 22738 15416 22744 15428
rect 18012 15388 22744 15416
rect 18012 15376 18018 15388
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13504 15320 13737 15348
rect 13504 15308 13510 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14550 15308 14556 15360
rect 14608 15308 14614 15360
rect 1104 15258 43884 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 43884 15258
rect 1104 15184 43884 15206
rect 1670 15104 1676 15156
rect 1728 15104 1734 15156
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2832 15116 2881 15144
rect 2832 15104 2838 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 3050 15104 3056 15156
rect 3108 15144 3114 15156
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 3108 15116 3617 15144
rect 3108 15104 3114 15116
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 3605 15107 3663 15113
rect 3970 15104 3976 15156
rect 4028 15104 4034 15156
rect 5445 15147 5503 15153
rect 5445 15113 5457 15147
rect 5491 15144 5503 15147
rect 6178 15144 6184 15156
rect 5491 15116 6184 15144
rect 5491 15113 5503 15116
rect 5445 15107 5503 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 7466 15144 7472 15156
rect 6564 15116 7472 15144
rect 2038 15036 2044 15088
rect 2096 15076 2102 15088
rect 2096 15048 5764 15076
rect 2096 15036 2102 15048
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3234 15008 3240 15020
rect 3099 14980 3240 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 4062 14968 4068 15020
rect 4120 14968 4126 15020
rect 4332 15011 4390 15017
rect 4332 14977 4344 15011
rect 4378 15008 4390 15011
rect 4614 15008 4620 15020
rect 4378 14980 4620 15008
rect 4378 14977 4390 14980
rect 4332 14971 4390 14977
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 5736 15017 5764 15048
rect 5810 15036 5816 15088
rect 5868 15076 5874 15088
rect 5905 15079 5963 15085
rect 5905 15076 5917 15079
rect 5868 15048 5917 15076
rect 5868 15036 5874 15048
rect 5905 15045 5917 15048
rect 5951 15045 5963 15079
rect 6564 15076 6592 15116
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 7558 15104 7564 15156
rect 7616 15104 7622 15156
rect 7653 15147 7711 15153
rect 7653 15113 7665 15147
rect 7699 15144 7711 15147
rect 8018 15144 8024 15156
rect 7699 15116 8024 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8481 15147 8539 15153
rect 8481 15113 8493 15147
rect 8527 15144 8539 15147
rect 8527 15116 8708 15144
rect 8527 15113 8539 15116
rect 8481 15107 8539 15113
rect 5905 15039 5963 15045
rect 6012 15048 6592 15076
rect 6012 15017 6040 15048
rect 6730 15036 6736 15088
rect 6788 15036 6794 15088
rect 7576 15076 7604 15104
rect 8680 15076 8708 15116
rect 9950 15104 9956 15156
rect 10008 15104 10014 15156
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10778 15144 10784 15156
rect 10459 15116 10784 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 12526 15144 12532 15156
rect 11440 15116 12532 15144
rect 8818 15079 8876 15085
rect 8818 15076 8830 15079
rect 7576 15048 8616 15076
rect 8680 15048 8830 15076
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 7009 15011 7067 15017
rect 7208 15014 7328 15030
rect 7009 14977 7021 15011
rect 7055 14998 7067 15011
rect 7122 15002 7328 15014
rect 7122 14998 7236 15002
rect 7055 14986 7236 14998
rect 7055 14977 7150 14986
rect 7009 14971 7150 14977
rect 7027 14970 7150 14971
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2363 14912 2774 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2746 14872 2774 14912
rect 3510 14900 3516 14952
rect 3568 14900 3574 14952
rect 5810 14900 5816 14952
rect 5868 14900 5874 14952
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 3528 14872 3556 14900
rect 2746 14844 3556 14872
rect 5828 14872 5856 14900
rect 6840 14872 6868 14900
rect 7300 14881 7328 15002
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7432 14980 8125 15008
rect 7432 14968 7438 14980
rect 8113 14977 8125 14980
rect 8159 15008 8171 15011
rect 8202 15008 8208 15020
rect 8159 14980 8208 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8478 15008 8484 15020
rect 8343 14980 8484 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8588 15017 8616 15048
rect 8818 15045 8830 15048
rect 8864 15045 8876 15079
rect 8818 15039 8876 15045
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11440 15008 11468 15116
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 12986 15144 12992 15156
rect 12943 15116 12992 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 14553 15147 14611 15153
rect 14553 15113 14565 15147
rect 14599 15144 14611 15147
rect 14734 15144 14740 15156
rect 14599 15116 14740 15144
rect 14599 15113 14611 15116
rect 14553 15107 14611 15113
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 15010 15104 15016 15156
rect 15068 15104 15074 15156
rect 11624 15048 14504 15076
rect 11195 14980 11468 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 11624 15008 11652 15048
rect 11790 15017 11796 15020
rect 11784 15008 11796 15017
rect 11572 14980 11652 15008
rect 11751 14980 11796 15008
rect 11572 14968 11578 14980
rect 11784 14971 11796 14980
rect 11790 14968 11796 14971
rect 11848 14968 11854 15020
rect 13188 15017 13216 15048
rect 14476 15020 14504 15048
rect 13446 15017 13452 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 14977 13231 15011
rect 13440 15008 13452 15017
rect 13407 14980 13452 15008
rect 13173 14971 13231 14977
rect 13440 14971 13452 14980
rect 13446 14968 13452 14971
rect 13504 14968 13510 15020
rect 14458 14968 14464 15020
rect 14516 14968 14522 15020
rect 7742 14900 7748 14952
rect 7800 14900 7806 14952
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 7929 14903 7987 14909
rect 10888 14912 10977 14940
rect 5828 14844 6868 14872
rect 7285 14875 7343 14881
rect 7285 14841 7297 14875
rect 7331 14841 7343 14875
rect 7285 14835 7343 14841
rect 2133 14807 2191 14813
rect 2133 14773 2145 14807
rect 2179 14804 2191 14807
rect 3234 14804 3240 14816
rect 2179 14776 3240 14804
rect 2179 14773 2191 14776
rect 2133 14767 2191 14773
rect 3234 14764 3240 14776
rect 3292 14804 3298 14816
rect 3694 14804 3700 14816
rect 3292 14776 3700 14804
rect 3292 14764 3298 14776
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5537 14807 5595 14813
rect 5537 14804 5549 14807
rect 4764 14776 5549 14804
rect 4764 14764 4770 14776
rect 5537 14773 5549 14776
rect 5583 14773 5595 14807
rect 5537 14767 5595 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 7944 14804 7972 14903
rect 10888 14816 10916 14912
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 7432 14776 7972 14804
rect 7432 14764 7438 14776
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11790 14804 11796 14816
rect 11379 14776 11796 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 1104 14714 43884 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 43884 14714
rect 1104 14640 43884 14662
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3292 14572 3525 14600
rect 3292 14560 3298 14572
rect 3513 14569 3525 14572
rect 3559 14569 3571 14603
rect 3513 14563 3571 14569
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4614 14600 4620 14612
rect 4203 14572 4620 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 6641 14603 6699 14609
rect 5276 14572 6597 14600
rect 4525 14535 4583 14541
rect 4525 14501 4537 14535
rect 4571 14532 4583 14535
rect 5166 14532 5172 14544
rect 4571 14504 5172 14532
rect 4571 14501 4583 14504
rect 4525 14495 4583 14501
rect 5166 14492 5172 14504
rect 5224 14532 5230 14544
rect 5276 14532 5304 14572
rect 5224 14504 5304 14532
rect 6569 14532 6597 14572
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 6914 14600 6920 14612
rect 6687 14572 6920 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 8110 14560 8116 14612
rect 8168 14560 8174 14612
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 8536 14572 9229 14600
rect 8536 14560 8542 14572
rect 9217 14569 9229 14572
rect 9263 14600 9275 14603
rect 10042 14600 10048 14612
rect 9263 14572 10048 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 10928 14572 11529 14600
rect 10928 14560 10934 14572
rect 11517 14569 11529 14572
rect 11563 14600 11575 14603
rect 13906 14600 13912 14612
rect 11563 14572 13912 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14274 14560 14280 14612
rect 14332 14560 14338 14612
rect 6569 14504 6684 14532
rect 5224 14492 5230 14504
rect 6656 14476 6684 14504
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9824 14504 9873 14532
rect 9824 14492 9830 14504
rect 9861 14501 9873 14504
rect 9907 14532 9919 14535
rect 13170 14532 13176 14544
rect 9907 14504 13176 14532
rect 9907 14501 9919 14504
rect 9861 14495 9919 14501
rect 13170 14492 13176 14504
rect 13228 14532 13234 14544
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 13228 14504 13369 14532
rect 13228 14492 13234 14504
rect 13357 14501 13369 14504
rect 13403 14501 13415 14535
rect 13357 14495 13415 14501
rect 1210 14424 1216 14476
rect 1268 14464 1274 14476
rect 1857 14467 1915 14473
rect 1857 14464 1869 14467
rect 1268 14436 1869 14464
rect 1268 14424 1274 14436
rect 1857 14433 1869 14436
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 3844 14436 4997 14464
rect 3844 14424 3850 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 4985 14427 5043 14433
rect 6638 14424 6644 14476
rect 6696 14424 6702 14476
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 3973 14399 4031 14405
rect 1627 14368 2774 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2746 14328 2774 14368
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4798 14396 4804 14408
rect 4019 14368 4804 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 6748 14396 6776 14427
rect 7006 14405 7012 14408
rect 7000 14396 7012 14405
rect 5316 14368 6776 14396
rect 6967 14368 7012 14396
rect 5316 14356 5322 14368
rect 5350 14328 5356 14340
rect 2746 14300 5356 14328
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 5528 14331 5586 14337
rect 5528 14297 5540 14331
rect 5574 14328 5586 14331
rect 6178 14328 6184 14340
rect 5574 14300 6184 14328
rect 5574 14297 5586 14300
rect 5528 14291 5586 14297
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 6748 14328 6776 14368
rect 7000 14359 7012 14368
rect 7006 14356 7012 14359
rect 7064 14356 7070 14408
rect 7558 14356 7564 14408
rect 7616 14356 7622 14408
rect 7576 14328 7604 14356
rect 6748 14300 7604 14328
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 7650 14260 7656 14272
rect 6144 14232 7656 14260
rect 6144 14220 6150 14232
rect 7650 14220 7656 14232
rect 7708 14260 7714 14272
rect 8110 14260 8116 14272
rect 7708 14232 8116 14260
rect 7708 14220 7714 14232
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 14550 14260 14556 14272
rect 13412 14232 14556 14260
rect 13412 14220 13418 14232
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 1104 14170 43884 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 43884 14170
rect 1104 14096 43884 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 1728 14028 2053 14056
rect 1728 14016 1734 14028
rect 2041 14025 2053 14028
rect 2087 14025 2099 14059
rect 2041 14019 2099 14025
rect 2498 14016 2504 14068
rect 2556 14056 2562 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 2556 14028 5181 14056
rect 2556 14016 2562 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 6178 14016 6184 14068
rect 6236 14016 6242 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 3234 13948 3240 14000
rect 3292 13988 3298 14000
rect 3329 13991 3387 13997
rect 3329 13988 3341 13991
rect 3292 13960 3341 13988
rect 3292 13948 3298 13960
rect 3329 13957 3341 13960
rect 3375 13988 3387 13991
rect 4065 13991 4123 13997
rect 4065 13988 4077 13991
rect 3375 13960 4077 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 4065 13957 4077 13960
rect 4111 13988 4123 13991
rect 4433 13991 4491 13997
rect 4433 13988 4445 13991
rect 4111 13960 4445 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 4433 13957 4445 13960
rect 4479 13988 4491 13991
rect 4614 13988 4620 14000
rect 4479 13960 4620 13988
rect 4479 13957 4491 13960
rect 4433 13951 4491 13957
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 4893 13991 4951 13997
rect 4893 13957 4905 13991
rect 4939 13988 4951 13991
rect 6086 13988 6092 14000
rect 4939 13960 6092 13988
rect 4939 13957 4951 13960
rect 4893 13951 4951 13957
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 3844 13892 5641 13920
rect 3844 13880 3850 13892
rect 5629 13889 5641 13892
rect 5675 13920 5687 13923
rect 5810 13920 5816 13932
rect 5675 13892 5816 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6380 13920 6408 14019
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 7098 14056 7104 14068
rect 6880 14028 7104 14056
rect 6880 14016 6886 14028
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 7834 14016 7840 14068
rect 7892 14016 7898 14068
rect 8110 14016 8116 14068
rect 8168 14016 8174 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8941 14059 8999 14065
rect 8941 14056 8953 14059
rect 8260 14028 8953 14056
rect 8260 14016 8266 14028
rect 8941 14025 8953 14028
rect 8987 14056 8999 14059
rect 10870 14056 10876 14068
rect 8987 14028 10876 14056
rect 8987 14025 8999 14028
rect 8941 14019 8999 14025
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 6972 13960 7236 13988
rect 6972 13948 6978 13960
rect 7208 13929 7236 13960
rect 6043 13892 6408 13920
rect 6733 13923 6791 13929
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7193 13923 7251 13929
rect 6779 13892 7144 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7116 13852 7144 13892
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 7852 13852 7880 14016
rect 7116 13824 7880 13852
rect 4614 13744 4620 13796
rect 4672 13744 4678 13796
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 7834 13784 7840 13796
rect 6788 13756 7840 13784
rect 6788 13744 6794 13756
rect 7834 13744 7840 13756
rect 7892 13784 7898 13796
rect 8573 13787 8631 13793
rect 8573 13784 8585 13787
rect 7892 13756 8585 13784
rect 7892 13744 7898 13756
rect 8573 13753 8585 13756
rect 8619 13753 8631 13787
rect 8573 13747 8631 13753
rect 4632 13716 4660 13744
rect 6914 13716 6920 13728
rect 4632 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13716 6978 13728
rect 7374 13716 7380 13728
rect 6972 13688 7380 13716
rect 6972 13676 6978 13688
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 1104 13626 43884 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 43884 13626
rect 1104 13552 43884 13574
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 3786 13512 3792 13524
rect 3651 13484 3792 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 3786 13472 3792 13484
rect 3844 13512 3850 13524
rect 4246 13512 4252 13524
rect 3844 13484 4252 13512
rect 3844 13472 3850 13484
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 4614 13472 4620 13524
rect 4672 13472 4678 13524
rect 5166 13472 5172 13524
rect 5224 13472 5230 13524
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13512 6055 13515
rect 6270 13512 6276 13524
rect 6043 13484 6276 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6411 13484 6929 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 6917 13481 6929 13484
rect 6963 13512 6975 13515
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 6963 13484 7481 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7469 13481 7481 13484
rect 7515 13512 7527 13515
rect 8478 13512 8484 13524
rect 7515 13484 8484 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 5537 13447 5595 13453
rect 5537 13413 5549 13447
rect 5583 13444 5595 13447
rect 6380 13444 6408 13475
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 5583 13416 6408 13444
rect 5583 13413 5595 13416
rect 5537 13407 5595 13413
rect 7374 13404 7380 13456
rect 7432 13444 7438 13456
rect 8113 13447 8171 13453
rect 8113 13444 8125 13447
rect 7432 13416 8125 13444
rect 7432 13404 7438 13416
rect 8113 13413 8125 13416
rect 8159 13413 8171 13447
rect 8113 13407 8171 13413
rect 1210 13336 1216 13388
rect 1268 13376 1274 13388
rect 1857 13379 1915 13385
rect 1857 13376 1869 13379
rect 1268 13348 1869 13376
rect 1268 13336 1274 13348
rect 1857 13345 1869 13348
rect 1903 13345 1915 13379
rect 1857 13339 1915 13345
rect 7834 13336 7840 13388
rect 7892 13336 7898 13388
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 4706 13308 4712 13320
rect 1627 13280 4712 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 1104 13082 43884 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 43884 13082
rect 1104 13008 43884 13030
rect 4246 12928 4252 12980
rect 4304 12928 4310 12980
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5224 12940 5917 12968
rect 5224 12928 5230 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6914 12968 6920 12980
rect 6687 12940 6920 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 5810 12860 5816 12912
rect 5868 12860 5874 12912
rect 6932 12900 6960 12928
rect 7653 12903 7711 12909
rect 7653 12900 7665 12903
rect 6932 12872 7665 12900
rect 7653 12869 7665 12872
rect 7699 12869 7711 12903
rect 7653 12863 7711 12869
rect 5828 12832 5856 12860
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 5828 12804 6929 12832
rect 6917 12801 6929 12804
rect 6963 12832 6975 12835
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6963 12804 7297 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 1104 12538 43884 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 43884 12538
rect 1104 12464 43884 12486
rect 1210 12248 1216 12300
rect 1268 12288 1274 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1268 12260 1869 12288
rect 1268 12248 1274 12260
rect 1857 12257 1869 12260
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12220 1639 12223
rect 6822 12220 6828 12232
rect 1627 12192 6828 12220
rect 1627 12189 1639 12192
rect 1581 12183 1639 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 1104 11994 43884 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 43884 11994
rect 1104 11920 43884 11942
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 11974 11744 11980 11756
rect 4672 11716 11980 11744
rect 4672 11704 4678 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 1104 11450 43884 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 43884 11450
rect 1104 11376 43884 11398
rect 1854 11160 1860 11212
rect 1912 11160 1918 11212
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 7742 11132 7748 11144
rect 1627 11104 7748 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 1104 10906 43884 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 43884 10906
rect 1104 10832 43884 10854
rect 1104 10362 43884 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 43884 10362
rect 1104 10288 43884 10310
rect 1210 10072 1216 10124
rect 1268 10112 1274 10124
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1268 10084 1869 10112
rect 1268 10072 1274 10084
rect 1857 10081 1869 10084
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 9398 10044 9404 10056
rect 1627 10016 9404 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 1104 9818 43884 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 43884 9818
rect 1104 9744 43884 9766
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 13354 9636 13360 9648
rect 11664 9608 13360 9636
rect 11664 9596 11670 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 1104 9274 43884 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 43884 9274
rect 1104 9200 43884 9222
rect 1210 8984 1216 9036
rect 1268 9024 1274 9036
rect 1857 9027 1915 9033
rect 1857 9024 1869 9027
rect 1268 8996 1869 9024
rect 1268 8984 1274 8996
rect 1857 8993 1869 8996
rect 1903 8993 1915 9027
rect 1857 8987 1915 8993
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 11146 8956 11152 8968
rect 1627 8928 11152 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 1104 8730 43884 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 43884 8730
rect 1104 8656 43884 8678
rect 1104 8186 43884 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 43884 8186
rect 1104 8112 43884 8134
rect 1210 7896 1216 7948
rect 1268 7936 1274 7948
rect 1857 7939 1915 7945
rect 1857 7936 1869 7939
rect 1268 7908 1869 7936
rect 1268 7896 1274 7908
rect 1857 7905 1869 7908
rect 1903 7905 1915 7939
rect 1857 7899 1915 7905
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 4614 7868 4620 7880
rect 1627 7840 4620 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 1104 7642 43884 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 43884 7642
rect 1104 7568 43884 7590
rect 1104 7098 43884 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 43884 7098
rect 1104 7024 43884 7046
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 1857 6851 1915 6857
rect 1857 6848 1869 6851
rect 1268 6820 1869 6848
rect 1268 6808 1274 6820
rect 1857 6817 1869 6820
rect 1903 6817 1915 6851
rect 1857 6811 1915 6817
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 11606 6780 11612 6792
rect 1627 6752 11612 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 1104 6554 43884 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 43884 6554
rect 1104 6480 43884 6502
rect 1104 6010 43884 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 43884 6010
rect 1104 5936 43884 5958
rect 1854 5720 1860 5772
rect 1912 5720 1918 5772
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1627 5664 3188 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 3160 5565 3188 5664
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 18506 5556 18512 5568
rect 3191 5528 18512 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 1104 5466 43884 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 43884 5466
rect 1104 5392 43884 5414
rect 1104 4922 43884 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 43884 4922
rect 1104 4848 43884 4870
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1857 4675 1915 4681
rect 1857 4672 1869 4675
rect 1268 4644 1869 4672
rect 1268 4632 1274 4644
rect 1857 4641 1869 4644
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 3160 4604 3188 4768
rect 1627 4576 3188 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1104 4378 43884 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 43884 4378
rect 1104 4304 43884 4326
rect 1104 3834 43884 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 43884 3834
rect 1104 3760 43884 3782
rect 3142 3680 3148 3732
rect 3200 3680 3206 3732
rect 1210 3544 1216 3596
rect 1268 3584 1274 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1268 3556 1869 3584
rect 1268 3544 1274 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 3160 3516 3188 3680
rect 1627 3488 3188 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1104 3290 43884 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 43884 3290
rect 1104 3216 43884 3238
rect 1104 2746 43884 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 43884 2746
rect 1104 2672 43884 2694
rect 24670 2592 24676 2644
rect 24728 2592 24734 2644
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 22741 2431 22799 2437
rect 22741 2397 22753 2431
rect 22787 2428 22799 2431
rect 24688 2428 24716 2592
rect 22787 2400 24716 2428
rect 22787 2397 22799 2400
rect 22741 2391 22799 2397
rect 1104 2202 43884 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 43884 2202
rect 1104 2128 43884 2150
<< via1 >>
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 24216 42304 24268 42356
rect 25412 42304 25464 42356
rect 26608 42304 26660 42356
rect 27804 42304 27856 42356
rect 29000 42304 29052 42356
rect 30196 42304 30248 42356
rect 31392 42304 31444 42356
rect 32588 42304 32640 42356
rect 36176 42304 36228 42356
rect 37372 42304 37424 42356
rect 34980 42236 35032 42288
rect 23940 42032 23992 42084
rect 24492 41964 24544 42016
rect 27344 41964 27396 42016
rect 27896 42007 27948 42016
rect 27896 41973 27905 42007
rect 27905 41973 27939 42007
rect 27939 41973 27948 42007
rect 27896 41964 27948 41973
rect 29092 42007 29144 42016
rect 29092 41973 29101 42007
rect 29101 41973 29135 42007
rect 29135 41973 29144 42007
rect 29092 41964 29144 41973
rect 31024 41964 31076 42016
rect 31484 42007 31536 42016
rect 31484 41973 31493 42007
rect 31493 41973 31527 42007
rect 31527 41973 31536 42007
rect 31484 41964 31536 41973
rect 32680 42007 32732 42016
rect 32680 41973 32689 42007
rect 32689 41973 32723 42007
rect 32723 41973 32732 42007
rect 32680 41964 32732 41973
rect 32772 41964 32824 42016
rect 36452 42007 36504 42016
rect 36452 41973 36461 42007
rect 36461 41973 36495 42007
rect 36495 41973 36504 42007
rect 36452 41964 36504 41973
rect 37648 42007 37700 42016
rect 37648 41973 37657 42007
rect 37657 41973 37691 42007
rect 37691 41973 37700 42007
rect 37648 41964 37700 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 17684 41760 17736 41812
rect 32772 41760 32824 41812
rect 940 41556 992 41608
rect 28724 41488 28776 41540
rect 29184 41420 29236 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 28816 41216 28868 41268
rect 29644 41216 29696 41268
rect 28356 41080 28408 41132
rect 8116 41055 8168 41064
rect 8116 41021 8125 41055
rect 8125 41021 8159 41055
rect 8159 41021 8168 41055
rect 8116 41012 8168 41021
rect 9128 41055 9180 41064
rect 9128 41021 9137 41055
rect 9137 41021 9171 41055
rect 9171 41021 9180 41055
rect 9128 41012 9180 41021
rect 10048 41055 10100 41064
rect 10048 41021 10057 41055
rect 10057 41021 10091 41055
rect 10091 41021 10100 41055
rect 10048 41012 10100 41021
rect 11152 41012 11204 41064
rect 12256 41055 12308 41064
rect 12256 41021 12265 41055
rect 12265 41021 12299 41055
rect 12299 41021 12308 41055
rect 12256 41012 12308 41021
rect 13544 41012 13596 41064
rect 27804 41012 27856 41064
rect 28724 41055 28776 41064
rect 28724 41021 28733 41055
rect 28733 41021 28767 41055
rect 28767 41021 28776 41055
rect 28724 41012 28776 41021
rect 28816 41055 28868 41064
rect 28816 41021 28825 41055
rect 28825 41021 28859 41055
rect 28859 41021 28868 41055
rect 28816 41012 28868 41021
rect 27712 40944 27764 40996
rect 29276 41055 29328 41064
rect 29276 41021 29285 41055
rect 29285 41021 29319 41055
rect 29319 41021 29328 41055
rect 29276 41012 29328 41021
rect 8668 40919 8720 40928
rect 8668 40885 8677 40919
rect 8677 40885 8711 40919
rect 8711 40885 8720 40919
rect 8668 40876 8720 40885
rect 9680 40876 9732 40928
rect 10600 40919 10652 40928
rect 10600 40885 10609 40919
rect 10609 40885 10643 40919
rect 10643 40885 10652 40919
rect 10600 40876 10652 40885
rect 11336 40919 11388 40928
rect 11336 40885 11345 40919
rect 11345 40885 11379 40919
rect 11379 40885 11388 40919
rect 11336 40876 11388 40885
rect 12808 40919 12860 40928
rect 12808 40885 12817 40919
rect 12817 40885 12851 40919
rect 12851 40885 12860 40919
rect 12808 40876 12860 40885
rect 12992 40876 13044 40928
rect 25044 40876 25096 40928
rect 28356 40919 28408 40928
rect 28356 40885 28365 40919
rect 28365 40885 28399 40919
rect 28399 40885 28408 40919
rect 28356 40876 28408 40885
rect 29460 40876 29512 40928
rect 29552 40876 29604 40928
rect 31208 40876 31260 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 12256 40672 12308 40724
rect 13268 40579 13320 40588
rect 13268 40545 13277 40579
rect 13277 40545 13311 40579
rect 13311 40545 13320 40579
rect 13268 40536 13320 40545
rect 23664 40536 23716 40588
rect 25044 40579 25096 40588
rect 25044 40545 25053 40579
rect 25053 40545 25087 40579
rect 25087 40545 25096 40579
rect 25044 40536 25096 40545
rect 940 40468 992 40520
rect 8576 40468 8628 40520
rect 8944 40511 8996 40520
rect 8944 40477 8953 40511
rect 8953 40477 8987 40511
rect 8987 40477 8996 40511
rect 8944 40468 8996 40477
rect 10416 40511 10468 40520
rect 10416 40477 10425 40511
rect 10425 40477 10459 40511
rect 10459 40477 10468 40511
rect 10416 40468 10468 40477
rect 11244 40511 11296 40520
rect 11244 40477 11253 40511
rect 11253 40477 11287 40511
rect 11287 40477 11296 40511
rect 11244 40468 11296 40477
rect 11888 40511 11940 40520
rect 11888 40477 11897 40511
rect 11897 40477 11931 40511
rect 11931 40477 11940 40511
rect 11888 40468 11940 40477
rect 14096 40511 14148 40520
rect 14096 40477 14105 40511
rect 14105 40477 14139 40511
rect 14139 40477 14148 40511
rect 14096 40468 14148 40477
rect 15108 40511 15160 40520
rect 15108 40477 15117 40511
rect 15117 40477 15151 40511
rect 15151 40477 15160 40511
rect 15108 40468 15160 40477
rect 15936 40511 15988 40520
rect 15936 40477 15945 40511
rect 15945 40477 15979 40511
rect 15979 40477 15988 40511
rect 15936 40468 15988 40477
rect 23480 40468 23532 40520
rect 24584 40511 24636 40520
rect 24584 40477 24593 40511
rect 24593 40477 24627 40511
rect 24627 40477 24636 40511
rect 24584 40468 24636 40477
rect 27896 40536 27948 40588
rect 29368 40672 29420 40724
rect 29736 40672 29788 40724
rect 8024 40400 8076 40452
rect 10876 40400 10928 40452
rect 24216 40443 24268 40452
rect 24216 40409 24225 40443
rect 24225 40409 24259 40443
rect 24259 40409 24268 40443
rect 24216 40400 24268 40409
rect 8852 40332 8904 40384
rect 10968 40375 11020 40384
rect 10968 40341 10977 40375
rect 10977 40341 11011 40375
rect 11011 40341 11020 40375
rect 10968 40332 11020 40341
rect 12440 40332 12492 40384
rect 13176 40332 13228 40384
rect 15752 40375 15804 40384
rect 15752 40341 15761 40375
rect 15761 40341 15795 40375
rect 15795 40341 15804 40375
rect 15752 40332 15804 40341
rect 16488 40375 16540 40384
rect 16488 40341 16497 40375
rect 16497 40341 16531 40375
rect 16531 40341 16540 40375
rect 16488 40332 16540 40341
rect 24768 40375 24820 40384
rect 24768 40341 24777 40375
rect 24777 40341 24811 40375
rect 24811 40341 24820 40375
rect 24768 40332 24820 40341
rect 26240 40400 26292 40452
rect 27436 40511 27488 40520
rect 27436 40477 27445 40511
rect 27445 40477 27479 40511
rect 27479 40477 27488 40511
rect 27436 40468 27488 40477
rect 29828 40536 29880 40588
rect 30104 40536 30156 40588
rect 29184 40511 29236 40520
rect 29184 40477 29193 40511
rect 29193 40477 29227 40511
rect 29227 40477 29236 40511
rect 29184 40468 29236 40477
rect 30748 40511 30800 40520
rect 30748 40477 30757 40511
rect 30757 40477 30791 40511
rect 30791 40477 30800 40511
rect 30748 40468 30800 40477
rect 31024 40511 31076 40520
rect 31024 40477 31033 40511
rect 31033 40477 31067 40511
rect 31067 40477 31076 40511
rect 31024 40468 31076 40477
rect 31484 40511 31536 40520
rect 31484 40477 31493 40511
rect 31493 40477 31527 40511
rect 31527 40477 31536 40511
rect 31484 40468 31536 40477
rect 26608 40332 26660 40384
rect 26700 40375 26752 40384
rect 26700 40341 26709 40375
rect 26709 40341 26743 40375
rect 26743 40341 26752 40375
rect 26700 40332 26752 40341
rect 27160 40375 27212 40384
rect 27160 40341 27169 40375
rect 27169 40341 27203 40375
rect 27203 40341 27212 40375
rect 27160 40332 27212 40341
rect 27620 40375 27672 40384
rect 27620 40341 27629 40375
rect 27629 40341 27663 40375
rect 27663 40341 27672 40375
rect 27620 40332 27672 40341
rect 27896 40375 27948 40384
rect 27896 40341 27905 40375
rect 27905 40341 27939 40375
rect 27939 40341 27948 40375
rect 27896 40332 27948 40341
rect 28816 40375 28868 40384
rect 28816 40341 28825 40375
rect 28825 40341 28859 40375
rect 28859 40341 28868 40375
rect 28816 40332 28868 40341
rect 29000 40332 29052 40384
rect 29368 40375 29420 40384
rect 29368 40341 29377 40375
rect 29377 40341 29411 40375
rect 29411 40341 29420 40375
rect 29368 40332 29420 40341
rect 29736 40332 29788 40384
rect 30380 40400 30432 40452
rect 30564 40332 30616 40384
rect 31300 40332 31352 40384
rect 31668 40375 31720 40384
rect 31668 40341 31677 40375
rect 31677 40341 31711 40375
rect 31711 40341 31720 40375
rect 31668 40332 31720 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 8116 40128 8168 40180
rect 10048 40128 10100 40180
rect 11336 40128 11388 40180
rect 14096 40128 14148 40180
rect 9588 40060 9640 40112
rect 12808 40060 12860 40112
rect 16488 40128 16540 40180
rect 27252 40128 27304 40180
rect 6276 39992 6328 40044
rect 8852 39992 8904 40044
rect 9496 39992 9548 40044
rect 13268 39992 13320 40044
rect 14740 39992 14792 40044
rect 6736 39924 6788 39976
rect 9220 39924 9272 39976
rect 9312 39967 9364 39976
rect 9312 39933 9321 39967
rect 9321 39933 9355 39967
rect 9355 39933 9364 39967
rect 9312 39924 9364 39933
rect 9404 39924 9456 39976
rect 10784 39924 10836 39976
rect 11980 39924 12032 39976
rect 7104 39831 7156 39840
rect 7104 39797 7113 39831
rect 7113 39797 7147 39831
rect 7147 39797 7156 39831
rect 7104 39788 7156 39797
rect 7840 39831 7892 39840
rect 7840 39797 7849 39831
rect 7849 39797 7883 39831
rect 7883 39797 7892 39831
rect 7840 39788 7892 39797
rect 9772 39788 9824 39840
rect 13636 39967 13688 39976
rect 13636 39933 13645 39967
rect 13645 39933 13679 39967
rect 13679 39933 13688 39967
rect 13636 39924 13688 39933
rect 15292 39924 15344 39976
rect 24216 40060 24268 40112
rect 24768 40060 24820 40112
rect 23940 40035 23992 40044
rect 23940 40001 23949 40035
rect 23949 40001 23983 40035
rect 23983 40001 23992 40035
rect 23940 39992 23992 40001
rect 26700 40060 26752 40112
rect 27620 40060 27672 40112
rect 27988 40060 28040 40112
rect 29644 40128 29696 40180
rect 30564 40128 30616 40180
rect 16856 39967 16908 39976
rect 16856 39933 16865 39967
rect 16865 39933 16899 39967
rect 16899 39933 16908 39967
rect 16856 39924 16908 39933
rect 17776 39967 17828 39976
rect 17776 39933 17785 39967
rect 17785 39933 17819 39967
rect 17819 39933 17828 39967
rect 17776 39924 17828 39933
rect 23480 39924 23532 39976
rect 26608 39992 26660 40044
rect 27436 39992 27488 40044
rect 29184 39992 29236 40044
rect 30380 39992 30432 40044
rect 13360 39788 13412 39840
rect 13820 39788 13872 39840
rect 15016 39831 15068 39840
rect 15016 39797 15025 39831
rect 15025 39797 15059 39831
rect 15059 39797 15068 39831
rect 15016 39788 15068 39797
rect 15568 39788 15620 39840
rect 17224 39788 17276 39840
rect 18328 39831 18380 39840
rect 18328 39797 18337 39831
rect 18337 39797 18371 39831
rect 18371 39797 18380 39831
rect 18328 39788 18380 39797
rect 23296 39788 23348 39840
rect 23664 39831 23716 39840
rect 23664 39797 23673 39831
rect 23673 39797 23707 39831
rect 23707 39797 23716 39831
rect 23664 39788 23716 39797
rect 24124 39831 24176 39840
rect 24124 39797 24133 39831
rect 24133 39797 24167 39831
rect 24167 39797 24176 39831
rect 24124 39788 24176 39797
rect 24492 39788 24544 39840
rect 25320 39788 25372 39840
rect 27528 39856 27580 39908
rect 28908 39924 28960 39976
rect 27436 39788 27488 39840
rect 27620 39788 27672 39840
rect 29092 39788 29144 39840
rect 30564 39856 30616 39908
rect 33232 39856 33284 39908
rect 33508 39788 33560 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1216 39448 1268 39500
rect 6368 39448 6420 39500
rect 9128 39584 9180 39636
rect 11152 39584 11204 39636
rect 13544 39627 13596 39636
rect 13544 39593 13553 39627
rect 13553 39593 13587 39627
rect 13587 39593 13596 39627
rect 13544 39584 13596 39593
rect 22376 39584 22428 39636
rect 7380 39491 7432 39500
rect 7380 39457 7389 39491
rect 7389 39457 7423 39491
rect 7423 39457 7432 39491
rect 7380 39448 7432 39457
rect 9772 39516 9824 39568
rect 6000 39423 6052 39432
rect 6000 39389 6009 39423
rect 6009 39389 6043 39423
rect 6043 39389 6052 39423
rect 6000 39380 6052 39389
rect 9680 39380 9732 39432
rect 9772 39380 9824 39432
rect 10600 39380 10652 39432
rect 11520 39423 11572 39432
rect 11520 39389 11529 39423
rect 11529 39389 11563 39423
rect 11563 39389 11572 39423
rect 11520 39380 11572 39389
rect 11980 39380 12032 39432
rect 12440 39423 12492 39432
rect 12440 39389 12474 39423
rect 12474 39389 12492 39423
rect 12440 39380 12492 39389
rect 14648 39423 14700 39432
rect 14648 39389 14657 39423
rect 14657 39389 14691 39423
rect 14691 39389 14700 39423
rect 14648 39380 14700 39389
rect 17132 39380 17184 39432
rect 17224 39380 17276 39432
rect 18144 39423 18196 39432
rect 18144 39389 18153 39423
rect 18153 39389 18187 39423
rect 18187 39389 18196 39423
rect 18144 39380 18196 39389
rect 24400 39423 24452 39432
rect 24400 39389 24409 39423
rect 24409 39389 24443 39423
rect 24443 39389 24452 39423
rect 24400 39380 24452 39389
rect 24492 39380 24544 39432
rect 26240 39584 26292 39636
rect 26332 39584 26384 39636
rect 27068 39516 27120 39568
rect 27620 39516 27672 39568
rect 25964 39448 26016 39500
rect 27896 39448 27948 39500
rect 28724 39448 28776 39500
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 26884 39380 26936 39432
rect 27068 39380 27120 39432
rect 27160 39380 27212 39432
rect 27252 39380 27304 39432
rect 6552 39287 6604 39296
rect 6552 39253 6561 39287
rect 6561 39253 6595 39287
rect 6595 39253 6604 39287
rect 6552 39244 6604 39253
rect 15752 39312 15804 39364
rect 9404 39287 9456 39296
rect 9404 39253 9413 39287
rect 9413 39253 9447 39287
rect 9447 39253 9456 39287
rect 9404 39244 9456 39253
rect 11336 39244 11388 39296
rect 12532 39244 12584 39296
rect 16028 39287 16080 39296
rect 16028 39253 16037 39287
rect 16037 39253 16071 39287
rect 16071 39253 16080 39287
rect 16028 39244 16080 39253
rect 16396 39287 16448 39296
rect 16396 39253 16405 39287
rect 16405 39253 16439 39287
rect 16439 39253 16448 39287
rect 22100 39355 22152 39364
rect 22100 39321 22109 39355
rect 22109 39321 22143 39355
rect 22143 39321 22152 39355
rect 22100 39312 22152 39321
rect 24124 39312 24176 39364
rect 24860 39312 24912 39364
rect 28908 39380 28960 39432
rect 31668 39380 31720 39432
rect 29368 39312 29420 39364
rect 43812 39312 43864 39364
rect 16396 39244 16448 39253
rect 17960 39287 18012 39296
rect 17960 39253 17969 39287
rect 17969 39253 18003 39287
rect 18003 39253 18012 39287
rect 17960 39244 18012 39253
rect 18696 39287 18748 39296
rect 18696 39253 18705 39287
rect 18705 39253 18739 39287
rect 18739 39253 18748 39287
rect 18696 39244 18748 39253
rect 21456 39287 21508 39296
rect 21456 39253 21465 39287
rect 21465 39253 21499 39287
rect 21499 39253 21508 39287
rect 21456 39244 21508 39253
rect 23204 39244 23256 39296
rect 23388 39244 23440 39296
rect 24308 39244 24360 39296
rect 25412 39244 25464 39296
rect 26240 39244 26292 39296
rect 27252 39244 27304 39296
rect 27344 39244 27396 39296
rect 28264 39244 28316 39296
rect 29184 39287 29236 39296
rect 29184 39253 29193 39287
rect 29193 39253 29227 39287
rect 29227 39253 29236 39287
rect 29184 39244 29236 39253
rect 30932 39287 30984 39296
rect 30932 39253 30941 39287
rect 30941 39253 30975 39287
rect 30975 39253 30984 39287
rect 30932 39244 30984 39253
rect 31944 39244 31996 39296
rect 32036 39244 32088 39296
rect 43536 39287 43588 39296
rect 43536 39253 43545 39287
rect 43545 39253 43579 39287
rect 43579 39253 43588 39287
rect 43536 39244 43588 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 6000 39040 6052 39092
rect 7104 39040 7156 39092
rect 8576 39040 8628 39092
rect 9680 39040 9732 39092
rect 11244 39083 11296 39092
rect 11244 39049 11253 39083
rect 11253 39049 11287 39083
rect 11287 39049 11296 39083
rect 11244 39040 11296 39049
rect 11520 39040 11572 39092
rect 11888 39083 11940 39092
rect 11888 39049 11897 39083
rect 11897 39049 11931 39083
rect 11931 39049 11940 39083
rect 11888 39040 11940 39049
rect 8668 38972 8720 39024
rect 9496 39015 9548 39024
rect 9496 38981 9505 39015
rect 9505 38981 9539 39015
rect 9539 38981 9548 39015
rect 9496 38972 9548 38981
rect 10968 38972 11020 39024
rect 13820 39040 13872 39092
rect 14096 39040 14148 39092
rect 15936 39040 15988 39092
rect 18144 39083 18196 39092
rect 18144 39049 18153 39083
rect 18153 39049 18187 39083
rect 18187 39049 18196 39083
rect 18144 39040 18196 39049
rect 18328 39040 18380 39092
rect 18696 39040 18748 39092
rect 24400 39040 24452 39092
rect 27252 39040 27304 39092
rect 12992 38972 13044 39024
rect 13176 39015 13228 39024
rect 13176 38981 13185 39015
rect 13185 38981 13219 39015
rect 13219 38981 13228 39015
rect 13176 38972 13228 38981
rect 13544 38972 13596 39024
rect 15016 38972 15068 39024
rect 23480 38972 23532 39024
rect 5632 38879 5684 38888
rect 5632 38845 5641 38879
rect 5641 38845 5675 38879
rect 5675 38845 5684 38879
rect 5632 38836 5684 38845
rect 5908 38836 5960 38888
rect 14648 38947 14700 38956
rect 14648 38913 14657 38947
rect 14657 38913 14691 38947
rect 14691 38913 14700 38947
rect 14648 38904 14700 38913
rect 17500 38904 17552 38956
rect 17960 38904 18012 38956
rect 19984 38904 20036 38956
rect 21364 38904 21416 38956
rect 21916 38904 21968 38956
rect 24308 38972 24360 39024
rect 24492 38972 24544 39024
rect 7380 38836 7432 38888
rect 9220 38836 9272 38888
rect 9496 38836 9548 38888
rect 9772 38836 9824 38888
rect 12348 38879 12400 38888
rect 12348 38845 12357 38879
rect 12357 38845 12391 38879
rect 12391 38845 12400 38879
rect 12348 38836 12400 38845
rect 13268 38879 13320 38888
rect 13268 38845 13277 38879
rect 13277 38845 13311 38879
rect 13311 38845 13320 38879
rect 13268 38836 13320 38845
rect 14280 38836 14332 38888
rect 17684 38836 17736 38888
rect 18788 38879 18840 38888
rect 18788 38845 18797 38879
rect 18797 38845 18831 38879
rect 18831 38845 18840 38879
rect 18788 38836 18840 38845
rect 21824 38879 21876 38888
rect 21824 38845 21833 38879
rect 21833 38845 21867 38879
rect 21867 38845 21876 38879
rect 21824 38836 21876 38845
rect 6184 38743 6236 38752
rect 6184 38709 6193 38743
rect 6193 38709 6227 38743
rect 6227 38709 6236 38743
rect 6184 38700 6236 38709
rect 7104 38700 7156 38752
rect 8208 38700 8260 38752
rect 11060 38700 11112 38752
rect 13360 38700 13412 38752
rect 15660 38700 15712 38752
rect 15844 38700 15896 38752
rect 16396 38743 16448 38752
rect 16396 38709 16405 38743
rect 16405 38709 16439 38743
rect 16439 38709 16448 38743
rect 16396 38700 16448 38709
rect 17776 38700 17828 38752
rect 19616 38743 19668 38752
rect 19616 38709 19625 38743
rect 19625 38709 19659 38743
rect 19659 38709 19668 38743
rect 19616 38700 19668 38709
rect 20260 38743 20312 38752
rect 20260 38709 20269 38743
rect 20269 38709 20303 38743
rect 20303 38709 20312 38743
rect 20260 38700 20312 38709
rect 20444 38700 20496 38752
rect 21272 38743 21324 38752
rect 21272 38709 21281 38743
rect 21281 38709 21315 38743
rect 21315 38709 21324 38743
rect 21272 38700 21324 38709
rect 21640 38743 21692 38752
rect 21640 38709 21649 38743
rect 21649 38709 21683 38743
rect 21683 38709 21692 38743
rect 21640 38700 21692 38709
rect 22100 38700 22152 38752
rect 23388 38836 23440 38888
rect 24584 38947 24636 38956
rect 24584 38913 24593 38947
rect 24593 38913 24627 38947
rect 24627 38913 24636 38947
rect 24584 38904 24636 38913
rect 24768 38947 24820 38956
rect 24768 38913 24777 38947
rect 24777 38913 24811 38947
rect 24811 38913 24820 38947
rect 24768 38904 24820 38913
rect 26884 38972 26936 39024
rect 29276 39040 29328 39092
rect 29368 39040 29420 39092
rect 29552 39040 29604 39092
rect 29644 39040 29696 39092
rect 30932 39040 30984 39092
rect 25412 38947 25464 38956
rect 25412 38913 25446 38947
rect 25446 38913 25464 38947
rect 23940 38836 23992 38888
rect 24216 38836 24268 38888
rect 23204 38700 23256 38752
rect 23480 38700 23532 38752
rect 25412 38904 25464 38913
rect 25964 38904 26016 38956
rect 27068 38904 27120 38956
rect 25320 38700 25372 38752
rect 27252 38904 27304 38956
rect 27528 38904 27580 38956
rect 28816 38836 28868 38888
rect 29368 38904 29420 38956
rect 29644 38904 29696 38956
rect 31208 38947 31260 38956
rect 31208 38913 31217 38947
rect 31217 38913 31251 38947
rect 31251 38913 31260 38947
rect 31208 38904 31260 38913
rect 31944 38904 31996 38956
rect 29920 38879 29972 38888
rect 29920 38845 29929 38879
rect 29929 38845 29963 38879
rect 29963 38845 29972 38879
rect 29920 38836 29972 38845
rect 29092 38700 29144 38752
rect 30840 38700 30892 38752
rect 31392 38768 31444 38820
rect 31576 38768 31628 38820
rect 33232 38768 33284 38820
rect 33600 38700 33652 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1216 38360 1268 38412
rect 6736 38496 6788 38548
rect 10232 38496 10284 38548
rect 10416 38496 10468 38548
rect 9220 38428 9272 38480
rect 11060 38496 11112 38548
rect 10784 38360 10836 38412
rect 12624 38496 12676 38548
rect 13636 38539 13688 38548
rect 13636 38505 13645 38539
rect 13645 38505 13679 38539
rect 13679 38505 13688 38539
rect 13636 38496 13688 38505
rect 15108 38496 15160 38548
rect 16856 38496 16908 38548
rect 17868 38496 17920 38548
rect 20168 38539 20220 38548
rect 20168 38505 20177 38539
rect 20177 38505 20211 38539
rect 20211 38505 20220 38539
rect 20168 38496 20220 38505
rect 21180 38496 21232 38548
rect 11980 38360 12032 38412
rect 12256 38403 12308 38412
rect 12256 38369 12265 38403
rect 12265 38369 12299 38403
rect 12299 38369 12308 38403
rect 12256 38360 12308 38369
rect 14188 38360 14240 38412
rect 15476 38360 15528 38412
rect 16028 38403 16080 38412
rect 16028 38369 16037 38403
rect 16037 38369 16071 38403
rect 16071 38369 16080 38403
rect 16028 38360 16080 38369
rect 17500 38360 17552 38412
rect 20260 38428 20312 38480
rect 20536 38428 20588 38480
rect 21548 38428 21600 38480
rect 24584 38496 24636 38548
rect 4160 38335 4212 38344
rect 4160 38301 4169 38335
rect 4169 38301 4203 38335
rect 4203 38301 4212 38335
rect 4160 38292 4212 38301
rect 4896 38335 4948 38344
rect 4896 38301 4905 38335
rect 4905 38301 4939 38335
rect 4939 38301 4948 38335
rect 4896 38292 4948 38301
rect 6552 38224 6604 38276
rect 7840 38292 7892 38344
rect 9036 38335 9088 38344
rect 9036 38301 9045 38335
rect 9045 38301 9079 38335
rect 9079 38301 9088 38335
rect 9036 38292 9088 38301
rect 7104 38224 7156 38276
rect 7472 38224 7524 38276
rect 10876 38335 10928 38344
rect 10876 38301 10885 38335
rect 10885 38301 10919 38335
rect 10919 38301 10928 38335
rect 10876 38292 10928 38301
rect 12532 38335 12584 38344
rect 12532 38301 12555 38335
rect 12555 38301 12584 38335
rect 11060 38224 11112 38276
rect 12532 38292 12584 38301
rect 13820 38292 13872 38344
rect 14372 38224 14424 38276
rect 18420 38335 18472 38344
rect 18420 38301 18429 38335
rect 18429 38301 18463 38335
rect 18463 38301 18472 38335
rect 18420 38292 18472 38301
rect 20720 38360 20772 38412
rect 23296 38428 23348 38480
rect 19616 38292 19668 38344
rect 22284 38403 22336 38412
rect 22284 38369 22293 38403
rect 22293 38369 22327 38403
rect 22327 38369 22336 38403
rect 22284 38360 22336 38369
rect 23664 38360 23716 38412
rect 29276 38496 29328 38548
rect 28724 38428 28776 38480
rect 31116 38496 31168 38548
rect 31576 38496 31628 38548
rect 14832 38224 14884 38276
rect 16856 38224 16908 38276
rect 17868 38224 17920 38276
rect 19984 38267 20036 38276
rect 19984 38233 19993 38267
rect 19993 38233 20027 38267
rect 20027 38233 20036 38267
rect 19984 38224 20036 38233
rect 4712 38199 4764 38208
rect 4712 38165 4721 38199
rect 4721 38165 4755 38199
rect 4755 38165 4764 38199
rect 4712 38156 4764 38165
rect 5448 38199 5500 38208
rect 5448 38165 5457 38199
rect 5457 38165 5491 38199
rect 5491 38165 5500 38199
rect 5448 38156 5500 38165
rect 6828 38156 6880 38208
rect 8760 38199 8812 38208
rect 8760 38165 8769 38199
rect 8769 38165 8803 38199
rect 8803 38165 8812 38199
rect 8760 38156 8812 38165
rect 9680 38199 9732 38208
rect 9680 38165 9689 38199
rect 9689 38165 9723 38199
rect 9723 38165 9732 38199
rect 9680 38156 9732 38165
rect 10416 38199 10468 38208
rect 10416 38165 10425 38199
rect 10425 38165 10459 38199
rect 10459 38165 10468 38199
rect 10416 38156 10468 38165
rect 12808 38156 12860 38208
rect 15108 38199 15160 38208
rect 15108 38165 15117 38199
rect 15117 38165 15151 38199
rect 15151 38165 15160 38199
rect 15108 38156 15160 38165
rect 15292 38156 15344 38208
rect 17684 38156 17736 38208
rect 18604 38156 18656 38208
rect 18696 38156 18748 38208
rect 20076 38156 20128 38208
rect 20352 38199 20404 38208
rect 20352 38165 20361 38199
rect 20361 38165 20395 38199
rect 20395 38165 20404 38199
rect 20352 38156 20404 38165
rect 21364 38335 21416 38344
rect 21364 38301 21373 38335
rect 21373 38301 21407 38335
rect 21407 38301 21416 38335
rect 21364 38292 21416 38301
rect 21272 38224 21324 38276
rect 21916 38292 21968 38344
rect 22192 38335 22244 38344
rect 22192 38301 22201 38335
rect 22201 38301 22235 38335
rect 22235 38301 22244 38335
rect 22192 38292 22244 38301
rect 23204 38292 23256 38344
rect 23480 38292 23532 38344
rect 24124 38292 24176 38344
rect 24492 38292 24544 38344
rect 28264 38360 28316 38412
rect 28908 38403 28960 38412
rect 28908 38369 28917 38403
rect 28917 38369 28951 38403
rect 28951 38369 28960 38403
rect 28908 38360 28960 38369
rect 30932 38428 30984 38480
rect 29368 38360 29420 38412
rect 30288 38360 30340 38412
rect 26148 38335 26200 38344
rect 26148 38301 26157 38335
rect 26157 38301 26191 38335
rect 26191 38301 26200 38335
rect 26148 38292 26200 38301
rect 26332 38292 26384 38344
rect 25412 38224 25464 38276
rect 21456 38156 21508 38208
rect 24032 38199 24084 38208
rect 24032 38165 24041 38199
rect 24041 38165 24075 38199
rect 24075 38165 24084 38199
rect 24032 38156 24084 38165
rect 25780 38199 25832 38208
rect 25780 38165 25789 38199
rect 25789 38165 25823 38199
rect 25823 38165 25832 38199
rect 25780 38156 25832 38165
rect 26516 38292 26568 38344
rect 27344 38335 27396 38344
rect 27344 38301 27353 38335
rect 27353 38301 27387 38335
rect 27387 38301 27396 38335
rect 27344 38292 27396 38301
rect 27528 38335 27580 38344
rect 27528 38301 27537 38335
rect 27537 38301 27571 38335
rect 27571 38301 27580 38335
rect 27528 38292 27580 38301
rect 28080 38335 28132 38344
rect 28080 38301 28089 38335
rect 28089 38301 28123 38335
rect 28123 38301 28132 38335
rect 28080 38292 28132 38301
rect 29184 38292 29236 38344
rect 27988 38267 28040 38276
rect 27988 38233 27997 38267
rect 27997 38233 28031 38267
rect 28031 38233 28040 38267
rect 27988 38224 28040 38233
rect 30012 38224 30064 38276
rect 30748 38292 30800 38344
rect 30840 38335 30892 38344
rect 30840 38301 30849 38335
rect 30849 38301 30883 38335
rect 30883 38301 30892 38335
rect 30840 38292 30892 38301
rect 31024 38335 31076 38344
rect 31024 38301 31033 38335
rect 31033 38301 31067 38335
rect 31067 38301 31076 38335
rect 31024 38292 31076 38301
rect 31116 38292 31168 38344
rect 37648 38360 37700 38412
rect 32312 38335 32364 38344
rect 32312 38301 32321 38335
rect 32321 38301 32355 38335
rect 32355 38301 32364 38335
rect 32312 38292 32364 38301
rect 32404 38292 32456 38344
rect 31944 38224 31996 38276
rect 32128 38267 32180 38276
rect 32128 38233 32137 38267
rect 32137 38233 32171 38267
rect 32171 38233 32180 38267
rect 32128 38224 32180 38233
rect 27160 38156 27212 38208
rect 31760 38156 31812 38208
rect 31852 38156 31904 38208
rect 32956 38199 33008 38208
rect 32956 38165 32965 38199
rect 32965 38165 32999 38199
rect 32999 38165 33008 38199
rect 32956 38156 33008 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4160 37952 4212 38004
rect 5632 37952 5684 38004
rect 6184 37952 6236 38004
rect 6736 37952 6788 38004
rect 6828 37927 6880 37936
rect 6828 37893 6837 37927
rect 6837 37893 6871 37927
rect 6871 37893 6880 37927
rect 6828 37884 6880 37893
rect 9312 37952 9364 38004
rect 9588 37952 9640 38004
rect 10416 37952 10468 38004
rect 11244 37952 11296 38004
rect 8024 37884 8076 37936
rect 8116 37884 8168 37936
rect 8300 37816 8352 37868
rect 10784 37816 10836 37868
rect 11796 37816 11848 37868
rect 12624 37859 12676 37868
rect 12624 37825 12633 37859
rect 12633 37825 12667 37859
rect 12667 37825 12676 37859
rect 12624 37816 12676 37825
rect 5264 37791 5316 37800
rect 5264 37757 5273 37791
rect 5273 37757 5307 37791
rect 5307 37757 5316 37791
rect 5264 37748 5316 37757
rect 5632 37680 5684 37732
rect 5908 37791 5960 37800
rect 5908 37757 5917 37791
rect 5917 37757 5951 37791
rect 5951 37757 5960 37791
rect 5908 37748 5960 37757
rect 6368 37748 6420 37800
rect 6920 37748 6972 37800
rect 7012 37791 7064 37800
rect 7012 37757 7021 37791
rect 7021 37757 7055 37791
rect 7055 37757 7064 37791
rect 7012 37748 7064 37757
rect 7472 37748 7524 37800
rect 8944 37748 8996 37800
rect 9404 37748 9456 37800
rect 6276 37612 6328 37664
rect 6460 37655 6512 37664
rect 6460 37621 6469 37655
rect 6469 37621 6503 37655
rect 6503 37621 6512 37655
rect 6460 37612 6512 37621
rect 10968 37791 11020 37800
rect 10968 37757 10977 37791
rect 10977 37757 11011 37791
rect 11011 37757 11020 37791
rect 10968 37748 11020 37757
rect 11152 37748 11204 37800
rect 12164 37791 12216 37800
rect 12164 37757 12173 37791
rect 12173 37757 12207 37791
rect 12207 37757 12216 37791
rect 12164 37748 12216 37757
rect 14648 37884 14700 37936
rect 12808 37816 12860 37868
rect 14924 37816 14976 37868
rect 16028 37952 16080 38004
rect 16212 37952 16264 38004
rect 15108 37884 15160 37936
rect 15384 37816 15436 37868
rect 15936 37816 15988 37868
rect 12256 37680 12308 37732
rect 15752 37791 15804 37800
rect 15752 37757 15761 37791
rect 15761 37757 15795 37791
rect 15795 37757 15804 37791
rect 15752 37748 15804 37757
rect 16212 37859 16264 37868
rect 16212 37825 16221 37859
rect 16221 37825 16255 37859
rect 16255 37825 16264 37859
rect 16212 37816 16264 37825
rect 16396 37748 16448 37800
rect 14464 37680 14516 37732
rect 17040 37859 17092 37868
rect 17040 37825 17049 37859
rect 17049 37825 17083 37859
rect 17083 37825 17092 37859
rect 17040 37816 17092 37825
rect 17132 37816 17184 37868
rect 18328 37952 18380 38004
rect 18696 37884 18748 37936
rect 19432 37884 19484 37936
rect 20076 37884 20128 37936
rect 20720 37952 20772 38004
rect 22376 37952 22428 38004
rect 24032 37952 24084 38004
rect 19248 37816 19300 37868
rect 16948 37748 17000 37800
rect 18420 37748 18472 37800
rect 18880 37748 18932 37800
rect 20168 37816 20220 37868
rect 20536 37816 20588 37868
rect 20720 37816 20772 37868
rect 17224 37723 17276 37732
rect 17224 37689 17233 37723
rect 17233 37689 17267 37723
rect 17267 37689 17276 37723
rect 17224 37680 17276 37689
rect 18328 37680 18380 37732
rect 22560 37816 22612 37868
rect 24860 37952 24912 38004
rect 25780 37952 25832 38004
rect 26148 37952 26200 38004
rect 28816 37995 28868 38004
rect 28816 37961 28825 37995
rect 28825 37961 28859 37995
rect 28859 37961 28868 37995
rect 28816 37952 28868 37961
rect 29644 37995 29696 38004
rect 29644 37961 29653 37995
rect 29653 37961 29687 37995
rect 29687 37961 29696 37995
rect 29644 37952 29696 37961
rect 24860 37816 24912 37868
rect 25044 37859 25096 37868
rect 25044 37825 25053 37859
rect 25053 37825 25087 37859
rect 25087 37825 25096 37859
rect 25044 37816 25096 37825
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 28448 37884 28500 37936
rect 32404 37952 32456 38004
rect 32956 37952 33008 38004
rect 33508 37995 33560 38004
rect 33508 37961 33517 37995
rect 33517 37961 33551 37995
rect 33551 37961 33560 37995
rect 33508 37952 33560 37961
rect 27436 37859 27488 37868
rect 27436 37825 27445 37859
rect 27445 37825 27479 37859
rect 27479 37825 27488 37859
rect 27436 37816 27488 37825
rect 27528 37816 27580 37868
rect 29092 37816 29144 37868
rect 29460 37816 29512 37868
rect 30288 37816 30340 37868
rect 30472 37859 30524 37868
rect 30472 37825 30506 37859
rect 30506 37825 30524 37859
rect 30472 37816 30524 37825
rect 33140 37816 33192 37868
rect 21364 37748 21416 37800
rect 21824 37748 21876 37800
rect 22100 37748 22152 37800
rect 9864 37612 9916 37664
rect 10416 37655 10468 37664
rect 10416 37621 10425 37655
rect 10425 37621 10459 37655
rect 10459 37621 10468 37655
rect 10416 37612 10468 37621
rect 11428 37612 11480 37664
rect 11520 37655 11572 37664
rect 11520 37621 11529 37655
rect 11529 37621 11563 37655
rect 11563 37621 11572 37655
rect 11520 37612 11572 37621
rect 13636 37612 13688 37664
rect 14096 37655 14148 37664
rect 14096 37621 14105 37655
rect 14105 37621 14139 37655
rect 14139 37621 14148 37655
rect 14096 37612 14148 37621
rect 14924 37612 14976 37664
rect 15200 37655 15252 37664
rect 15200 37621 15209 37655
rect 15209 37621 15243 37655
rect 15243 37621 15252 37655
rect 15200 37612 15252 37621
rect 15384 37612 15436 37664
rect 16488 37612 16540 37664
rect 16672 37612 16724 37664
rect 18512 37612 18564 37664
rect 18788 37612 18840 37664
rect 20536 37612 20588 37664
rect 20812 37680 20864 37732
rect 22192 37680 22244 37732
rect 25780 37748 25832 37800
rect 24216 37680 24268 37732
rect 26332 37748 26384 37800
rect 28908 37791 28960 37800
rect 28908 37757 28917 37791
rect 28917 37757 28951 37791
rect 28951 37757 28960 37791
rect 28908 37748 28960 37757
rect 21272 37612 21324 37664
rect 21548 37655 21600 37664
rect 21548 37621 21557 37655
rect 21557 37621 21591 37655
rect 21591 37621 21600 37655
rect 21548 37612 21600 37621
rect 23756 37612 23808 37664
rect 24768 37655 24820 37664
rect 24768 37621 24777 37655
rect 24777 37621 24811 37655
rect 24811 37621 24820 37655
rect 24768 37612 24820 37621
rect 25228 37612 25280 37664
rect 26240 37612 26292 37664
rect 26700 37612 26752 37664
rect 31208 37748 31260 37800
rect 32680 37748 32732 37800
rect 31300 37680 31352 37732
rect 27712 37612 27764 37664
rect 29552 37655 29604 37664
rect 29552 37621 29561 37655
rect 29561 37621 29595 37655
rect 29595 37621 29604 37655
rect 29552 37612 29604 37621
rect 30012 37612 30064 37664
rect 31852 37655 31904 37664
rect 31852 37621 31861 37655
rect 31861 37621 31895 37655
rect 31895 37621 31904 37655
rect 31852 37612 31904 37621
rect 32220 37612 32272 37664
rect 33232 37612 33284 37664
rect 33968 37655 34020 37664
rect 33968 37621 33977 37655
rect 33977 37621 34011 37655
rect 34011 37621 34020 37655
rect 33968 37612 34020 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5632 37408 5684 37460
rect 8392 37408 8444 37460
rect 9036 37408 9088 37460
rect 11060 37408 11112 37460
rect 6736 37315 6788 37324
rect 6736 37281 6745 37315
rect 6745 37281 6779 37315
rect 6779 37281 6788 37315
rect 6736 37272 6788 37281
rect 8484 37272 8536 37324
rect 1216 37068 1268 37120
rect 4160 37247 4212 37256
rect 4160 37213 4169 37247
rect 4169 37213 4203 37247
rect 4203 37213 4212 37247
rect 4160 37204 4212 37213
rect 7472 37204 7524 37256
rect 8576 37204 8628 37256
rect 4712 37136 4764 37188
rect 5724 37136 5776 37188
rect 5816 37068 5868 37120
rect 6092 37111 6144 37120
rect 6092 37077 6101 37111
rect 6101 37077 6135 37111
rect 6135 37077 6144 37111
rect 6092 37068 6144 37077
rect 6460 37136 6512 37188
rect 8668 37136 8720 37188
rect 9772 37204 9824 37256
rect 11336 37408 11388 37460
rect 12900 37408 12952 37460
rect 14004 37408 14056 37460
rect 11428 37340 11480 37392
rect 12164 37272 12216 37324
rect 13268 37340 13320 37392
rect 13912 37340 13964 37392
rect 14280 37451 14332 37460
rect 14280 37417 14289 37451
rect 14289 37417 14323 37451
rect 14323 37417 14332 37451
rect 14280 37408 14332 37417
rect 14464 37451 14516 37460
rect 14464 37417 14473 37451
rect 14473 37417 14507 37451
rect 14507 37417 14516 37451
rect 14464 37408 14516 37417
rect 17040 37408 17092 37460
rect 18052 37408 18104 37460
rect 17500 37383 17552 37392
rect 17500 37349 17509 37383
rect 17509 37349 17543 37383
rect 17543 37349 17552 37383
rect 17500 37340 17552 37349
rect 19800 37408 19852 37460
rect 13636 37315 13688 37324
rect 13636 37281 13645 37315
rect 13645 37281 13679 37315
rect 13679 37281 13688 37315
rect 13636 37272 13688 37281
rect 14188 37272 14240 37324
rect 14648 37315 14700 37324
rect 14648 37281 14657 37315
rect 14657 37281 14691 37315
rect 14691 37281 14700 37315
rect 14648 37272 14700 37281
rect 16488 37272 16540 37324
rect 11796 37204 11848 37256
rect 13176 37247 13228 37256
rect 13176 37213 13185 37247
rect 13185 37213 13219 37247
rect 13219 37213 13228 37247
rect 13176 37204 13228 37213
rect 13360 37204 13412 37256
rect 14924 37247 14976 37256
rect 14924 37213 14958 37247
rect 14958 37213 14976 37247
rect 9680 37136 9732 37188
rect 10968 37136 11020 37188
rect 11060 37136 11112 37188
rect 14924 37204 14976 37213
rect 6644 37111 6696 37120
rect 6644 37077 6653 37111
rect 6653 37077 6687 37111
rect 6687 37077 6696 37111
rect 6644 37068 6696 37077
rect 8944 37111 8996 37120
rect 8944 37077 8953 37111
rect 8953 37077 8987 37111
rect 8987 37077 8996 37111
rect 8944 37068 8996 37077
rect 9404 37111 9456 37120
rect 9404 37077 9413 37111
rect 9413 37077 9447 37111
rect 9447 37077 9456 37111
rect 9404 37068 9456 37077
rect 11336 37111 11388 37120
rect 11336 37077 11345 37111
rect 11345 37077 11379 37111
rect 11379 37077 11388 37111
rect 11336 37068 11388 37077
rect 11888 37068 11940 37120
rect 12164 37111 12216 37120
rect 12164 37077 12173 37111
rect 12173 37077 12207 37111
rect 12207 37077 12216 37111
rect 12164 37068 12216 37077
rect 12532 37111 12584 37120
rect 12532 37077 12541 37111
rect 12541 37077 12575 37111
rect 12575 37077 12584 37111
rect 12532 37068 12584 37077
rect 12992 37111 13044 37120
rect 12992 37077 13001 37111
rect 13001 37077 13035 37111
rect 13035 37077 13044 37111
rect 12992 37068 13044 37077
rect 13176 37068 13228 37120
rect 14556 37136 14608 37188
rect 14832 37068 14884 37120
rect 16304 37068 16356 37120
rect 16488 37068 16540 37120
rect 19248 37272 19300 37324
rect 29552 37408 29604 37460
rect 20444 37272 20496 37324
rect 21548 37272 21600 37324
rect 17224 37204 17276 37256
rect 17592 37204 17644 37256
rect 18788 37204 18840 37256
rect 16856 37136 16908 37188
rect 17040 37136 17092 37188
rect 17408 37136 17460 37188
rect 17868 37068 17920 37120
rect 17960 37068 18012 37120
rect 19800 37204 19852 37256
rect 19248 37136 19300 37188
rect 24216 37340 24268 37392
rect 25228 37340 25280 37392
rect 26240 37340 26292 37392
rect 28724 37340 28776 37392
rect 33140 37408 33192 37460
rect 33600 37451 33652 37460
rect 33600 37417 33609 37451
rect 33609 37417 33643 37451
rect 33643 37417 33652 37451
rect 33600 37408 33652 37417
rect 23296 37272 23348 37324
rect 24768 37315 24820 37324
rect 24768 37281 24777 37315
rect 24777 37281 24811 37315
rect 24811 37281 24820 37315
rect 24768 37272 24820 37281
rect 19156 37068 19208 37120
rect 20812 37111 20864 37120
rect 20812 37077 20821 37111
rect 20821 37077 20855 37111
rect 20855 37077 20864 37111
rect 20812 37068 20864 37077
rect 20996 37068 21048 37120
rect 21732 37068 21784 37120
rect 22284 37204 22336 37256
rect 22468 37136 22520 37188
rect 22836 37179 22888 37188
rect 22836 37145 22845 37179
rect 22845 37145 22879 37179
rect 22879 37145 22888 37179
rect 22836 37136 22888 37145
rect 23848 37136 23900 37188
rect 24032 37247 24084 37256
rect 24032 37213 24041 37247
rect 24041 37213 24075 37247
rect 24075 37213 24084 37247
rect 24032 37204 24084 37213
rect 24124 37247 24176 37256
rect 24124 37213 24133 37247
rect 24133 37213 24167 37247
rect 24167 37213 24176 37247
rect 24124 37204 24176 37213
rect 24400 37204 24452 37256
rect 24216 37136 24268 37188
rect 24952 37247 25004 37256
rect 24952 37213 24961 37247
rect 24961 37213 24995 37247
rect 24995 37213 25004 37247
rect 24952 37204 25004 37213
rect 22284 37068 22336 37120
rect 22560 37068 22612 37120
rect 23112 37068 23164 37120
rect 23572 37111 23624 37120
rect 23572 37077 23581 37111
rect 23581 37077 23615 37111
rect 23615 37077 23624 37111
rect 23572 37068 23624 37077
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 25044 37068 25096 37120
rect 27436 37272 27488 37324
rect 29276 37272 29328 37324
rect 29552 37272 29604 37324
rect 26700 37204 26752 37256
rect 26792 37247 26844 37256
rect 26792 37213 26801 37247
rect 26801 37213 26835 37247
rect 26835 37213 26844 37247
rect 26792 37204 26844 37213
rect 26976 37204 27028 37256
rect 29644 37204 29696 37256
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 31208 37272 31260 37324
rect 30932 37204 30984 37256
rect 31116 37247 31168 37256
rect 31116 37213 31125 37247
rect 31125 37213 31159 37247
rect 31159 37213 31168 37247
rect 31116 37204 31168 37213
rect 31392 37204 31444 37256
rect 26516 37068 26568 37120
rect 26608 37111 26660 37120
rect 26608 37077 26617 37111
rect 26617 37077 26651 37111
rect 26651 37077 26660 37111
rect 26608 37068 26660 37077
rect 27068 37068 27120 37120
rect 27620 37068 27672 37120
rect 30012 37136 30064 37188
rect 33968 37204 34020 37256
rect 29276 37068 29328 37120
rect 30380 37068 30432 37120
rect 31116 37068 31168 37120
rect 32036 37068 32088 37120
rect 33324 37111 33376 37120
rect 33324 37077 33333 37111
rect 33333 37077 33367 37111
rect 33367 37077 33376 37111
rect 33324 37068 33376 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 5448 36796 5500 36848
rect 6644 36864 6696 36916
rect 9680 36864 9732 36916
rect 11336 36864 11388 36916
rect 4160 36771 4212 36780
rect 4160 36737 4169 36771
rect 4169 36737 4203 36771
rect 4203 36737 4212 36771
rect 4160 36728 4212 36737
rect 5632 36728 5684 36780
rect 6644 36660 6696 36712
rect 7012 36728 7064 36780
rect 8208 36728 8260 36780
rect 9588 36728 9640 36780
rect 9772 36771 9824 36780
rect 9772 36737 9781 36771
rect 9781 36737 9815 36771
rect 9815 36737 9824 36771
rect 9772 36728 9824 36737
rect 11060 36728 11112 36780
rect 11520 36796 11572 36848
rect 12992 36864 13044 36916
rect 13544 36864 13596 36916
rect 14556 36864 14608 36916
rect 13912 36796 13964 36848
rect 13360 36728 13412 36780
rect 7104 36592 7156 36644
rect 8116 36660 8168 36712
rect 9496 36660 9548 36712
rect 12072 36703 12124 36712
rect 4068 36567 4120 36576
rect 4068 36533 4077 36567
rect 4077 36533 4111 36567
rect 4111 36533 4120 36567
rect 4068 36524 4120 36533
rect 6092 36567 6144 36576
rect 6092 36533 6101 36567
rect 6101 36533 6135 36567
rect 6135 36533 6144 36567
rect 6092 36524 6144 36533
rect 6736 36524 6788 36576
rect 8760 36524 8812 36576
rect 9036 36524 9088 36576
rect 12072 36669 12081 36703
rect 12081 36669 12115 36703
rect 12115 36669 12124 36703
rect 12072 36660 12124 36669
rect 12624 36660 12676 36712
rect 14096 36771 14148 36780
rect 14096 36737 14105 36771
rect 14105 36737 14139 36771
rect 14139 36737 14148 36771
rect 14096 36728 14148 36737
rect 17592 36864 17644 36916
rect 17960 36864 18012 36916
rect 18420 36864 18472 36916
rect 19156 36864 19208 36916
rect 16856 36796 16908 36848
rect 13636 36592 13688 36644
rect 14556 36660 14608 36712
rect 11520 36567 11572 36576
rect 11520 36533 11529 36567
rect 11529 36533 11563 36567
rect 11563 36533 11572 36567
rect 11520 36524 11572 36533
rect 11888 36524 11940 36576
rect 13176 36567 13228 36576
rect 13176 36533 13185 36567
rect 13185 36533 13219 36567
rect 13219 36533 13228 36567
rect 13176 36524 13228 36533
rect 13912 36567 13964 36576
rect 13912 36533 13921 36567
rect 13921 36533 13955 36567
rect 13955 36533 13964 36567
rect 13912 36524 13964 36533
rect 14924 36660 14976 36712
rect 15752 36728 15804 36780
rect 15844 36728 15896 36780
rect 16488 36728 16540 36780
rect 14924 36524 14976 36576
rect 16304 36660 16356 36712
rect 17224 36703 17276 36712
rect 17224 36669 17233 36703
rect 17233 36669 17267 36703
rect 17267 36669 17276 36703
rect 17224 36660 17276 36669
rect 17408 36728 17460 36780
rect 20812 36864 20864 36916
rect 22192 36864 22244 36916
rect 22836 36864 22888 36916
rect 24584 36864 24636 36916
rect 21640 36796 21692 36848
rect 24860 36796 24912 36848
rect 18604 36703 18656 36712
rect 18604 36669 18613 36703
rect 18613 36669 18647 36703
rect 18647 36669 18656 36703
rect 18604 36660 18656 36669
rect 18696 36703 18748 36712
rect 18696 36669 18705 36703
rect 18705 36669 18739 36703
rect 18739 36669 18748 36703
rect 18696 36660 18748 36669
rect 15660 36592 15712 36644
rect 17132 36592 17184 36644
rect 17960 36592 18012 36644
rect 19248 36703 19300 36712
rect 19248 36669 19257 36703
rect 19257 36669 19291 36703
rect 19291 36669 19300 36703
rect 19248 36660 19300 36669
rect 21456 36703 21508 36712
rect 21456 36669 21465 36703
rect 21465 36669 21499 36703
rect 21499 36669 21508 36703
rect 21456 36660 21508 36669
rect 19156 36592 19208 36644
rect 18512 36524 18564 36576
rect 19340 36524 19392 36576
rect 20352 36524 20404 36576
rect 20628 36567 20680 36576
rect 20628 36533 20637 36567
rect 20637 36533 20671 36567
rect 20671 36533 20680 36567
rect 20628 36524 20680 36533
rect 23112 36771 23164 36780
rect 23112 36737 23121 36771
rect 23121 36737 23155 36771
rect 23155 36737 23164 36771
rect 23112 36728 23164 36737
rect 23204 36728 23256 36780
rect 26976 36796 27028 36848
rect 26240 36728 26292 36780
rect 26424 36771 26476 36780
rect 26424 36737 26433 36771
rect 26433 36737 26467 36771
rect 26467 36737 26476 36771
rect 26424 36728 26476 36737
rect 24400 36660 24452 36712
rect 26332 36635 26384 36644
rect 26332 36601 26341 36635
rect 26341 36601 26375 36635
rect 26375 36601 26384 36635
rect 26792 36728 26844 36780
rect 27160 36728 27212 36780
rect 26332 36592 26384 36601
rect 27620 36771 27672 36780
rect 27620 36737 27629 36771
rect 27629 36737 27663 36771
rect 27663 36737 27672 36771
rect 27620 36728 27672 36737
rect 27712 36703 27764 36712
rect 27712 36669 27721 36703
rect 27721 36669 27755 36703
rect 27755 36669 27764 36703
rect 27712 36660 27764 36669
rect 28080 36771 28132 36780
rect 28080 36737 28089 36771
rect 28089 36737 28123 36771
rect 28123 36737 28132 36771
rect 28080 36728 28132 36737
rect 28356 36728 28408 36780
rect 28632 36771 28684 36780
rect 28632 36737 28641 36771
rect 28641 36737 28675 36771
rect 28675 36737 28684 36771
rect 28632 36728 28684 36737
rect 29184 36796 29236 36848
rect 29736 36864 29788 36916
rect 30196 36864 30248 36916
rect 33140 36907 33192 36916
rect 33140 36873 33149 36907
rect 33149 36873 33183 36907
rect 33183 36873 33192 36907
rect 33140 36864 33192 36873
rect 33232 36864 33284 36916
rect 28540 36660 28592 36712
rect 29000 36728 29052 36780
rect 29368 36771 29420 36780
rect 29368 36737 29377 36771
rect 29377 36737 29411 36771
rect 29411 36737 29420 36771
rect 29368 36728 29420 36737
rect 29460 36771 29512 36780
rect 29460 36737 29469 36771
rect 29469 36737 29503 36771
rect 29503 36737 29512 36771
rect 29460 36728 29512 36737
rect 31300 36796 31352 36848
rect 30012 36771 30064 36780
rect 30012 36737 30021 36771
rect 30021 36737 30055 36771
rect 30055 36737 30064 36771
rect 30012 36728 30064 36737
rect 23664 36524 23716 36576
rect 24308 36524 24360 36576
rect 25872 36524 25924 36576
rect 28908 36592 28960 36644
rect 29000 36524 29052 36576
rect 29092 36567 29144 36576
rect 29092 36533 29101 36567
rect 29101 36533 29135 36567
rect 29135 36533 29144 36567
rect 29092 36524 29144 36533
rect 29736 36592 29788 36644
rect 31760 36660 31812 36712
rect 30380 36524 30432 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4068 36320 4120 36372
rect 4896 36320 4948 36372
rect 5632 36320 5684 36372
rect 8484 36320 8536 36372
rect 10968 36363 11020 36372
rect 10968 36329 10977 36363
rect 10977 36329 11011 36363
rect 11011 36329 11020 36363
rect 10968 36320 11020 36329
rect 11060 36320 11112 36372
rect 940 36116 992 36168
rect 4436 36159 4488 36168
rect 4436 36125 4445 36159
rect 4445 36125 4479 36159
rect 4479 36125 4488 36159
rect 4436 36116 4488 36125
rect 5632 36227 5684 36236
rect 5632 36193 5641 36227
rect 5641 36193 5675 36227
rect 5675 36193 5684 36227
rect 5632 36184 5684 36193
rect 6000 36159 6052 36168
rect 6000 36125 6009 36159
rect 6009 36125 6043 36159
rect 6043 36125 6052 36159
rect 6000 36116 6052 36125
rect 5908 36048 5960 36100
rect 9036 36252 9088 36304
rect 9772 36252 9824 36304
rect 7656 36184 7708 36236
rect 7380 36116 7432 36168
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 8116 36159 8168 36168
rect 8116 36125 8125 36159
rect 8125 36125 8159 36159
rect 8159 36125 8168 36159
rect 8116 36116 8168 36125
rect 9036 36116 9088 36168
rect 9312 36159 9364 36168
rect 9312 36125 9321 36159
rect 9321 36125 9355 36159
rect 9355 36125 9364 36159
rect 9312 36116 9364 36125
rect 10416 36227 10468 36236
rect 10416 36193 10425 36227
rect 10425 36193 10459 36227
rect 10459 36193 10468 36227
rect 10416 36184 10468 36193
rect 12164 36320 12216 36372
rect 13360 36363 13412 36372
rect 13360 36329 13369 36363
rect 13369 36329 13403 36363
rect 13403 36329 13412 36363
rect 13360 36320 13412 36329
rect 13912 36320 13964 36372
rect 11980 36227 12032 36236
rect 11980 36193 11989 36227
rect 11989 36193 12023 36227
rect 12023 36193 12032 36227
rect 11980 36184 12032 36193
rect 6920 36048 6972 36100
rect 12072 36116 12124 36168
rect 13820 36116 13872 36168
rect 16212 36320 16264 36372
rect 16856 36320 16908 36372
rect 17316 36320 17368 36372
rect 19248 36363 19300 36372
rect 19248 36329 19257 36363
rect 19257 36329 19291 36363
rect 19291 36329 19300 36363
rect 19248 36320 19300 36329
rect 20260 36320 20312 36372
rect 22468 36363 22520 36372
rect 22468 36329 22477 36363
rect 22477 36329 22511 36363
rect 22511 36329 22520 36363
rect 22468 36320 22520 36329
rect 25872 36320 25924 36372
rect 26608 36320 26660 36372
rect 14740 36227 14792 36236
rect 14740 36193 14749 36227
rect 14749 36193 14783 36227
rect 14783 36193 14792 36227
rect 14740 36184 14792 36193
rect 15660 36227 15712 36236
rect 15660 36193 15669 36227
rect 15669 36193 15703 36227
rect 15703 36193 15712 36227
rect 15660 36184 15712 36193
rect 10140 36048 10192 36100
rect 10968 36048 11020 36100
rect 13728 36048 13780 36100
rect 16120 36116 16172 36168
rect 16948 36184 17000 36236
rect 17776 36116 17828 36168
rect 17960 36159 18012 36168
rect 17960 36125 17969 36159
rect 17969 36125 18003 36159
rect 18003 36125 18012 36159
rect 17960 36116 18012 36125
rect 18512 36159 18564 36168
rect 18512 36125 18521 36159
rect 18521 36125 18555 36159
rect 18555 36125 18564 36159
rect 18512 36116 18564 36125
rect 18604 36116 18656 36168
rect 15384 36048 15436 36100
rect 17040 36048 17092 36100
rect 17500 36048 17552 36100
rect 22100 36184 22152 36236
rect 25596 36252 25648 36304
rect 24308 36184 24360 36236
rect 25964 36184 26016 36236
rect 21456 36116 21508 36168
rect 21824 36159 21876 36168
rect 21824 36125 21833 36159
rect 21833 36125 21867 36159
rect 21867 36125 21876 36159
rect 21824 36116 21876 36125
rect 24768 36116 24820 36168
rect 25044 36159 25096 36168
rect 25044 36125 25053 36159
rect 25053 36125 25087 36159
rect 25087 36125 25096 36159
rect 25044 36116 25096 36125
rect 20628 36048 20680 36100
rect 25320 36048 25372 36100
rect 25412 36048 25464 36100
rect 26332 36048 26384 36100
rect 26700 36227 26752 36236
rect 26700 36193 26709 36227
rect 26709 36193 26743 36227
rect 26743 36193 26752 36227
rect 26700 36184 26752 36193
rect 28080 36320 28132 36372
rect 28172 36320 28224 36372
rect 28724 36320 28776 36372
rect 4988 36023 5040 36032
rect 4988 35989 4997 36023
rect 4997 35989 5031 36023
rect 5031 35989 5040 36023
rect 4988 35980 5040 35989
rect 6552 36023 6604 36032
rect 6552 35989 6561 36023
rect 6561 35989 6595 36023
rect 6595 35989 6604 36023
rect 6552 35980 6604 35989
rect 7288 36023 7340 36032
rect 7288 35989 7297 36023
rect 7297 35989 7331 36023
rect 7331 35989 7340 36023
rect 7288 35980 7340 35989
rect 8760 36023 8812 36032
rect 8760 35989 8769 36023
rect 8769 35989 8803 36023
rect 8803 35989 8812 36023
rect 8760 35980 8812 35989
rect 9496 35980 9548 36032
rect 12808 35980 12860 36032
rect 13084 35980 13136 36032
rect 13452 36023 13504 36032
rect 13452 35989 13461 36023
rect 13461 35989 13495 36023
rect 13495 35989 13504 36023
rect 13452 35980 13504 35989
rect 13820 36023 13872 36032
rect 13820 35989 13829 36023
rect 13829 35989 13863 36023
rect 13863 35989 13872 36023
rect 13820 35980 13872 35989
rect 14280 35980 14332 36032
rect 16212 35980 16264 36032
rect 17408 36023 17460 36032
rect 17408 35989 17417 36023
rect 17417 35989 17451 36023
rect 17451 35989 17460 36023
rect 17408 35980 17460 35989
rect 18144 35980 18196 36032
rect 20168 35980 20220 36032
rect 21732 35980 21784 36032
rect 25504 35980 25556 36032
rect 26056 36023 26108 36032
rect 26056 35989 26065 36023
rect 26065 35989 26099 36023
rect 26099 35989 26108 36023
rect 26056 35980 26108 35989
rect 26424 36023 26476 36032
rect 26424 35989 26433 36023
rect 26433 35989 26467 36023
rect 26467 35989 26476 36023
rect 26424 35980 26476 35989
rect 26976 36048 27028 36100
rect 28816 36252 28868 36304
rect 28448 36227 28500 36236
rect 28448 36193 28457 36227
rect 28457 36193 28491 36227
rect 28491 36193 28500 36227
rect 28448 36184 28500 36193
rect 28540 36227 28592 36236
rect 28540 36193 28549 36227
rect 28549 36193 28583 36227
rect 28583 36193 28592 36227
rect 28540 36184 28592 36193
rect 28632 36184 28684 36236
rect 28908 36184 28960 36236
rect 29460 36320 29512 36372
rect 29736 36320 29788 36372
rect 32128 36184 32180 36236
rect 33048 36184 33100 36236
rect 29092 36159 29144 36168
rect 29092 36125 29101 36159
rect 29101 36125 29135 36159
rect 29135 36125 29144 36159
rect 29092 36116 29144 36125
rect 27896 35980 27948 36032
rect 27988 36023 28040 36032
rect 27988 35989 27997 36023
rect 27997 35989 28031 36023
rect 28031 35989 28040 36023
rect 27988 35980 28040 35989
rect 28356 36023 28408 36032
rect 28356 35989 28365 36023
rect 28365 35989 28399 36023
rect 28399 35989 28408 36023
rect 28356 35980 28408 35989
rect 28540 35980 28592 36032
rect 28724 35980 28776 36032
rect 30104 36116 30156 36168
rect 30288 36116 30340 36168
rect 32312 36091 32364 36100
rect 32312 36057 32321 36091
rect 32321 36057 32355 36091
rect 32355 36057 32364 36091
rect 32312 36048 32364 36057
rect 30380 35980 30432 36032
rect 31944 36023 31996 36032
rect 31944 35989 31953 36023
rect 31953 35989 31987 36023
rect 31987 35989 31996 36023
rect 31944 35980 31996 35989
rect 32680 36023 32732 36032
rect 32680 35989 32689 36023
rect 32689 35989 32723 36023
rect 32723 35989 32732 36023
rect 32680 35980 32732 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4436 35776 4488 35828
rect 6000 35776 6052 35828
rect 7288 35776 7340 35828
rect 7380 35776 7432 35828
rect 7472 35776 7524 35828
rect 8116 35776 8168 35828
rect 8760 35776 8812 35828
rect 9404 35776 9456 35828
rect 12532 35819 12584 35828
rect 12532 35785 12541 35819
rect 12541 35785 12575 35819
rect 12575 35785 12584 35819
rect 12532 35776 12584 35785
rect 12624 35819 12676 35828
rect 12624 35785 12633 35819
rect 12633 35785 12667 35819
rect 12667 35785 12676 35819
rect 12624 35776 12676 35785
rect 13176 35776 13228 35828
rect 13728 35776 13780 35828
rect 13820 35776 13872 35828
rect 16396 35776 16448 35828
rect 18328 35776 18380 35828
rect 5632 35708 5684 35760
rect 5264 35615 5316 35624
rect 5264 35581 5273 35615
rect 5273 35581 5307 35615
rect 5307 35581 5316 35615
rect 5264 35572 5316 35581
rect 5908 35615 5960 35624
rect 5908 35581 5917 35615
rect 5917 35581 5951 35615
rect 5951 35581 5960 35615
rect 5908 35572 5960 35581
rect 7748 35708 7800 35760
rect 8300 35708 8352 35760
rect 6276 35504 6328 35556
rect 7012 35615 7064 35624
rect 7012 35581 7021 35615
rect 7021 35581 7055 35615
rect 7055 35581 7064 35615
rect 7012 35572 7064 35581
rect 8852 35640 8904 35692
rect 9036 35640 9088 35692
rect 10140 35708 10192 35760
rect 11336 35708 11388 35760
rect 8024 35572 8076 35624
rect 9404 35572 9456 35624
rect 9680 35640 9732 35692
rect 9772 35683 9824 35692
rect 9772 35649 9781 35683
rect 9781 35649 9815 35683
rect 9815 35649 9824 35683
rect 9772 35640 9824 35649
rect 11152 35683 11204 35692
rect 11152 35649 11161 35683
rect 11161 35649 11195 35683
rect 11195 35649 11204 35683
rect 11152 35640 11204 35649
rect 11888 35683 11940 35692
rect 11888 35649 11897 35683
rect 11897 35649 11931 35683
rect 11931 35649 11940 35683
rect 11888 35640 11940 35649
rect 12716 35708 12768 35760
rect 14648 35708 14700 35760
rect 14004 35640 14056 35692
rect 16212 35708 16264 35760
rect 18512 35776 18564 35828
rect 21824 35776 21876 35828
rect 23204 35819 23256 35828
rect 23204 35785 23213 35819
rect 23213 35785 23247 35819
rect 23247 35785 23256 35819
rect 23204 35776 23256 35785
rect 23756 35819 23808 35828
rect 23756 35785 23765 35819
rect 23765 35785 23799 35819
rect 23799 35785 23808 35819
rect 23756 35776 23808 35785
rect 25412 35776 25464 35828
rect 25780 35776 25832 35828
rect 26056 35776 26108 35828
rect 26516 35776 26568 35828
rect 26700 35776 26752 35828
rect 14832 35640 14884 35692
rect 18328 35640 18380 35692
rect 11428 35572 11480 35624
rect 13268 35615 13320 35624
rect 13268 35581 13277 35615
rect 13277 35581 13311 35615
rect 13311 35581 13320 35615
rect 13268 35572 13320 35581
rect 16948 35615 17000 35624
rect 16948 35581 16957 35615
rect 16957 35581 16991 35615
rect 16991 35581 17000 35615
rect 16948 35572 17000 35581
rect 11612 35504 11664 35556
rect 12808 35504 12860 35556
rect 13820 35504 13872 35556
rect 14188 35504 14240 35556
rect 16580 35504 16632 35556
rect 17684 35572 17736 35624
rect 19340 35640 19392 35692
rect 20536 35708 20588 35760
rect 23572 35708 23624 35760
rect 24492 35708 24544 35760
rect 20168 35683 20220 35692
rect 20168 35649 20177 35683
rect 20177 35649 20211 35683
rect 20211 35649 20220 35683
rect 20168 35640 20220 35649
rect 21456 35640 21508 35692
rect 24308 35683 24360 35692
rect 23480 35572 23532 35624
rect 24308 35649 24317 35683
rect 24317 35649 24351 35683
rect 24351 35649 24360 35683
rect 24308 35640 24360 35649
rect 24400 35640 24452 35692
rect 24676 35572 24728 35624
rect 25136 35683 25188 35692
rect 25136 35649 25145 35683
rect 25145 35649 25179 35683
rect 25179 35649 25188 35683
rect 25136 35640 25188 35649
rect 25596 35640 25648 35692
rect 27344 35640 27396 35692
rect 28264 35683 28316 35692
rect 28264 35649 28273 35683
rect 28273 35649 28307 35683
rect 28307 35649 28316 35683
rect 28264 35640 28316 35649
rect 25320 35572 25372 35624
rect 17868 35504 17920 35556
rect 6460 35436 6512 35488
rect 7196 35479 7248 35488
rect 7196 35445 7205 35479
rect 7205 35445 7239 35479
rect 7239 35445 7248 35479
rect 7196 35436 7248 35445
rect 9588 35436 9640 35488
rect 9864 35436 9916 35488
rect 9956 35479 10008 35488
rect 9956 35445 9965 35479
rect 9965 35445 9999 35479
rect 9999 35445 10008 35479
rect 9956 35436 10008 35445
rect 10508 35479 10560 35488
rect 10508 35445 10517 35479
rect 10517 35445 10551 35479
rect 10551 35445 10560 35479
rect 10508 35436 10560 35445
rect 12348 35436 12400 35488
rect 12992 35436 13044 35488
rect 16120 35479 16172 35488
rect 16120 35445 16129 35479
rect 16129 35445 16163 35479
rect 16163 35445 16172 35479
rect 16120 35436 16172 35445
rect 18144 35436 18196 35488
rect 25136 35504 25188 35556
rect 19156 35436 19208 35488
rect 24860 35479 24912 35488
rect 24860 35445 24869 35479
rect 24869 35445 24903 35479
rect 24903 35445 24912 35479
rect 24860 35436 24912 35445
rect 25228 35436 25280 35488
rect 26792 35572 26844 35624
rect 26148 35504 26200 35556
rect 27160 35572 27212 35624
rect 28172 35572 28224 35624
rect 29184 35776 29236 35828
rect 29276 35819 29328 35828
rect 29276 35785 29285 35819
rect 29285 35785 29319 35819
rect 29319 35785 29328 35819
rect 29276 35776 29328 35785
rect 29736 35776 29788 35828
rect 33048 35819 33100 35828
rect 33048 35785 33057 35819
rect 33057 35785 33091 35819
rect 33091 35785 33100 35819
rect 33048 35776 33100 35785
rect 29092 35751 29144 35760
rect 29092 35717 29101 35751
rect 29101 35717 29135 35751
rect 29135 35717 29144 35751
rect 29092 35708 29144 35717
rect 29000 35640 29052 35692
rect 30380 35640 30432 35692
rect 31024 35708 31076 35760
rect 32220 35640 32272 35692
rect 29736 35572 29788 35624
rect 30288 35572 30340 35624
rect 28908 35504 28960 35556
rect 25964 35436 26016 35488
rect 26240 35479 26292 35488
rect 26240 35445 26249 35479
rect 26249 35445 26283 35479
rect 26283 35445 26292 35479
rect 26240 35436 26292 35445
rect 28172 35479 28224 35488
rect 28172 35445 28181 35479
rect 28181 35445 28215 35479
rect 28215 35445 28224 35479
rect 28172 35436 28224 35445
rect 28816 35479 28868 35488
rect 28816 35445 28825 35479
rect 28825 35445 28859 35479
rect 28859 35445 28868 35479
rect 28816 35436 28868 35445
rect 29092 35436 29144 35488
rect 30104 35436 30156 35488
rect 31760 35436 31812 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5632 35275 5684 35284
rect 5632 35241 5641 35275
rect 5641 35241 5675 35275
rect 5675 35241 5684 35275
rect 5632 35232 5684 35241
rect 6092 35232 6144 35284
rect 7380 35232 7432 35284
rect 8668 35232 8720 35284
rect 9864 35232 9916 35284
rect 11152 35232 11204 35284
rect 11704 35232 11756 35284
rect 12716 35275 12768 35284
rect 12716 35241 12725 35275
rect 12725 35241 12759 35275
rect 12759 35241 12768 35275
rect 12716 35232 12768 35241
rect 12808 35232 12860 35284
rect 12992 35232 13044 35284
rect 7656 35207 7708 35216
rect 7656 35173 7665 35207
rect 7665 35173 7699 35207
rect 7699 35173 7708 35207
rect 7656 35164 7708 35173
rect 9036 35164 9088 35216
rect 940 35028 992 35080
rect 7012 35028 7064 35080
rect 7564 35071 7616 35080
rect 7564 35037 7573 35071
rect 7573 35037 7607 35071
rect 7607 35037 7616 35071
rect 7564 35028 7616 35037
rect 8576 35139 8628 35148
rect 8576 35105 8585 35139
rect 8585 35105 8619 35139
rect 8619 35105 8628 35139
rect 8576 35096 8628 35105
rect 8944 35139 8996 35148
rect 8944 35105 8953 35139
rect 8953 35105 8987 35139
rect 8987 35105 8996 35139
rect 8944 35096 8996 35105
rect 4988 34960 5040 35012
rect 6552 34960 6604 35012
rect 6828 34960 6880 35012
rect 11336 35164 11388 35216
rect 12624 35207 12676 35216
rect 12624 35173 12633 35207
rect 12633 35173 12667 35207
rect 12667 35173 12676 35207
rect 12624 35164 12676 35173
rect 9772 35139 9824 35148
rect 9772 35105 9781 35139
rect 9781 35105 9815 35139
rect 9815 35105 9824 35139
rect 9772 35096 9824 35105
rect 9220 35028 9272 35080
rect 10324 35071 10376 35080
rect 10324 35037 10333 35071
rect 10333 35037 10367 35071
rect 10367 35037 10376 35071
rect 10324 35028 10376 35037
rect 10508 35071 10560 35080
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 10876 35028 10928 35080
rect 11428 35096 11480 35148
rect 11796 35071 11848 35080
rect 11796 35037 11805 35071
rect 11805 35037 11839 35071
rect 11839 35037 11848 35071
rect 11796 35028 11848 35037
rect 13360 35164 13412 35216
rect 13452 35096 13504 35148
rect 3332 34892 3384 34944
rect 4620 34892 4672 34944
rect 8208 34892 8260 34944
rect 9864 34892 9916 34944
rect 11244 34960 11296 35012
rect 13176 35071 13228 35080
rect 13176 35037 13185 35071
rect 13185 35037 13219 35071
rect 13219 35037 13228 35071
rect 13176 35028 13228 35037
rect 14372 35232 14424 35284
rect 15384 35232 15436 35284
rect 15568 35164 15620 35216
rect 16764 35164 16816 35216
rect 15752 35096 15804 35148
rect 17040 35164 17092 35216
rect 17224 35164 17276 35216
rect 18328 35232 18380 35284
rect 24492 35232 24544 35284
rect 24676 35232 24728 35284
rect 25228 35275 25280 35284
rect 25228 35241 25237 35275
rect 25237 35241 25271 35275
rect 25271 35241 25280 35275
rect 25228 35232 25280 35241
rect 17132 35139 17184 35148
rect 17132 35105 17141 35139
rect 17141 35105 17175 35139
rect 17175 35105 17184 35139
rect 17132 35096 17184 35105
rect 12256 35003 12308 35012
rect 12256 34969 12265 35003
rect 12265 34969 12299 35003
rect 12299 34969 12308 35003
rect 12256 34960 12308 34969
rect 10968 34935 11020 34944
rect 10968 34901 10977 34935
rect 10977 34901 11011 34935
rect 11011 34901 11020 34935
rect 10968 34892 11020 34901
rect 12808 34892 12860 34944
rect 13636 35071 13688 35080
rect 13636 35037 13645 35071
rect 13645 35037 13679 35071
rect 13679 35037 13688 35071
rect 13636 35028 13688 35037
rect 13912 35028 13964 35080
rect 14648 35028 14700 35080
rect 14924 34960 14976 35012
rect 14096 34892 14148 34944
rect 14188 34892 14240 34944
rect 16488 35028 16540 35080
rect 18696 35164 18748 35216
rect 19432 35164 19484 35216
rect 20076 35164 20128 35216
rect 20996 35164 21048 35216
rect 18512 35071 18564 35080
rect 18512 35037 18521 35071
rect 18521 35037 18555 35071
rect 18555 35037 18564 35071
rect 18512 35028 18564 35037
rect 20076 35071 20128 35080
rect 20076 35037 20085 35071
rect 20085 35037 20119 35071
rect 20119 35037 20128 35071
rect 20076 35028 20128 35037
rect 20904 34960 20956 35012
rect 16580 34892 16632 34944
rect 17132 34892 17184 34944
rect 18604 34892 18656 34944
rect 19064 34892 19116 34944
rect 20720 34935 20772 34944
rect 20720 34901 20729 34935
rect 20729 34901 20763 34935
rect 20763 34901 20772 34935
rect 20720 34892 20772 34901
rect 21088 35071 21140 35080
rect 21088 35037 21097 35071
rect 21097 35037 21131 35071
rect 21131 35037 21140 35071
rect 21088 35028 21140 35037
rect 22192 35096 22244 35148
rect 21364 35071 21416 35080
rect 21364 35037 21373 35071
rect 21373 35037 21407 35071
rect 21407 35037 21416 35071
rect 21364 35028 21416 35037
rect 24400 35164 24452 35216
rect 26700 35232 26752 35284
rect 27620 35232 27672 35284
rect 28632 35232 28684 35284
rect 30932 35232 30984 35284
rect 32220 35275 32272 35284
rect 32220 35241 32229 35275
rect 32229 35241 32263 35275
rect 32263 35241 32272 35275
rect 32220 35232 32272 35241
rect 23480 35096 23532 35148
rect 25872 35164 25924 35216
rect 27896 35207 27948 35216
rect 27896 35173 27905 35207
rect 27905 35173 27939 35207
rect 27939 35173 27948 35207
rect 27896 35164 27948 35173
rect 28264 35164 28316 35216
rect 30012 35164 30064 35216
rect 21824 35003 21876 35012
rect 21824 34969 21833 35003
rect 21833 34969 21867 35003
rect 21867 34969 21876 35003
rect 21824 34960 21876 34969
rect 22008 34960 22060 35012
rect 21088 34892 21140 34944
rect 22284 34935 22336 34944
rect 22284 34901 22293 34935
rect 22293 34901 22327 34935
rect 22327 34901 22336 34935
rect 22284 34892 22336 34901
rect 22652 34935 22704 34944
rect 22652 34901 22661 34935
rect 22661 34901 22695 34935
rect 22695 34901 22704 34935
rect 22652 34892 22704 34901
rect 24860 35096 24912 35148
rect 24952 35096 25004 35148
rect 25228 35028 25280 35080
rect 25504 35028 25556 35080
rect 25964 35028 26016 35080
rect 26884 35028 26936 35080
rect 28356 35096 28408 35148
rect 28908 35139 28960 35148
rect 28908 35105 28917 35139
rect 28917 35105 28951 35139
rect 28951 35105 28960 35139
rect 28908 35096 28960 35105
rect 25780 35003 25832 35012
rect 25780 34969 25789 35003
rect 25789 34969 25823 35003
rect 25823 34969 25832 35003
rect 25780 34960 25832 34969
rect 26056 34892 26108 34944
rect 26700 34892 26752 34944
rect 28080 35071 28132 35080
rect 28080 35037 28089 35071
rect 28089 35037 28123 35071
rect 28123 35037 28132 35071
rect 28080 35028 28132 35037
rect 28724 35028 28776 35080
rect 29828 35096 29880 35148
rect 28448 34935 28500 34944
rect 28448 34901 28457 34935
rect 28457 34901 28491 34935
rect 28491 34901 28500 34935
rect 28448 34892 28500 34901
rect 28540 34892 28592 34944
rect 30012 35003 30064 35012
rect 30012 34969 30021 35003
rect 30021 34969 30055 35003
rect 30055 34969 30064 35003
rect 30012 34960 30064 34969
rect 30196 35071 30248 35080
rect 30196 35037 30205 35071
rect 30205 35037 30239 35071
rect 30239 35037 30248 35071
rect 30196 35028 30248 35037
rect 32680 35164 32732 35216
rect 31024 35139 31076 35148
rect 31024 35105 31033 35139
rect 31033 35105 31067 35139
rect 31067 35105 31076 35139
rect 31024 35096 31076 35105
rect 31760 35139 31812 35148
rect 31760 35105 31769 35139
rect 31769 35105 31803 35139
rect 31803 35105 31812 35139
rect 31760 35096 31812 35105
rect 30840 35028 30892 35080
rect 30656 34960 30708 35012
rect 32312 35028 32364 35080
rect 32128 34960 32180 35012
rect 29920 34935 29972 34944
rect 29920 34901 29929 34935
rect 29929 34901 29963 34935
rect 29963 34901 29972 34935
rect 29920 34892 29972 34901
rect 31392 34892 31444 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4712 34688 4764 34740
rect 7748 34731 7800 34740
rect 7748 34697 7757 34731
rect 7757 34697 7791 34731
rect 7791 34697 7800 34731
rect 7748 34688 7800 34697
rect 4988 34552 5040 34604
rect 6920 34552 6972 34604
rect 7012 34552 7064 34604
rect 1768 34527 1820 34536
rect 1768 34493 1777 34527
rect 1777 34493 1811 34527
rect 1811 34493 1820 34527
rect 1768 34484 1820 34493
rect 2136 34527 2188 34536
rect 2136 34493 2145 34527
rect 2145 34493 2179 34527
rect 2179 34493 2188 34527
rect 2136 34484 2188 34493
rect 2228 34484 2280 34536
rect 2872 34527 2924 34536
rect 2872 34493 2881 34527
rect 2881 34493 2915 34527
rect 2915 34493 2924 34527
rect 2872 34484 2924 34493
rect 3516 34527 3568 34536
rect 3516 34493 3525 34527
rect 3525 34493 3559 34527
rect 3559 34493 3568 34527
rect 3516 34484 3568 34493
rect 9404 34620 9456 34672
rect 9588 34663 9640 34672
rect 9588 34629 9597 34663
rect 9597 34629 9631 34663
rect 9631 34629 9640 34663
rect 9588 34620 9640 34629
rect 8668 34484 8720 34536
rect 9220 34527 9272 34536
rect 9220 34493 9229 34527
rect 9229 34493 9263 34527
rect 9263 34493 9272 34527
rect 9220 34484 9272 34493
rect 9588 34484 9640 34536
rect 9956 34688 10008 34740
rect 10140 34688 10192 34740
rect 11428 34688 11480 34740
rect 11980 34688 12032 34740
rect 9864 34595 9916 34604
rect 9864 34561 9873 34595
rect 9873 34561 9907 34595
rect 9907 34561 9916 34595
rect 9864 34552 9916 34561
rect 9956 34595 10008 34604
rect 9956 34561 9965 34595
rect 9965 34561 9999 34595
rect 9999 34561 10008 34595
rect 9956 34552 10008 34561
rect 10140 34552 10192 34604
rect 13084 34688 13136 34740
rect 13912 34688 13964 34740
rect 14096 34688 14148 34740
rect 14924 34731 14976 34740
rect 14924 34697 14933 34731
rect 14933 34697 14967 34731
rect 14967 34697 14976 34731
rect 14924 34688 14976 34697
rect 15108 34688 15160 34740
rect 15476 34688 15528 34740
rect 16212 34688 16264 34740
rect 16396 34731 16448 34740
rect 16396 34697 16405 34731
rect 16405 34697 16439 34731
rect 16439 34697 16448 34731
rect 16396 34688 16448 34697
rect 11796 34484 11848 34536
rect 12164 34595 12216 34604
rect 12164 34561 12173 34595
rect 12173 34561 12207 34595
rect 12207 34561 12216 34595
rect 12164 34552 12216 34561
rect 12808 34552 12860 34604
rect 14188 34663 14240 34672
rect 14188 34629 14197 34663
rect 14197 34629 14231 34663
rect 14231 34629 14240 34663
rect 14188 34620 14240 34629
rect 14464 34620 14516 34672
rect 13084 34484 13136 34536
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 14096 34552 14148 34604
rect 16948 34688 17000 34740
rect 17500 34688 17552 34740
rect 20076 34688 20128 34740
rect 20720 34688 20772 34740
rect 20904 34688 20956 34740
rect 21824 34688 21876 34740
rect 22192 34731 22244 34740
rect 22192 34697 22201 34731
rect 22201 34697 22235 34731
rect 22235 34697 22244 34731
rect 22192 34688 22244 34697
rect 22652 34688 22704 34740
rect 23020 34688 23072 34740
rect 26700 34688 26752 34740
rect 14280 34527 14332 34536
rect 14280 34493 14289 34527
rect 14289 34493 14323 34527
rect 14323 34493 14332 34527
rect 14280 34484 14332 34493
rect 14556 34484 14608 34536
rect 15844 34552 15896 34604
rect 16672 34620 16724 34672
rect 16764 34620 16816 34672
rect 16488 34595 16540 34604
rect 16488 34561 16497 34595
rect 16497 34561 16531 34595
rect 16531 34561 16540 34595
rect 16488 34552 16540 34561
rect 19432 34620 19484 34672
rect 19064 34552 19116 34604
rect 15292 34484 15344 34536
rect 16580 34484 16632 34536
rect 18696 34484 18748 34536
rect 19156 34527 19208 34536
rect 19156 34493 19165 34527
rect 19165 34493 19199 34527
rect 19199 34493 19208 34527
rect 19156 34484 19208 34493
rect 19892 34552 19944 34604
rect 20628 34552 20680 34604
rect 6184 34459 6236 34468
rect 6184 34425 6193 34459
rect 6193 34425 6227 34459
rect 6227 34425 6236 34459
rect 6184 34416 6236 34425
rect 10324 34416 10376 34468
rect 3424 34391 3476 34400
rect 3424 34357 3433 34391
rect 3433 34357 3467 34391
rect 3467 34357 3476 34391
rect 3424 34348 3476 34357
rect 5356 34348 5408 34400
rect 6000 34348 6052 34400
rect 6552 34348 6604 34400
rect 7104 34348 7156 34400
rect 10876 34348 10928 34400
rect 10968 34391 11020 34400
rect 10968 34357 10977 34391
rect 10977 34357 11011 34391
rect 11011 34357 11020 34391
rect 10968 34348 11020 34357
rect 12808 34416 12860 34468
rect 12440 34391 12492 34400
rect 12440 34357 12449 34391
rect 12449 34357 12483 34391
rect 12483 34357 12492 34391
rect 12440 34348 12492 34357
rect 12992 34391 13044 34400
rect 12992 34357 13001 34391
rect 13001 34357 13035 34391
rect 13035 34357 13044 34391
rect 12992 34348 13044 34357
rect 15108 34416 15160 34468
rect 15476 34416 15528 34468
rect 17040 34348 17092 34400
rect 19708 34527 19760 34536
rect 19708 34493 19717 34527
rect 19717 34493 19751 34527
rect 19751 34493 19760 34527
rect 19708 34484 19760 34493
rect 21272 34552 21324 34604
rect 20720 34348 20772 34400
rect 20996 34348 21048 34400
rect 21272 34348 21324 34400
rect 21824 34595 21876 34604
rect 21824 34561 21833 34595
rect 21833 34561 21867 34595
rect 21867 34561 21876 34595
rect 21824 34552 21876 34561
rect 22284 34552 22336 34604
rect 22376 34527 22428 34536
rect 22376 34493 22385 34527
rect 22385 34493 22419 34527
rect 22419 34493 22428 34527
rect 22376 34484 22428 34493
rect 23296 34527 23348 34536
rect 23296 34493 23305 34527
rect 23305 34493 23339 34527
rect 23339 34493 23348 34527
rect 23296 34484 23348 34493
rect 23756 34620 23808 34672
rect 24676 34620 24728 34672
rect 24768 34663 24820 34672
rect 24768 34629 24777 34663
rect 24777 34629 24811 34663
rect 24811 34629 24820 34663
rect 24768 34620 24820 34629
rect 24492 34552 24544 34604
rect 25412 34595 25464 34604
rect 25412 34561 25421 34595
rect 25421 34561 25455 34595
rect 25455 34561 25464 34595
rect 25412 34552 25464 34561
rect 25688 34620 25740 34672
rect 26424 34620 26476 34672
rect 25872 34552 25924 34604
rect 26056 34552 26108 34604
rect 27712 34688 27764 34740
rect 28172 34688 28224 34740
rect 28356 34731 28408 34740
rect 28356 34697 28365 34731
rect 28365 34697 28399 34731
rect 28399 34697 28408 34731
rect 28356 34688 28408 34697
rect 28448 34688 28500 34740
rect 29552 34688 29604 34740
rect 29920 34688 29972 34740
rect 30288 34688 30340 34740
rect 32312 34731 32364 34740
rect 32312 34697 32321 34731
rect 32321 34697 32355 34731
rect 32355 34697 32364 34731
rect 32312 34688 32364 34697
rect 26976 34595 27028 34604
rect 26976 34561 26985 34595
rect 26985 34561 27019 34595
rect 27019 34561 27028 34595
rect 26976 34552 27028 34561
rect 27528 34552 27580 34604
rect 24860 34484 24912 34536
rect 25044 34484 25096 34536
rect 26148 34484 26200 34536
rect 26884 34484 26936 34536
rect 24400 34416 24452 34468
rect 23020 34391 23072 34400
rect 23020 34357 23029 34391
rect 23029 34357 23063 34391
rect 23063 34357 23072 34391
rect 23020 34348 23072 34357
rect 23848 34348 23900 34400
rect 25136 34391 25188 34400
rect 25136 34357 25145 34391
rect 25145 34357 25179 34391
rect 25179 34357 25188 34391
rect 25136 34348 25188 34357
rect 26424 34459 26476 34468
rect 26424 34425 26433 34459
rect 26433 34425 26467 34459
rect 26467 34425 26476 34459
rect 26424 34416 26476 34425
rect 26516 34459 26568 34468
rect 26516 34425 26525 34459
rect 26525 34425 26559 34459
rect 26559 34425 26568 34459
rect 26516 34416 26568 34425
rect 28080 34484 28132 34536
rect 28908 34484 28960 34536
rect 29368 34527 29420 34536
rect 29368 34493 29377 34527
rect 29377 34493 29411 34527
rect 29411 34493 29420 34527
rect 29368 34484 29420 34493
rect 25596 34348 25648 34400
rect 27160 34348 27212 34400
rect 27344 34348 27396 34400
rect 28540 34348 28592 34400
rect 30564 34348 30616 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2136 34144 2188 34196
rect 4620 34144 4672 34196
rect 6828 34144 6880 34196
rect 7564 34144 7616 34196
rect 8576 34144 8628 34196
rect 9128 34144 9180 34196
rect 9312 34144 9364 34196
rect 9772 34144 9824 34196
rect 9956 34144 10008 34196
rect 10968 34144 11020 34196
rect 11244 34144 11296 34196
rect 12256 34144 12308 34196
rect 13544 34144 13596 34196
rect 15200 34144 15252 34196
rect 4988 34119 5040 34128
rect 4988 34085 4997 34119
rect 4997 34085 5031 34119
rect 5031 34085 5040 34119
rect 4988 34076 5040 34085
rect 1952 34008 2004 34060
rect 3332 34051 3384 34060
rect 3332 34017 3341 34051
rect 3341 34017 3375 34051
rect 3375 34017 3384 34051
rect 3332 34008 3384 34017
rect 4068 34008 4120 34060
rect 5540 34076 5592 34128
rect 6276 34008 6328 34060
rect 6460 34051 6512 34060
rect 6460 34017 6469 34051
rect 6469 34017 6503 34051
rect 6503 34017 6512 34051
rect 6460 34008 6512 34017
rect 6644 34051 6696 34060
rect 6644 34017 6653 34051
rect 6653 34017 6687 34051
rect 6687 34017 6696 34051
rect 6644 34008 6696 34017
rect 940 33940 992 33992
rect 2044 33983 2096 33992
rect 2044 33949 2053 33983
rect 2053 33949 2087 33983
rect 2087 33949 2096 33983
rect 2044 33940 2096 33949
rect 3424 33872 3476 33924
rect 7196 33940 7248 33992
rect 7472 33940 7524 33992
rect 12624 34076 12676 34128
rect 8668 34008 8720 34060
rect 8760 33940 8812 33992
rect 10876 34051 10928 34060
rect 10876 34017 10885 34051
rect 10885 34017 10919 34051
rect 10919 34017 10928 34051
rect 10876 34008 10928 34017
rect 7012 33872 7064 33924
rect 9588 33872 9640 33924
rect 10508 33915 10560 33924
rect 10508 33881 10517 33915
rect 10517 33881 10551 33915
rect 10551 33881 10560 33915
rect 10508 33872 10560 33881
rect 2596 33847 2648 33856
rect 2596 33813 2605 33847
rect 2605 33813 2639 33847
rect 2639 33813 2648 33847
rect 2596 33804 2648 33813
rect 3608 33804 3660 33856
rect 3884 33804 3936 33856
rect 5448 33847 5500 33856
rect 5448 33813 5457 33847
rect 5457 33813 5491 33847
rect 5491 33813 5500 33847
rect 5448 33804 5500 33813
rect 7288 33804 7340 33856
rect 11060 33983 11112 33992
rect 11060 33949 11069 33983
rect 11069 33949 11103 33983
rect 11103 33949 11112 33983
rect 11060 33940 11112 33949
rect 11244 33804 11296 33856
rect 11704 34051 11756 34060
rect 11704 34017 11713 34051
rect 11713 34017 11747 34051
rect 11747 34017 11756 34051
rect 11704 34008 11756 34017
rect 12072 33983 12124 33992
rect 12072 33949 12081 33983
rect 12081 33949 12115 33983
rect 12115 33949 12124 33983
rect 12072 33940 12124 33949
rect 12164 33983 12216 33992
rect 12164 33949 12173 33983
rect 12173 33949 12207 33983
rect 12207 33949 12216 33983
rect 12164 33940 12216 33949
rect 12440 33983 12492 33992
rect 12440 33949 12449 33983
rect 12449 33949 12483 33983
rect 12483 33949 12492 33983
rect 12440 33940 12492 33949
rect 12808 33940 12860 33992
rect 15108 34076 15160 34128
rect 13268 34051 13320 34060
rect 13268 34017 13277 34051
rect 13277 34017 13311 34051
rect 13311 34017 13320 34051
rect 13268 34008 13320 34017
rect 13912 34008 13964 34060
rect 13084 33983 13136 33992
rect 13084 33949 13093 33983
rect 13093 33949 13127 33983
rect 13127 33949 13136 33983
rect 13084 33940 13136 33949
rect 12716 33872 12768 33924
rect 13544 33940 13596 33992
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 14832 34008 14884 34060
rect 17408 34144 17460 34196
rect 19616 34144 19668 34196
rect 22376 34144 22428 34196
rect 23204 34144 23256 34196
rect 24584 34144 24636 34196
rect 24865 34144 24917 34196
rect 26424 34144 26476 34196
rect 26516 34144 26568 34196
rect 27068 34144 27120 34196
rect 29184 34144 29236 34196
rect 31392 34187 31444 34196
rect 31392 34153 31401 34187
rect 31401 34153 31435 34187
rect 31435 34153 31444 34187
rect 31392 34144 31444 34153
rect 14556 33983 14608 33992
rect 14556 33949 14565 33983
rect 14565 33949 14599 33983
rect 14599 33949 14608 33983
rect 14556 33940 14608 33949
rect 15016 33940 15068 33992
rect 15108 33940 15160 33992
rect 15384 33940 15436 33992
rect 16028 34076 16080 34128
rect 17132 34119 17184 34128
rect 17132 34085 17141 34119
rect 17141 34085 17175 34119
rect 17175 34085 17184 34119
rect 17132 34076 17184 34085
rect 15844 34051 15896 34060
rect 15844 34017 15853 34051
rect 15853 34017 15887 34051
rect 15887 34017 15896 34051
rect 15844 34008 15896 34017
rect 15936 33983 15988 33992
rect 15936 33949 15945 33983
rect 15945 33949 15979 33983
rect 15979 33949 15988 33983
rect 15936 33940 15988 33949
rect 14740 33872 14792 33924
rect 16396 33872 16448 33924
rect 17040 33872 17092 33924
rect 17592 33983 17644 33992
rect 17592 33949 17601 33983
rect 17601 33949 17635 33983
rect 17635 33949 17644 33983
rect 17592 33940 17644 33949
rect 17776 33983 17828 33992
rect 17776 33949 17785 33983
rect 17785 33949 17819 33983
rect 17819 33949 17828 33983
rect 17776 33940 17828 33949
rect 17960 33872 18012 33924
rect 18604 34051 18656 34060
rect 18604 34017 18613 34051
rect 18613 34017 18647 34051
rect 18647 34017 18656 34051
rect 18604 34008 18656 34017
rect 20352 34076 20404 34128
rect 22652 34076 22704 34128
rect 25044 34076 25096 34128
rect 26240 34076 26292 34128
rect 27620 34076 27672 34128
rect 27712 34076 27764 34128
rect 18788 33940 18840 33992
rect 22192 34008 22244 34060
rect 18972 33983 19024 33992
rect 18972 33949 18981 33983
rect 18981 33949 19015 33983
rect 19015 33949 19024 33983
rect 18972 33940 19024 33949
rect 19616 33983 19668 33992
rect 19616 33949 19625 33983
rect 19625 33949 19659 33983
rect 19659 33949 19668 33983
rect 19616 33940 19668 33949
rect 19892 33940 19944 33992
rect 20352 33940 20404 33992
rect 21364 33940 21416 33992
rect 21640 33940 21692 33992
rect 22744 33940 22796 33992
rect 26516 34008 26568 34060
rect 23848 33940 23900 33992
rect 21916 33872 21968 33924
rect 13820 33804 13872 33856
rect 17408 33804 17460 33856
rect 18788 33804 18840 33856
rect 19708 33804 19760 33856
rect 21364 33847 21416 33856
rect 21364 33813 21373 33847
rect 21373 33813 21407 33847
rect 21407 33813 21416 33847
rect 21364 33804 21416 33813
rect 22928 33872 22980 33924
rect 24032 33872 24084 33924
rect 22652 33804 22704 33856
rect 22744 33804 22796 33856
rect 23388 33804 23440 33856
rect 24308 33872 24360 33924
rect 24676 33804 24728 33856
rect 24952 33804 25004 33856
rect 25044 33804 25096 33856
rect 25504 33940 25556 33992
rect 25872 33940 25924 33992
rect 26148 33983 26200 33992
rect 26148 33949 26157 33983
rect 26157 33949 26191 33983
rect 26191 33949 26200 33983
rect 26148 33940 26200 33949
rect 25688 33872 25740 33924
rect 25964 33847 26016 33856
rect 25964 33813 25973 33847
rect 25973 33813 26007 33847
rect 26007 33813 26016 33847
rect 25964 33804 26016 33813
rect 26056 33804 26108 33856
rect 26700 33940 26752 33992
rect 27068 33983 27120 33992
rect 27068 33949 27077 33983
rect 27077 33949 27111 33983
rect 27111 33949 27120 33983
rect 27068 33940 27120 33949
rect 27160 33983 27212 33992
rect 27160 33949 27169 33983
rect 27169 33949 27203 33983
rect 27203 33949 27212 33983
rect 27160 33940 27212 33949
rect 27988 34051 28040 34060
rect 27988 34017 27997 34051
rect 27997 34017 28031 34051
rect 28031 34017 28040 34051
rect 27988 34008 28040 34017
rect 28356 34008 28408 34060
rect 28816 34008 28868 34060
rect 27528 33940 27580 33992
rect 27436 33915 27488 33924
rect 27436 33881 27445 33915
rect 27445 33881 27479 33915
rect 27479 33881 27488 33915
rect 27436 33872 27488 33881
rect 27896 33940 27948 33992
rect 28080 33983 28132 33992
rect 28080 33949 28089 33983
rect 28089 33949 28123 33983
rect 28123 33949 28132 33983
rect 28080 33940 28132 33949
rect 28264 33940 28316 33992
rect 28908 33983 28960 33992
rect 28908 33949 28917 33983
rect 28917 33949 28951 33983
rect 28951 33949 28960 33983
rect 28908 33940 28960 33949
rect 30564 34008 30616 34060
rect 30656 34051 30708 34060
rect 30656 34017 30665 34051
rect 30665 34017 30699 34051
rect 30699 34017 30708 34051
rect 30656 34008 30708 34017
rect 29460 33940 29512 33992
rect 27160 33804 27212 33856
rect 27620 33847 27672 33856
rect 27620 33813 27629 33847
rect 27629 33813 27663 33847
rect 27663 33813 27672 33847
rect 27620 33804 27672 33813
rect 27712 33847 27764 33856
rect 27712 33813 27721 33847
rect 27721 33813 27755 33847
rect 27755 33813 27764 33847
rect 27712 33804 27764 33813
rect 28080 33804 28132 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1952 33643 2004 33652
rect 1952 33609 1961 33643
rect 1961 33609 1995 33643
rect 1995 33609 2004 33643
rect 1952 33600 2004 33609
rect 2044 33600 2096 33652
rect 2596 33600 2648 33652
rect 3516 33600 3568 33652
rect 5448 33600 5500 33652
rect 8668 33643 8720 33652
rect 8668 33609 8677 33643
rect 8677 33609 8711 33643
rect 8711 33609 8720 33643
rect 8668 33600 8720 33609
rect 8760 33643 8812 33652
rect 8760 33609 8769 33643
rect 8769 33609 8803 33643
rect 8803 33609 8812 33643
rect 8760 33600 8812 33609
rect 9588 33600 9640 33652
rect 11060 33600 11112 33652
rect 1860 33396 1912 33448
rect 4712 33464 4764 33516
rect 6000 33464 6052 33516
rect 6644 33464 6696 33516
rect 11520 33600 11572 33652
rect 12164 33600 12216 33652
rect 12532 33600 12584 33652
rect 13084 33643 13136 33652
rect 13084 33609 13093 33643
rect 13093 33609 13127 33643
rect 13127 33609 13136 33643
rect 13084 33600 13136 33609
rect 13176 33600 13228 33652
rect 3976 33439 4028 33448
rect 3976 33405 3985 33439
rect 3985 33405 4019 33439
rect 4019 33405 4028 33439
rect 3976 33396 4028 33405
rect 4068 33439 4120 33448
rect 4068 33405 4077 33439
rect 4077 33405 4111 33439
rect 4111 33405 4120 33439
rect 4068 33396 4120 33405
rect 4896 33439 4948 33448
rect 4896 33405 4905 33439
rect 4905 33405 4939 33439
rect 4939 33405 4948 33439
rect 4896 33396 4948 33405
rect 3884 33328 3936 33380
rect 7380 33439 7432 33448
rect 7380 33405 7389 33439
rect 7389 33405 7423 33439
rect 7423 33405 7432 33439
rect 7380 33396 7432 33405
rect 9128 33464 9180 33516
rect 9220 33507 9272 33516
rect 9220 33473 9229 33507
rect 9229 33473 9263 33507
rect 9263 33473 9272 33507
rect 9220 33464 9272 33473
rect 9312 33464 9364 33516
rect 10600 33507 10652 33516
rect 10600 33473 10609 33507
rect 10609 33473 10643 33507
rect 10643 33473 10652 33507
rect 10600 33464 10652 33473
rect 10692 33507 10744 33516
rect 10692 33473 10701 33507
rect 10701 33473 10735 33507
rect 10735 33473 10744 33507
rect 10692 33464 10744 33473
rect 11060 33396 11112 33448
rect 11244 33464 11296 33516
rect 11704 33507 11756 33516
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 10968 33328 11020 33380
rect 3424 33260 3476 33312
rect 5356 33260 5408 33312
rect 5632 33260 5684 33312
rect 7932 33303 7984 33312
rect 7932 33269 7941 33303
rect 7941 33269 7975 33303
rect 7975 33269 7984 33303
rect 7932 33260 7984 33269
rect 8392 33303 8444 33312
rect 8392 33269 8401 33303
rect 8401 33269 8435 33303
rect 8435 33269 8444 33303
rect 8392 33260 8444 33269
rect 10876 33260 10928 33312
rect 11336 33396 11388 33448
rect 12164 33464 12216 33516
rect 12256 33507 12308 33516
rect 12256 33473 12265 33507
rect 12265 33473 12299 33507
rect 12299 33473 12308 33507
rect 12256 33464 12308 33473
rect 12348 33507 12400 33516
rect 12348 33473 12357 33507
rect 12357 33473 12391 33507
rect 12391 33473 12400 33507
rect 12348 33464 12400 33473
rect 12716 33464 12768 33516
rect 12900 33507 12952 33516
rect 12900 33473 12909 33507
rect 12909 33473 12943 33507
rect 12943 33473 12952 33507
rect 14004 33643 14056 33652
rect 14004 33609 14013 33643
rect 14013 33609 14047 33643
rect 14047 33609 14056 33643
rect 14004 33600 14056 33609
rect 15936 33600 15988 33652
rect 16212 33600 16264 33652
rect 16304 33600 16356 33652
rect 16764 33600 16816 33652
rect 18052 33600 18104 33652
rect 18144 33600 18196 33652
rect 18972 33600 19024 33652
rect 20812 33600 20864 33652
rect 14464 33532 14516 33584
rect 12900 33464 12952 33473
rect 13636 33464 13688 33516
rect 15108 33532 15160 33584
rect 15292 33532 15344 33584
rect 12532 33328 12584 33380
rect 12808 33328 12860 33380
rect 12164 33260 12216 33312
rect 14188 33396 14240 33448
rect 14648 33464 14700 33516
rect 15200 33464 15252 33516
rect 15660 33464 15712 33516
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 17500 33575 17552 33584
rect 17500 33541 17509 33575
rect 17509 33541 17543 33575
rect 17543 33541 17552 33575
rect 17500 33532 17552 33541
rect 21364 33600 21416 33652
rect 16580 33464 16632 33516
rect 17224 33507 17276 33516
rect 17224 33473 17233 33507
rect 17233 33473 17267 33507
rect 17267 33473 17276 33507
rect 17224 33464 17276 33473
rect 17868 33464 17920 33516
rect 14924 33396 14976 33448
rect 16212 33396 16264 33448
rect 17960 33396 18012 33448
rect 18512 33439 18564 33448
rect 18512 33405 18521 33439
rect 18521 33405 18555 33439
rect 18555 33405 18564 33439
rect 18512 33396 18564 33405
rect 19064 33507 19116 33516
rect 19064 33473 19073 33507
rect 19073 33473 19107 33507
rect 19107 33473 19116 33507
rect 19064 33464 19116 33473
rect 19156 33464 19208 33516
rect 19432 33464 19484 33516
rect 20444 33464 20496 33516
rect 21088 33464 21140 33516
rect 22376 33600 22428 33652
rect 24400 33643 24452 33652
rect 24400 33609 24409 33643
rect 24409 33609 24443 33643
rect 24443 33609 24452 33643
rect 24400 33600 24452 33609
rect 22008 33532 22060 33584
rect 23020 33532 23072 33584
rect 24216 33532 24268 33584
rect 27712 33600 27764 33652
rect 28080 33600 28132 33652
rect 24860 33532 24912 33584
rect 26792 33532 26844 33584
rect 27252 33532 27304 33584
rect 21548 33507 21600 33516
rect 21548 33473 21557 33507
rect 21557 33473 21591 33507
rect 21591 33473 21600 33507
rect 21548 33464 21600 33473
rect 23204 33464 23256 33516
rect 23664 33507 23716 33516
rect 23664 33473 23673 33507
rect 23673 33473 23707 33507
rect 23707 33473 23716 33507
rect 23664 33464 23716 33473
rect 20904 33396 20956 33448
rect 21916 33396 21968 33448
rect 24584 33507 24636 33516
rect 24584 33473 24593 33507
rect 24593 33473 24627 33507
rect 24627 33473 24636 33507
rect 24584 33464 24636 33473
rect 25228 33464 25280 33516
rect 25412 33464 25464 33516
rect 25596 33464 25648 33516
rect 24860 33396 24912 33448
rect 25688 33396 25740 33448
rect 25872 33439 25924 33448
rect 25872 33405 25881 33439
rect 25881 33405 25915 33439
rect 25915 33405 25924 33439
rect 25872 33396 25924 33405
rect 26240 33507 26292 33516
rect 26240 33473 26249 33507
rect 26249 33473 26283 33507
rect 26283 33473 26292 33507
rect 26240 33464 26292 33473
rect 26516 33396 26568 33448
rect 28908 33575 28960 33584
rect 28908 33541 28917 33575
rect 28917 33541 28951 33575
rect 28951 33541 28960 33575
rect 28908 33532 28960 33541
rect 29736 33532 29788 33584
rect 27804 33464 27856 33516
rect 28172 33507 28224 33516
rect 28172 33473 28181 33507
rect 28181 33473 28215 33507
rect 28215 33473 28224 33507
rect 28172 33464 28224 33473
rect 14740 33328 14792 33380
rect 13360 33303 13412 33312
rect 13360 33269 13369 33303
rect 13369 33269 13403 33303
rect 13403 33269 13412 33303
rect 13360 33260 13412 33269
rect 13728 33260 13780 33312
rect 14648 33260 14700 33312
rect 15568 33260 15620 33312
rect 26240 33328 26292 33380
rect 26332 33328 26384 33380
rect 27344 33328 27396 33380
rect 28540 33396 28592 33448
rect 29000 33464 29052 33516
rect 16856 33260 16908 33312
rect 18880 33260 18932 33312
rect 19984 33260 20036 33312
rect 20536 33260 20588 33312
rect 22376 33260 22428 33312
rect 23572 33303 23624 33312
rect 23572 33269 23581 33303
rect 23581 33269 23615 33303
rect 23615 33269 23624 33303
rect 23572 33260 23624 33269
rect 25688 33260 25740 33312
rect 26884 33260 26936 33312
rect 27712 33260 27764 33312
rect 28264 33260 28316 33312
rect 28632 33328 28684 33380
rect 29460 33303 29512 33312
rect 29460 33269 29469 33303
rect 29469 33269 29503 33303
rect 29503 33269 29512 33303
rect 29460 33260 29512 33269
rect 29920 33260 29972 33312
rect 30472 33260 30524 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2872 33056 2924 33108
rect 3976 33056 4028 33108
rect 6276 33056 6328 33108
rect 6644 33056 6696 33108
rect 9220 33056 9272 33108
rect 9404 33099 9456 33108
rect 9404 33065 9413 33099
rect 9413 33065 9447 33099
rect 9447 33065 9456 33099
rect 9404 33056 9456 33065
rect 10508 33056 10560 33108
rect 10600 33056 10652 33108
rect 1768 32920 1820 32972
rect 1860 32895 1912 32904
rect 1860 32861 1869 32895
rect 1869 32861 1903 32895
rect 1903 32861 1912 32895
rect 1860 32852 1912 32861
rect 8668 32920 8720 32972
rect 2688 32852 2740 32904
rect 4528 32852 4580 32904
rect 940 32716 992 32768
rect 2136 32827 2188 32836
rect 2136 32793 2170 32827
rect 2170 32793 2188 32827
rect 2136 32784 2188 32793
rect 7012 32852 7064 32904
rect 7932 32852 7984 32904
rect 4712 32784 4764 32836
rect 8392 32852 8444 32904
rect 8852 32852 8904 32904
rect 11704 33056 11756 33108
rect 11244 33031 11296 33040
rect 11244 32997 11253 33031
rect 11253 32997 11287 33031
rect 11287 32997 11296 33031
rect 11244 32988 11296 32997
rect 9220 32852 9272 32904
rect 9772 32895 9824 32904
rect 9772 32861 9781 32895
rect 9781 32861 9815 32895
rect 9815 32861 9824 32895
rect 9772 32852 9824 32861
rect 12716 33056 12768 33108
rect 13360 33056 13412 33108
rect 13636 33056 13688 33108
rect 12256 32920 12308 32972
rect 12900 32920 12952 32972
rect 13268 32963 13320 32972
rect 13268 32929 13277 32963
rect 13277 32929 13311 32963
rect 13311 32929 13320 32963
rect 13268 32920 13320 32929
rect 3976 32759 4028 32768
rect 3976 32725 3985 32759
rect 3985 32725 4019 32759
rect 4019 32725 4028 32759
rect 3976 32716 4028 32725
rect 4068 32716 4120 32768
rect 5356 32716 5408 32768
rect 5908 32716 5960 32768
rect 7472 32716 7524 32768
rect 8300 32716 8352 32768
rect 8852 32716 8904 32768
rect 10324 32784 10376 32836
rect 11060 32852 11112 32904
rect 11612 32852 11664 32904
rect 11520 32784 11572 32836
rect 11796 32852 11848 32904
rect 12164 32852 12216 32904
rect 16304 33056 16356 33108
rect 16856 33056 16908 33108
rect 13912 32852 13964 32904
rect 14096 32895 14148 32904
rect 12348 32784 12400 32836
rect 12532 32784 12584 32836
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 15660 32852 15712 32904
rect 16396 32988 16448 33040
rect 19984 33056 20036 33108
rect 20076 33056 20128 33108
rect 21824 33056 21876 33108
rect 22192 33056 22244 33108
rect 24676 33056 24728 33108
rect 25964 33056 26016 33108
rect 26148 33056 26200 33108
rect 26424 33056 26476 33108
rect 26792 33056 26844 33108
rect 27896 33099 27948 33108
rect 27896 33065 27905 33099
rect 27905 33065 27939 33099
rect 27939 33065 27948 33099
rect 27896 33056 27948 33065
rect 28540 33099 28592 33108
rect 28540 33065 28549 33099
rect 28549 33065 28583 33099
rect 28583 33065 28592 33099
rect 28540 33056 28592 33065
rect 29276 33056 29328 33108
rect 29552 33056 29604 33108
rect 16212 32920 16264 32972
rect 18144 32988 18196 33040
rect 18604 32988 18656 33040
rect 15936 32852 15988 32904
rect 16488 32852 16540 32904
rect 17776 32852 17828 32904
rect 18420 32895 18472 32904
rect 18420 32861 18429 32895
rect 18429 32861 18463 32895
rect 18463 32861 18472 32895
rect 18420 32852 18472 32861
rect 19064 32852 19116 32904
rect 19156 32852 19208 32904
rect 19984 32920 20036 32972
rect 20168 32920 20220 32972
rect 20536 32920 20588 32972
rect 10692 32716 10744 32768
rect 12072 32716 12124 32768
rect 18512 32784 18564 32836
rect 20904 32895 20956 32904
rect 20904 32861 20913 32895
rect 20913 32861 20947 32895
rect 20947 32861 20956 32895
rect 20904 32852 20956 32861
rect 22376 32963 22428 32972
rect 22376 32929 22385 32963
rect 22385 32929 22419 32963
rect 22419 32929 22428 32963
rect 22376 32920 22428 32929
rect 23204 32852 23256 32904
rect 23940 32852 23992 32904
rect 24492 32895 24544 32904
rect 24492 32861 24501 32895
rect 24501 32861 24535 32895
rect 24535 32861 24544 32895
rect 24492 32852 24544 32861
rect 27344 32920 27396 32972
rect 12808 32759 12860 32768
rect 12808 32725 12817 32759
rect 12817 32725 12851 32759
rect 12851 32725 12860 32759
rect 12808 32716 12860 32725
rect 15660 32716 15712 32768
rect 16948 32716 17000 32768
rect 17040 32759 17092 32768
rect 17040 32725 17049 32759
rect 17049 32725 17083 32759
rect 17083 32725 17092 32759
rect 17040 32716 17092 32725
rect 17132 32716 17184 32768
rect 17868 32759 17920 32768
rect 17868 32725 17877 32759
rect 17877 32725 17911 32759
rect 17911 32725 17920 32759
rect 17868 32716 17920 32725
rect 19064 32759 19116 32768
rect 19064 32725 19073 32759
rect 19073 32725 19107 32759
rect 19107 32725 19116 32759
rect 19064 32716 19116 32725
rect 19984 32716 20036 32768
rect 20076 32716 20128 32768
rect 24860 32784 24912 32836
rect 25504 32852 25556 32904
rect 25780 32852 25832 32904
rect 26240 32852 26292 32904
rect 26424 32852 26476 32904
rect 26976 32852 27028 32904
rect 27620 32920 27672 32972
rect 28908 32920 28960 32972
rect 29276 32920 29328 32972
rect 29368 32920 29420 32972
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 27712 32895 27764 32904
rect 27712 32861 27721 32895
rect 27721 32861 27755 32895
rect 27755 32861 27764 32895
rect 27712 32852 27764 32861
rect 27804 32895 27856 32904
rect 27804 32861 27813 32895
rect 27813 32861 27847 32895
rect 27847 32861 27856 32895
rect 27804 32852 27856 32861
rect 28448 32852 28500 32904
rect 29092 32895 29144 32904
rect 29092 32861 29101 32895
rect 29101 32861 29135 32895
rect 29135 32861 29144 32895
rect 29092 32852 29144 32861
rect 29736 32852 29788 32904
rect 30380 32852 30432 32904
rect 24584 32716 24636 32768
rect 25044 32759 25096 32768
rect 25044 32725 25053 32759
rect 25053 32725 25087 32759
rect 25087 32725 25096 32759
rect 25044 32716 25096 32725
rect 26424 32716 26476 32768
rect 29000 32784 29052 32836
rect 29276 32784 29328 32836
rect 29368 32827 29420 32836
rect 29368 32793 29377 32827
rect 29377 32793 29411 32827
rect 29411 32793 29420 32827
rect 29368 32784 29420 32793
rect 29644 32784 29696 32836
rect 26700 32716 26752 32768
rect 26884 32716 26936 32768
rect 27252 32759 27304 32768
rect 27252 32725 27261 32759
rect 27261 32725 27295 32759
rect 27295 32725 27304 32759
rect 27252 32716 27304 32725
rect 28172 32716 28224 32768
rect 28724 32716 28776 32768
rect 28816 32759 28868 32768
rect 28816 32725 28825 32759
rect 28825 32725 28859 32759
rect 28859 32725 28868 32759
rect 28816 32716 28868 32725
rect 29920 32716 29972 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 7380 32512 7432 32564
rect 8300 32555 8352 32564
rect 8300 32521 8309 32555
rect 8309 32521 8343 32555
rect 8343 32521 8352 32555
rect 8300 32512 8352 32521
rect 1676 32376 1728 32428
rect 1492 32308 1544 32360
rect 2964 32351 3016 32360
rect 2964 32317 2973 32351
rect 2973 32317 3007 32351
rect 3007 32317 3016 32351
rect 2964 32308 3016 32317
rect 5632 32376 5684 32428
rect 7380 32376 7432 32428
rect 9312 32512 9364 32564
rect 8668 32444 8720 32496
rect 9220 32444 9272 32496
rect 11152 32512 11204 32564
rect 11704 32512 11756 32564
rect 13636 32555 13688 32564
rect 13636 32521 13645 32555
rect 13645 32521 13679 32555
rect 13679 32521 13688 32555
rect 13636 32512 13688 32521
rect 14924 32512 14976 32564
rect 3516 32215 3568 32224
rect 3516 32181 3525 32215
rect 3525 32181 3559 32215
rect 3559 32181 3568 32215
rect 3516 32172 3568 32181
rect 4068 32172 4120 32224
rect 5908 32240 5960 32292
rect 6276 32240 6328 32292
rect 7840 32308 7892 32360
rect 8208 32240 8260 32292
rect 7012 32172 7064 32224
rect 10324 32376 10376 32428
rect 13544 32444 13596 32496
rect 15568 32555 15620 32564
rect 15568 32521 15577 32555
rect 15577 32521 15611 32555
rect 15611 32521 15620 32555
rect 15568 32512 15620 32521
rect 15660 32555 15712 32564
rect 15660 32521 15669 32555
rect 15669 32521 15703 32555
rect 15703 32521 15712 32555
rect 15660 32512 15712 32521
rect 15936 32512 15988 32564
rect 13912 32376 13964 32428
rect 14004 32419 14056 32428
rect 14004 32385 14013 32419
rect 14013 32385 14047 32419
rect 14047 32385 14056 32419
rect 14004 32376 14056 32385
rect 14280 32419 14332 32428
rect 14280 32385 14289 32419
rect 14289 32385 14323 32419
rect 14323 32385 14332 32419
rect 14280 32376 14332 32385
rect 14372 32419 14424 32428
rect 14372 32385 14381 32419
rect 14381 32385 14415 32419
rect 14415 32385 14424 32419
rect 14372 32376 14424 32385
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 14556 32419 14608 32428
rect 14556 32385 14591 32419
rect 14591 32385 14608 32419
rect 14556 32376 14608 32385
rect 8576 32351 8628 32360
rect 8576 32317 8585 32351
rect 8585 32317 8619 32351
rect 8619 32317 8628 32351
rect 8576 32308 8628 32317
rect 9312 32308 9364 32360
rect 9496 32351 9548 32360
rect 9496 32317 9505 32351
rect 9505 32317 9539 32351
rect 9539 32317 9548 32351
rect 9496 32308 9548 32317
rect 10232 32308 10284 32360
rect 10508 32308 10560 32360
rect 9128 32283 9180 32292
rect 9128 32249 9137 32283
rect 9137 32249 9171 32283
rect 9171 32249 9180 32283
rect 9128 32240 9180 32249
rect 10324 32215 10376 32224
rect 10324 32181 10333 32215
rect 10333 32181 10367 32215
rect 10367 32181 10376 32215
rect 10324 32172 10376 32181
rect 10968 32283 11020 32292
rect 10968 32249 10977 32283
rect 10977 32249 11011 32283
rect 11011 32249 11020 32283
rect 10968 32240 11020 32249
rect 14740 32351 14792 32360
rect 14740 32317 14749 32351
rect 14749 32317 14783 32351
rect 14783 32317 14792 32351
rect 14740 32308 14792 32317
rect 16028 32444 16080 32496
rect 16304 32512 16356 32564
rect 16488 32555 16540 32564
rect 16488 32521 16497 32555
rect 16497 32521 16531 32555
rect 16531 32521 16540 32555
rect 16488 32512 16540 32521
rect 17040 32512 17092 32564
rect 17868 32512 17920 32564
rect 20076 32512 20128 32564
rect 20444 32512 20496 32564
rect 20720 32512 20772 32564
rect 22468 32555 22520 32564
rect 22468 32521 22477 32555
rect 22477 32521 22511 32555
rect 22511 32521 22520 32555
rect 22468 32512 22520 32521
rect 24492 32512 24544 32564
rect 24860 32555 24912 32564
rect 24860 32521 24869 32555
rect 24869 32521 24903 32555
rect 24903 32521 24912 32555
rect 24860 32512 24912 32521
rect 25044 32512 25096 32564
rect 15660 32376 15712 32428
rect 15936 32376 15988 32428
rect 16764 32444 16816 32496
rect 19432 32444 19484 32496
rect 20904 32444 20956 32496
rect 18512 32376 18564 32428
rect 19248 32376 19300 32428
rect 16580 32308 16632 32360
rect 16948 32308 17000 32360
rect 17224 32351 17276 32360
rect 17224 32317 17233 32351
rect 17233 32317 17267 32351
rect 17267 32317 17276 32351
rect 17224 32308 17276 32317
rect 19340 32308 19392 32360
rect 19984 32419 20036 32428
rect 19984 32385 19993 32419
rect 19993 32385 20027 32419
rect 20027 32385 20036 32419
rect 19984 32376 20036 32385
rect 20444 32376 20496 32428
rect 12072 32215 12124 32224
rect 12072 32181 12081 32215
rect 12081 32181 12115 32215
rect 12115 32181 12124 32215
rect 12072 32172 12124 32181
rect 13728 32172 13780 32224
rect 17960 32240 18012 32292
rect 20628 32351 20680 32360
rect 20628 32317 20637 32351
rect 20637 32317 20671 32351
rect 20671 32317 20680 32351
rect 20628 32308 20680 32317
rect 20812 32419 20864 32428
rect 20812 32385 20821 32419
rect 20821 32385 20855 32419
rect 20855 32385 20864 32419
rect 26424 32444 26476 32496
rect 20812 32376 20864 32385
rect 23756 32376 23808 32428
rect 20996 32308 21048 32360
rect 22100 32308 22152 32360
rect 23848 32308 23900 32360
rect 24124 32376 24176 32428
rect 24308 32351 24360 32360
rect 24308 32317 24317 32351
rect 24317 32317 24351 32351
rect 24351 32317 24360 32351
rect 24308 32308 24360 32317
rect 24584 32419 24636 32428
rect 24584 32385 24593 32419
rect 24593 32385 24627 32419
rect 24627 32385 24636 32419
rect 24584 32376 24636 32385
rect 24860 32376 24912 32428
rect 24952 32376 25004 32428
rect 25412 32376 25464 32428
rect 25504 32419 25556 32428
rect 25504 32385 25513 32419
rect 25513 32385 25547 32419
rect 25547 32385 25556 32419
rect 25504 32376 25556 32385
rect 25872 32376 25924 32428
rect 26056 32419 26108 32428
rect 26056 32385 26065 32419
rect 26065 32385 26099 32419
rect 26099 32385 26108 32419
rect 26056 32376 26108 32385
rect 26240 32419 26292 32428
rect 26240 32385 26249 32419
rect 26249 32385 26283 32419
rect 26283 32385 26292 32419
rect 26240 32376 26292 32385
rect 26884 32512 26936 32564
rect 27344 32512 27396 32564
rect 28264 32512 28316 32564
rect 28724 32512 28776 32564
rect 29460 32512 29512 32564
rect 29644 32555 29696 32564
rect 29644 32521 29653 32555
rect 29653 32521 29687 32555
rect 29687 32521 29696 32555
rect 29644 32512 29696 32521
rect 30012 32512 30064 32564
rect 16396 32172 16448 32224
rect 16672 32172 16724 32224
rect 18604 32172 18656 32224
rect 24124 32240 24176 32292
rect 24676 32240 24728 32292
rect 25136 32351 25188 32360
rect 25136 32317 25145 32351
rect 25145 32317 25179 32351
rect 25179 32317 25188 32351
rect 25136 32308 25188 32317
rect 18972 32172 19024 32224
rect 20076 32172 20128 32224
rect 20352 32172 20404 32224
rect 21272 32215 21324 32224
rect 21272 32181 21281 32215
rect 21281 32181 21315 32215
rect 21315 32181 21324 32215
rect 21272 32172 21324 32181
rect 22008 32215 22060 32224
rect 22008 32181 22017 32215
rect 22017 32181 22051 32215
rect 22051 32181 22060 32215
rect 22008 32172 22060 32181
rect 23940 32215 23992 32224
rect 23940 32181 23949 32215
rect 23949 32181 23983 32215
rect 23983 32181 23992 32215
rect 23940 32172 23992 32181
rect 25228 32172 25280 32224
rect 25596 32172 25648 32224
rect 26332 32215 26384 32224
rect 26332 32181 26341 32215
rect 26341 32181 26375 32215
rect 26375 32181 26384 32215
rect 26332 32172 26384 32181
rect 26516 32283 26568 32292
rect 26516 32249 26525 32283
rect 26525 32249 26559 32283
rect 26559 32249 26568 32283
rect 26516 32240 26568 32249
rect 26884 32376 26936 32428
rect 27252 32376 27304 32428
rect 27804 32376 27856 32428
rect 28172 32419 28224 32428
rect 28172 32385 28181 32419
rect 28181 32385 28215 32419
rect 28215 32385 28224 32419
rect 28172 32376 28224 32385
rect 28356 32419 28408 32428
rect 28356 32385 28365 32419
rect 28365 32385 28399 32419
rect 28399 32385 28408 32419
rect 28356 32376 28408 32385
rect 26976 32308 27028 32360
rect 27344 32308 27396 32360
rect 27528 32351 27580 32360
rect 27528 32317 27537 32351
rect 27537 32317 27571 32351
rect 27571 32317 27580 32351
rect 28724 32376 28776 32428
rect 29000 32376 29052 32428
rect 27528 32308 27580 32317
rect 28816 32308 28868 32360
rect 26976 32215 27028 32224
rect 26976 32181 26985 32215
rect 26985 32181 27019 32215
rect 27019 32181 27028 32215
rect 26976 32172 27028 32181
rect 27988 32283 28040 32292
rect 27988 32249 27997 32283
rect 27997 32249 28031 32283
rect 28031 32249 28040 32283
rect 27988 32240 28040 32249
rect 30012 32419 30064 32428
rect 30012 32385 30021 32419
rect 30021 32385 30055 32419
rect 30055 32385 30064 32419
rect 30012 32376 30064 32385
rect 30748 32512 30800 32564
rect 32220 32512 32272 32564
rect 33048 32444 33100 32496
rect 30380 32376 30432 32428
rect 31392 32376 31444 32428
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 30472 32240 30524 32292
rect 29368 32172 29420 32224
rect 30840 32172 30892 32224
rect 32128 32215 32180 32224
rect 32128 32181 32137 32215
rect 32137 32181 32171 32215
rect 32171 32181 32180 32215
rect 32128 32172 32180 32181
rect 32772 32172 32824 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1860 31968 1912 32020
rect 3516 31968 3568 32020
rect 4712 31968 4764 32020
rect 4896 31968 4948 32020
rect 5356 31968 5408 32020
rect 4344 31875 4396 31884
rect 4344 31841 4353 31875
rect 4353 31841 4387 31875
rect 4387 31841 4396 31875
rect 4344 31832 4396 31841
rect 4896 31832 4948 31884
rect 7380 32011 7432 32020
rect 7380 31977 7389 32011
rect 7389 31977 7423 32011
rect 7423 31977 7432 32011
rect 7380 31968 7432 31977
rect 8576 31968 8628 32020
rect 9312 31968 9364 32020
rect 11796 31968 11848 32020
rect 12256 31968 12308 32020
rect 11612 31900 11664 31952
rect 14188 31968 14240 32020
rect 14280 31968 14332 32020
rect 16580 31968 16632 32020
rect 17960 31968 18012 32020
rect 5356 31875 5408 31884
rect 5356 31841 5365 31875
rect 5365 31841 5399 31875
rect 5399 31841 5408 31875
rect 5356 31832 5408 31841
rect 5448 31832 5500 31884
rect 6368 31807 6420 31816
rect 6368 31773 6377 31807
rect 6377 31773 6411 31807
rect 6411 31773 6420 31807
rect 6368 31764 6420 31773
rect 7012 31832 7064 31884
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 7564 31764 7616 31816
rect 8024 31807 8076 31816
rect 8024 31773 8033 31807
rect 8033 31773 8067 31807
rect 8067 31773 8076 31807
rect 8024 31764 8076 31773
rect 8208 31764 8260 31816
rect 9588 31764 9640 31816
rect 10968 31764 11020 31816
rect 12992 31900 13044 31952
rect 13544 31900 13596 31952
rect 14556 31832 14608 31884
rect 12348 31764 12400 31816
rect 15476 31832 15528 31884
rect 16028 31832 16080 31884
rect 3424 31739 3476 31748
rect 3424 31705 3433 31739
rect 3433 31705 3467 31739
rect 3467 31705 3476 31739
rect 3424 31696 3476 31705
rect 4160 31739 4212 31748
rect 4160 31705 4169 31739
rect 4169 31705 4203 31739
rect 4203 31705 4212 31739
rect 4160 31696 4212 31705
rect 5908 31696 5960 31748
rect 8484 31696 8536 31748
rect 15752 31764 15804 31816
rect 18052 31900 18104 31952
rect 18144 31875 18196 31884
rect 18144 31841 18153 31875
rect 18153 31841 18187 31875
rect 18187 31841 18196 31875
rect 18144 31832 18196 31841
rect 18512 31968 18564 32020
rect 19064 31968 19116 32020
rect 19616 31968 19668 32020
rect 20260 31968 20312 32020
rect 19156 31900 19208 31952
rect 19432 31832 19484 31884
rect 3884 31628 3936 31680
rect 4988 31628 5040 31680
rect 5172 31671 5224 31680
rect 5172 31637 5181 31671
rect 5181 31637 5215 31671
rect 5215 31637 5224 31671
rect 5172 31628 5224 31637
rect 7472 31628 7524 31680
rect 8760 31671 8812 31680
rect 8760 31637 8769 31671
rect 8769 31637 8803 31671
rect 8803 31637 8812 31671
rect 8760 31628 8812 31637
rect 9496 31628 9548 31680
rect 10048 31628 10100 31680
rect 12072 31628 12124 31680
rect 13544 31671 13596 31680
rect 13544 31637 13553 31671
rect 13553 31637 13587 31671
rect 13587 31637 13596 31671
rect 13544 31628 13596 31637
rect 13728 31628 13780 31680
rect 14188 31628 14240 31680
rect 14464 31628 14516 31680
rect 15476 31696 15528 31748
rect 16672 31739 16724 31748
rect 16672 31705 16706 31739
rect 16706 31705 16724 31739
rect 16672 31696 16724 31705
rect 16764 31696 16816 31748
rect 17592 31696 17644 31748
rect 19892 31807 19944 31816
rect 19892 31773 19926 31807
rect 19926 31773 19944 31807
rect 19892 31764 19944 31773
rect 24676 31968 24728 32020
rect 20996 31943 21048 31952
rect 20996 31909 21005 31943
rect 21005 31909 21039 31943
rect 21039 31909 21048 31943
rect 20996 31900 21048 31909
rect 20904 31832 20956 31884
rect 22100 31875 22152 31884
rect 22100 31841 22109 31875
rect 22109 31841 22143 31875
rect 22143 31841 22152 31875
rect 22100 31832 22152 31841
rect 15568 31628 15620 31680
rect 15752 31628 15804 31680
rect 16396 31628 16448 31680
rect 20260 31696 20312 31748
rect 20536 31696 20588 31748
rect 21272 31696 21324 31748
rect 23296 31764 23348 31816
rect 25136 31943 25188 31952
rect 25136 31909 25145 31943
rect 25145 31909 25179 31943
rect 25179 31909 25188 31943
rect 25136 31900 25188 31909
rect 26240 31968 26292 32020
rect 26792 31968 26844 32020
rect 26332 31900 26384 31952
rect 23848 31832 23900 31884
rect 24400 31807 24452 31816
rect 24400 31773 24409 31807
rect 24409 31773 24443 31807
rect 24443 31773 24452 31807
rect 24400 31764 24452 31773
rect 24768 31764 24820 31816
rect 26240 31832 26292 31884
rect 25228 31764 25280 31816
rect 25780 31764 25832 31816
rect 25872 31764 25924 31816
rect 26148 31764 26200 31816
rect 27804 31900 27856 31952
rect 27988 31900 28040 31952
rect 30104 31900 30156 31952
rect 26884 31875 26936 31884
rect 26884 31841 26893 31875
rect 26893 31841 26927 31875
rect 26927 31841 26936 31875
rect 26884 31832 26936 31841
rect 27344 31832 27396 31884
rect 28632 31832 28684 31884
rect 29092 31832 29144 31884
rect 23664 31696 23716 31748
rect 19524 31628 19576 31680
rect 21088 31671 21140 31680
rect 21088 31637 21097 31671
rect 21097 31637 21131 31671
rect 21131 31637 21140 31671
rect 21088 31628 21140 31637
rect 21456 31628 21508 31680
rect 21548 31628 21600 31680
rect 21916 31671 21968 31680
rect 21916 31637 21925 31671
rect 21925 31637 21959 31671
rect 21959 31637 21968 31671
rect 21916 31628 21968 31637
rect 23480 31628 23532 31680
rect 25596 31628 25648 31680
rect 26792 31807 26844 31816
rect 26792 31773 26801 31807
rect 26801 31773 26835 31807
rect 26835 31773 26844 31807
rect 26792 31764 26844 31773
rect 27068 31764 27120 31816
rect 27252 31696 27304 31748
rect 26976 31628 27028 31680
rect 27068 31628 27120 31680
rect 27620 31764 27672 31816
rect 28080 31764 28132 31816
rect 28816 31807 28868 31816
rect 28816 31773 28825 31807
rect 28825 31773 28859 31807
rect 28859 31773 28868 31807
rect 28816 31764 28868 31773
rect 28908 31807 28960 31816
rect 28908 31773 28917 31807
rect 28917 31773 28951 31807
rect 28951 31773 28960 31807
rect 28908 31764 28960 31773
rect 29552 31764 29604 31816
rect 31392 32011 31444 32020
rect 31392 31977 31401 32011
rect 31401 31977 31435 32011
rect 31435 31977 31444 32011
rect 31392 31968 31444 31977
rect 33048 32011 33100 32020
rect 33048 31977 33057 32011
rect 33057 31977 33091 32011
rect 33091 31977 33100 32011
rect 33048 31968 33100 31977
rect 30840 31875 30892 31884
rect 30840 31841 30849 31875
rect 30849 31841 30883 31875
rect 30883 31841 30892 31875
rect 30840 31832 30892 31841
rect 31024 31832 31076 31884
rect 32220 31875 32272 31884
rect 32220 31841 32229 31875
rect 32229 31841 32263 31875
rect 32263 31841 32272 31875
rect 32220 31832 32272 31841
rect 27712 31696 27764 31748
rect 28172 31628 28224 31680
rect 29092 31628 29144 31680
rect 29368 31628 29420 31680
rect 32404 31807 32456 31816
rect 32404 31773 32413 31807
rect 32413 31773 32447 31807
rect 32447 31773 32456 31807
rect 32404 31764 32456 31773
rect 30380 31628 30432 31680
rect 32128 31671 32180 31680
rect 32128 31637 32137 31671
rect 32137 31637 32171 31671
rect 32171 31637 32180 31671
rect 32128 31628 32180 31637
rect 32220 31628 32272 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2964 31424 3016 31476
rect 6828 31467 6880 31476
rect 6828 31433 6837 31467
rect 6837 31433 6871 31467
rect 6871 31433 6880 31467
rect 6828 31424 6880 31433
rect 3148 31356 3200 31408
rect 5448 31356 5500 31408
rect 6920 31356 6972 31408
rect 7564 31356 7616 31408
rect 7748 31356 7800 31408
rect 1952 31331 2004 31340
rect 1952 31297 1961 31331
rect 1961 31297 1995 31331
rect 1995 31297 2004 31331
rect 1952 31288 2004 31297
rect 2504 31288 2556 31340
rect 3884 31288 3936 31340
rect 4896 31331 4948 31340
rect 4896 31297 4905 31331
rect 4905 31297 4939 31331
rect 4939 31297 4948 31331
rect 4896 31288 4948 31297
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 4988 31288 5040 31297
rect 4068 31152 4120 31204
rect 4344 31263 4396 31272
rect 4344 31229 4353 31263
rect 4353 31229 4387 31263
rect 4387 31229 4396 31263
rect 4344 31220 4396 31229
rect 4804 31220 4856 31272
rect 6460 31288 6512 31340
rect 7104 31331 7156 31340
rect 7104 31297 7113 31331
rect 7113 31297 7147 31331
rect 7147 31297 7156 31331
rect 7104 31288 7156 31297
rect 8484 31467 8536 31476
rect 8484 31433 8493 31467
rect 8493 31433 8527 31467
rect 8527 31433 8536 31467
rect 8484 31424 8536 31433
rect 10140 31424 10192 31476
rect 11520 31424 11572 31476
rect 13544 31424 13596 31476
rect 8116 31399 8168 31408
rect 8116 31365 8125 31399
rect 8125 31365 8159 31399
rect 8159 31365 8168 31399
rect 8116 31356 8168 31365
rect 5540 31263 5592 31272
rect 5540 31229 5549 31263
rect 5549 31229 5583 31263
rect 5583 31229 5592 31263
rect 5540 31220 5592 31229
rect 7472 31263 7524 31272
rect 7472 31229 7481 31263
rect 7481 31229 7515 31263
rect 7515 31229 7524 31263
rect 7472 31220 7524 31229
rect 8208 31331 8260 31340
rect 8208 31297 8217 31331
rect 8217 31297 8251 31331
rect 8251 31297 8260 31331
rect 8208 31288 8260 31297
rect 8760 31288 8812 31340
rect 8668 31152 8720 31204
rect 8944 31331 8996 31340
rect 8944 31297 8953 31331
rect 8953 31297 8987 31331
rect 8987 31297 8996 31331
rect 8944 31288 8996 31297
rect 9588 31331 9640 31340
rect 9588 31297 9597 31331
rect 9597 31297 9631 31331
rect 9631 31297 9640 31331
rect 9588 31288 9640 31297
rect 11612 31288 11664 31340
rect 13728 31288 13780 31340
rect 15476 31356 15528 31408
rect 9312 31263 9364 31272
rect 9312 31229 9321 31263
rect 9321 31229 9355 31263
rect 9355 31229 9364 31263
rect 9312 31220 9364 31229
rect 9864 31263 9916 31272
rect 9864 31229 9873 31263
rect 9873 31229 9907 31263
rect 9907 31229 9916 31263
rect 9864 31220 9916 31229
rect 14280 31220 14332 31272
rect 17224 31424 17276 31476
rect 17868 31467 17920 31476
rect 17868 31433 17877 31467
rect 17877 31433 17911 31467
rect 17911 31433 17920 31467
rect 17868 31424 17920 31433
rect 18420 31467 18472 31476
rect 18420 31433 18429 31467
rect 18429 31433 18463 31467
rect 18463 31433 18472 31467
rect 18420 31424 18472 31433
rect 18604 31424 18656 31476
rect 15660 31356 15712 31408
rect 16028 31220 16080 31272
rect 16396 31220 16448 31272
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 17868 31288 17920 31340
rect 18328 31356 18380 31408
rect 18788 31399 18840 31408
rect 18788 31365 18797 31399
rect 18797 31365 18831 31399
rect 18831 31365 18840 31399
rect 18788 31356 18840 31365
rect 19248 31424 19300 31476
rect 19423 31424 19475 31476
rect 19984 31424 20036 31476
rect 20536 31424 20588 31476
rect 18512 31288 18564 31340
rect 19156 31331 19208 31340
rect 19156 31297 19165 31331
rect 19165 31297 19199 31331
rect 19199 31297 19208 31331
rect 19156 31288 19208 31297
rect 17224 31220 17276 31272
rect 18052 31220 18104 31272
rect 19064 31263 19116 31272
rect 19064 31229 19073 31263
rect 19073 31229 19107 31263
rect 19107 31229 19116 31263
rect 19064 31220 19116 31229
rect 19708 31288 19760 31340
rect 19984 31288 20036 31340
rect 20076 31331 20128 31340
rect 20076 31297 20085 31331
rect 20085 31297 20119 31331
rect 20119 31297 20128 31331
rect 20076 31288 20128 31297
rect 21088 31356 21140 31408
rect 21180 31356 21232 31408
rect 23480 31424 23532 31476
rect 23664 31467 23716 31476
rect 23664 31433 23673 31467
rect 23673 31433 23707 31467
rect 23707 31433 23716 31467
rect 23664 31424 23716 31433
rect 24400 31467 24452 31476
rect 24400 31433 24409 31467
rect 24409 31433 24443 31467
rect 24443 31433 24452 31467
rect 24400 31424 24452 31433
rect 24492 31467 24544 31476
rect 24492 31433 24501 31467
rect 24501 31433 24535 31467
rect 24535 31433 24544 31467
rect 24492 31424 24544 31433
rect 24584 31424 24636 31476
rect 20628 31288 20680 31340
rect 21824 31331 21876 31340
rect 21824 31297 21833 31331
rect 21833 31297 21867 31331
rect 21867 31297 21876 31331
rect 21824 31288 21876 31297
rect 22192 31288 22244 31340
rect 20444 31220 20496 31272
rect 3700 31084 3752 31136
rect 4620 31127 4672 31136
rect 4620 31093 4629 31127
rect 4629 31093 4663 31127
rect 4663 31093 4672 31127
rect 4620 31084 4672 31093
rect 7656 31084 7708 31136
rect 10784 31084 10836 31136
rect 10968 31127 11020 31136
rect 10968 31093 10977 31127
rect 10977 31093 11011 31127
rect 11011 31093 11020 31127
rect 10968 31084 11020 31093
rect 11704 31084 11756 31136
rect 12440 31084 12492 31136
rect 14556 31127 14608 31136
rect 14556 31093 14565 31127
rect 14565 31093 14599 31127
rect 14599 31093 14608 31127
rect 14556 31084 14608 31093
rect 14832 31084 14884 31136
rect 16396 31127 16448 31136
rect 16396 31093 16405 31127
rect 16405 31093 16439 31127
rect 16439 31093 16448 31127
rect 16396 31084 16448 31093
rect 17132 31084 17184 31136
rect 17868 31084 17920 31136
rect 18420 31084 18472 31136
rect 19156 31152 19208 31204
rect 19248 31152 19300 31204
rect 20812 31152 20864 31204
rect 20996 31263 21048 31272
rect 20996 31229 21005 31263
rect 21005 31229 21039 31263
rect 21039 31229 21048 31263
rect 20996 31220 21048 31229
rect 22560 31152 22612 31204
rect 22744 31331 22796 31340
rect 22744 31297 22753 31331
rect 22753 31297 22787 31331
rect 22787 31297 22796 31331
rect 22744 31288 22796 31297
rect 22928 31331 22980 31340
rect 22928 31297 22937 31331
rect 22937 31297 22971 31331
rect 22971 31297 22980 31331
rect 22928 31288 22980 31297
rect 23848 31288 23900 31340
rect 24768 31399 24820 31408
rect 24768 31365 24777 31399
rect 24777 31365 24811 31399
rect 24811 31365 24820 31399
rect 24768 31356 24820 31365
rect 24860 31399 24912 31408
rect 24860 31365 24869 31399
rect 24869 31365 24903 31399
rect 24903 31365 24912 31399
rect 24860 31356 24912 31365
rect 24952 31288 25004 31340
rect 25320 31356 25372 31408
rect 25872 31424 25924 31476
rect 25964 31424 26016 31476
rect 28356 31424 28408 31476
rect 24400 31220 24452 31272
rect 25596 31288 25648 31340
rect 26240 31356 26292 31408
rect 26332 31331 26384 31340
rect 26332 31297 26341 31331
rect 26341 31297 26375 31331
rect 26375 31297 26384 31331
rect 26332 31288 26384 31297
rect 26516 31288 26568 31340
rect 26700 31288 26752 31340
rect 27344 31288 27396 31340
rect 27620 31288 27672 31340
rect 27712 31288 27764 31340
rect 27804 31288 27856 31340
rect 28080 31331 28132 31340
rect 28080 31297 28089 31331
rect 28089 31297 28123 31331
rect 28123 31297 28132 31331
rect 28080 31288 28132 31297
rect 28356 31288 28408 31340
rect 26148 31263 26200 31272
rect 26148 31229 26157 31263
rect 26157 31229 26191 31263
rect 26191 31229 26200 31263
rect 26148 31220 26200 31229
rect 25964 31195 26016 31204
rect 25964 31161 25973 31195
rect 25973 31161 26007 31195
rect 26007 31161 26016 31195
rect 25964 31152 26016 31161
rect 28908 31220 28960 31272
rect 29552 31331 29604 31340
rect 29552 31297 29561 31331
rect 29561 31297 29595 31331
rect 29595 31297 29604 31331
rect 29552 31288 29604 31297
rect 32128 31288 32180 31340
rect 20536 31084 20588 31136
rect 21180 31084 21232 31136
rect 21364 31084 21416 31136
rect 21640 31127 21692 31136
rect 21640 31093 21649 31127
rect 21649 31093 21683 31127
rect 21683 31093 21692 31127
rect 21640 31084 21692 31093
rect 22284 31084 22336 31136
rect 23756 31084 23808 31136
rect 25320 31084 25372 31136
rect 25872 31084 25924 31136
rect 26056 31084 26108 31136
rect 26424 31084 26476 31136
rect 27252 31084 27304 31136
rect 27620 31084 27672 31136
rect 27896 31084 27948 31136
rect 28908 31084 28960 31136
rect 29552 31084 29604 31136
rect 30288 31084 30340 31136
rect 30932 31152 30984 31204
rect 30748 31084 30800 31136
rect 31024 31127 31076 31136
rect 31024 31093 31033 31127
rect 31033 31093 31067 31127
rect 31067 31093 31076 31127
rect 31024 31084 31076 31093
rect 31668 31084 31720 31136
rect 31760 31127 31812 31136
rect 31760 31093 31769 31127
rect 31769 31093 31803 31127
rect 31803 31093 31812 31127
rect 31760 31084 31812 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2504 30880 2556 30932
rect 3976 30923 4028 30932
rect 3976 30889 3985 30923
rect 3985 30889 4019 30923
rect 4019 30889 4028 30923
rect 3976 30880 4028 30889
rect 4068 30880 4120 30932
rect 4804 30880 4856 30932
rect 4988 30880 5040 30932
rect 6920 30880 6972 30932
rect 7104 30923 7156 30932
rect 7104 30889 7113 30923
rect 7113 30889 7147 30923
rect 7147 30889 7156 30923
rect 7104 30880 7156 30889
rect 8944 30880 8996 30932
rect 9864 30880 9916 30932
rect 10600 30880 10652 30932
rect 11612 30880 11664 30932
rect 13728 30880 13780 30932
rect 14556 30880 14608 30932
rect 15016 30880 15068 30932
rect 15476 30880 15528 30932
rect 1216 30744 1268 30796
rect 2044 30744 2096 30796
rect 5448 30812 5500 30864
rect 5540 30855 5592 30864
rect 5540 30821 5549 30855
rect 5549 30821 5583 30855
rect 5583 30821 5592 30855
rect 5540 30812 5592 30821
rect 6460 30812 6512 30864
rect 7656 30855 7708 30864
rect 7656 30821 7665 30855
rect 7665 30821 7699 30855
rect 7699 30821 7708 30855
rect 7656 30812 7708 30821
rect 8208 30812 8260 30864
rect 13636 30812 13688 30864
rect 14832 30812 14884 30864
rect 15108 30812 15160 30864
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 3424 30676 3476 30728
rect 3700 30676 3752 30728
rect 3976 30676 4028 30728
rect 4528 30676 4580 30728
rect 4620 30676 4672 30728
rect 4896 30676 4948 30728
rect 4988 30719 5040 30728
rect 4988 30685 4997 30719
rect 4997 30685 5031 30719
rect 5031 30685 5040 30719
rect 4988 30676 5040 30685
rect 3332 30651 3384 30660
rect 3332 30617 3341 30651
rect 3341 30617 3375 30651
rect 3375 30617 3384 30651
rect 3332 30608 3384 30617
rect 5356 30719 5408 30728
rect 5356 30685 5365 30719
rect 5365 30685 5399 30719
rect 5399 30685 5408 30719
rect 5356 30676 5408 30685
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 3056 30540 3108 30592
rect 3976 30540 4028 30592
rect 5264 30608 5316 30660
rect 7564 30719 7616 30728
rect 7564 30685 7573 30719
rect 7573 30685 7607 30719
rect 7607 30685 7616 30719
rect 7564 30676 7616 30685
rect 7748 30719 7800 30728
rect 7748 30685 7757 30719
rect 7757 30685 7791 30719
rect 7791 30685 7800 30719
rect 7748 30676 7800 30685
rect 8576 30744 8628 30796
rect 10600 30744 10652 30796
rect 10784 30744 10836 30796
rect 11888 30744 11940 30796
rect 12992 30744 13044 30796
rect 14924 30744 14976 30796
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 17316 30880 17368 30932
rect 17592 30880 17644 30932
rect 18144 30880 18196 30932
rect 18604 30880 18656 30932
rect 18696 30923 18748 30932
rect 18696 30889 18705 30923
rect 18705 30889 18739 30923
rect 18739 30889 18748 30923
rect 18696 30880 18748 30889
rect 9220 30719 9272 30728
rect 9220 30685 9229 30719
rect 9229 30685 9263 30719
rect 9263 30685 9272 30719
rect 9220 30676 9272 30685
rect 9496 30676 9548 30728
rect 10048 30719 10100 30728
rect 10048 30685 10057 30719
rect 10057 30685 10091 30719
rect 10091 30685 10100 30719
rect 10048 30676 10100 30685
rect 12164 30719 12216 30728
rect 12164 30685 12173 30719
rect 12173 30685 12207 30719
rect 12207 30685 12216 30719
rect 12164 30676 12216 30685
rect 12716 30719 12768 30728
rect 12716 30685 12725 30719
rect 12725 30685 12759 30719
rect 12759 30685 12768 30719
rect 12716 30676 12768 30685
rect 9312 30608 9364 30660
rect 10876 30608 10928 30660
rect 12072 30608 12124 30660
rect 12256 30608 12308 30660
rect 4528 30540 4580 30592
rect 6460 30540 6512 30592
rect 6920 30540 6972 30592
rect 7104 30540 7156 30592
rect 7840 30540 7892 30592
rect 8944 30540 8996 30592
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 18696 30744 18748 30796
rect 17316 30719 17368 30728
rect 17316 30685 17325 30719
rect 17325 30685 17359 30719
rect 17359 30685 17368 30719
rect 17316 30676 17368 30685
rect 17776 30719 17828 30728
rect 17776 30685 17785 30719
rect 17785 30685 17819 30719
rect 17819 30685 17828 30719
rect 17776 30676 17828 30685
rect 17960 30719 18012 30728
rect 17960 30685 17969 30719
rect 17969 30685 18003 30719
rect 18003 30685 18012 30719
rect 17960 30676 18012 30685
rect 13728 30540 13780 30592
rect 13912 30540 13964 30592
rect 14004 30540 14056 30592
rect 14372 30540 14424 30592
rect 14464 30583 14516 30592
rect 14464 30549 14473 30583
rect 14473 30549 14507 30583
rect 14507 30549 14516 30583
rect 14464 30540 14516 30549
rect 15660 30583 15712 30592
rect 15660 30549 15669 30583
rect 15669 30549 15703 30583
rect 15703 30549 15712 30583
rect 15660 30540 15712 30549
rect 17684 30608 17736 30660
rect 18328 30719 18380 30728
rect 18328 30685 18337 30719
rect 18337 30685 18371 30719
rect 18371 30685 18380 30719
rect 18328 30676 18380 30685
rect 18420 30676 18472 30728
rect 19340 30744 19392 30796
rect 19248 30719 19300 30728
rect 19248 30685 19257 30719
rect 19257 30685 19291 30719
rect 19291 30685 19300 30719
rect 19248 30676 19300 30685
rect 20444 30812 20496 30864
rect 22468 30880 22520 30932
rect 22928 30880 22980 30932
rect 24308 30880 24360 30932
rect 24400 30880 24452 30932
rect 24492 30880 24544 30932
rect 24584 30880 24636 30932
rect 23940 30812 23992 30864
rect 24124 30812 24176 30864
rect 20352 30744 20404 30796
rect 20720 30744 20772 30796
rect 20904 30787 20956 30796
rect 20904 30753 20913 30787
rect 20913 30753 20947 30787
rect 20947 30753 20956 30787
rect 20904 30744 20956 30753
rect 18512 30608 18564 30660
rect 18604 30608 18656 30660
rect 18788 30608 18840 30660
rect 19340 30608 19392 30660
rect 22008 30676 22060 30728
rect 23480 30744 23532 30796
rect 23572 30744 23624 30796
rect 24584 30744 24636 30796
rect 24676 30787 24728 30796
rect 24676 30753 24685 30787
rect 24685 30753 24719 30787
rect 24719 30753 24728 30787
rect 24676 30744 24728 30753
rect 24768 30787 24820 30796
rect 24768 30753 24777 30787
rect 24777 30753 24811 30787
rect 24811 30753 24820 30787
rect 24768 30744 24820 30753
rect 24952 30787 25004 30796
rect 24952 30753 24961 30787
rect 24961 30753 24995 30787
rect 24995 30753 25004 30787
rect 24952 30744 25004 30753
rect 23848 30719 23900 30728
rect 23848 30685 23857 30719
rect 23857 30685 23891 30719
rect 23891 30685 23900 30719
rect 23848 30676 23900 30685
rect 25780 30812 25832 30864
rect 25320 30719 25372 30728
rect 25320 30685 25329 30719
rect 25329 30685 25363 30719
rect 25363 30685 25372 30719
rect 25320 30676 25372 30685
rect 25412 30719 25464 30728
rect 25412 30685 25421 30719
rect 25421 30685 25455 30719
rect 25455 30685 25464 30719
rect 25412 30676 25464 30685
rect 26148 30880 26200 30932
rect 28172 30923 28224 30932
rect 28172 30889 28181 30923
rect 28181 30889 28215 30923
rect 28215 30889 28224 30923
rect 28172 30880 28224 30889
rect 28448 30923 28500 30932
rect 28448 30889 28457 30923
rect 28457 30889 28491 30923
rect 28491 30889 28500 30923
rect 28448 30880 28500 30889
rect 29552 30923 29604 30932
rect 29552 30889 29561 30923
rect 29561 30889 29595 30923
rect 29595 30889 29604 30923
rect 29552 30880 29604 30889
rect 32404 30880 32456 30932
rect 26332 30855 26384 30864
rect 26332 30821 26341 30855
rect 26341 30821 26375 30855
rect 26375 30821 26384 30855
rect 26332 30812 26384 30821
rect 26516 30812 26568 30864
rect 26976 30812 27028 30864
rect 27620 30812 27672 30864
rect 28724 30812 28776 30864
rect 20720 30608 20772 30660
rect 17132 30540 17184 30592
rect 19156 30540 19208 30592
rect 19248 30540 19300 30592
rect 20076 30540 20128 30592
rect 20444 30540 20496 30592
rect 20536 30583 20588 30592
rect 20536 30549 20545 30583
rect 20545 30549 20579 30583
rect 20579 30549 20588 30583
rect 20536 30540 20588 30549
rect 20904 30540 20956 30592
rect 22744 30540 22796 30592
rect 23112 30540 23164 30592
rect 24492 30608 24544 30660
rect 25044 30608 25096 30660
rect 23664 30540 23716 30592
rect 24400 30540 24452 30592
rect 24768 30540 24820 30592
rect 25504 30651 25556 30660
rect 25504 30617 25513 30651
rect 25513 30617 25547 30651
rect 25547 30617 25556 30651
rect 25504 30608 25556 30617
rect 26056 30608 26108 30660
rect 26700 30540 26752 30592
rect 27528 30787 27580 30796
rect 27528 30753 27537 30787
rect 27537 30753 27571 30787
rect 27571 30753 27580 30787
rect 27528 30744 27580 30753
rect 28632 30744 28684 30796
rect 28816 30744 28868 30796
rect 28448 30608 28500 30660
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 29276 30744 29328 30796
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 30472 30719 30524 30728
rect 30472 30685 30481 30719
rect 30481 30685 30515 30719
rect 30515 30685 30524 30719
rect 30472 30676 30524 30685
rect 30656 30608 30708 30660
rect 30932 30676 30984 30728
rect 32220 30676 32272 30728
rect 31760 30608 31812 30660
rect 33508 30676 33560 30728
rect 28816 30583 28868 30592
rect 28816 30549 28825 30583
rect 28825 30549 28859 30583
rect 28859 30549 28868 30583
rect 28816 30540 28868 30549
rect 30012 30540 30064 30592
rect 31392 30540 31444 30592
rect 31944 30540 31996 30592
rect 32312 30540 32364 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 2044 30379 2096 30388
rect 2044 30345 2053 30379
rect 2053 30345 2087 30379
rect 2087 30345 2096 30379
rect 2044 30336 2096 30345
rect 3332 30336 3384 30388
rect 2136 30243 2188 30252
rect 2136 30209 2145 30243
rect 2145 30209 2179 30243
rect 2179 30209 2188 30243
rect 2136 30200 2188 30209
rect 2412 30200 2464 30252
rect 2504 30243 2556 30252
rect 2504 30209 2513 30243
rect 2513 30209 2547 30243
rect 2547 30209 2556 30243
rect 2504 30200 2556 30209
rect 2872 30200 2924 30252
rect 3240 30268 3292 30320
rect 3976 30311 4028 30320
rect 3976 30277 3985 30311
rect 3985 30277 4019 30311
rect 4019 30277 4028 30311
rect 3976 30268 4028 30277
rect 4160 30268 4212 30320
rect 4804 30336 4856 30388
rect 4344 30311 4396 30320
rect 4344 30277 4353 30311
rect 4353 30277 4387 30311
rect 4387 30277 4396 30311
rect 4344 30268 4396 30277
rect 4712 30268 4764 30320
rect 5448 30379 5500 30388
rect 5448 30345 5457 30379
rect 5457 30345 5491 30379
rect 5491 30345 5500 30379
rect 5448 30336 5500 30345
rect 5632 30336 5684 30388
rect 6920 30379 6972 30388
rect 6920 30345 6929 30379
rect 6929 30345 6963 30379
rect 6963 30345 6972 30379
rect 6920 30336 6972 30345
rect 7840 30379 7892 30388
rect 7840 30345 7849 30379
rect 7849 30345 7883 30379
rect 7883 30345 7892 30379
rect 7840 30336 7892 30345
rect 8116 30336 8168 30388
rect 9588 30336 9640 30388
rect 9864 30336 9916 30388
rect 10600 30336 10652 30388
rect 10784 30336 10836 30388
rect 2688 30064 2740 30116
rect 3148 30200 3200 30252
rect 3516 30200 3568 30252
rect 4160 30132 4212 30184
rect 4528 30132 4580 30184
rect 3332 30064 3384 30116
rect 4252 30064 4304 30116
rect 4620 30064 4672 30116
rect 4896 30200 4948 30252
rect 5264 30268 5316 30320
rect 7104 30311 7156 30320
rect 7104 30277 7113 30311
rect 7113 30277 7147 30311
rect 7147 30277 7156 30311
rect 7104 30268 7156 30277
rect 11888 30336 11940 30388
rect 12164 30336 12216 30388
rect 12348 30336 12400 30388
rect 6184 30200 6236 30252
rect 5172 30175 5224 30184
rect 5172 30141 5181 30175
rect 5181 30141 5215 30175
rect 5215 30141 5224 30175
rect 5172 30132 5224 30141
rect 5356 30132 5408 30184
rect 6828 30200 6880 30252
rect 7748 30200 7800 30252
rect 5540 30064 5592 30116
rect 7564 30175 7616 30184
rect 7564 30141 7573 30175
rect 7573 30141 7607 30175
rect 7607 30141 7616 30175
rect 7564 30132 7616 30141
rect 8116 30132 8168 30184
rect 8208 30132 8260 30184
rect 8668 30243 8720 30252
rect 8668 30209 8677 30243
rect 8677 30209 8711 30243
rect 8711 30209 8720 30243
rect 8668 30200 8720 30209
rect 9220 30200 9272 30252
rect 9956 30200 10008 30252
rect 10416 30200 10468 30252
rect 10876 30200 10928 30252
rect 11336 30243 11388 30252
rect 11336 30209 11345 30243
rect 11345 30209 11379 30243
rect 11379 30209 11388 30243
rect 11336 30200 11388 30209
rect 11520 30243 11572 30252
rect 11520 30209 11529 30243
rect 11529 30209 11563 30243
rect 11563 30209 11572 30243
rect 11520 30200 11572 30209
rect 11612 30243 11664 30252
rect 11612 30209 11622 30243
rect 11622 30209 11656 30243
rect 11656 30209 11664 30243
rect 11612 30200 11664 30209
rect 11980 30200 12032 30252
rect 12992 30379 13044 30388
rect 12992 30345 13001 30379
rect 13001 30345 13035 30379
rect 13035 30345 13044 30379
rect 12992 30336 13044 30345
rect 9312 30132 9364 30184
rect 9496 30132 9548 30184
rect 2964 29996 3016 30048
rect 4160 29996 4212 30048
rect 5264 30039 5316 30048
rect 5264 30005 5273 30039
rect 5273 30005 5307 30039
rect 5307 30005 5316 30039
rect 5264 29996 5316 30005
rect 6368 29996 6420 30048
rect 7656 30039 7708 30048
rect 7656 30005 7665 30039
rect 7665 30005 7699 30039
rect 7699 30005 7708 30039
rect 7656 29996 7708 30005
rect 11336 30064 11388 30116
rect 12256 29996 12308 30048
rect 12440 30132 12492 30184
rect 14004 30336 14056 30388
rect 14280 30379 14332 30388
rect 14280 30345 14289 30379
rect 14289 30345 14323 30379
rect 14323 30345 14332 30379
rect 14280 30336 14332 30345
rect 15660 30336 15712 30388
rect 17776 30336 17828 30388
rect 14832 30268 14884 30320
rect 12532 30064 12584 30116
rect 12624 29996 12676 30048
rect 13084 30064 13136 30116
rect 15108 30200 15160 30252
rect 15476 30243 15528 30252
rect 15476 30209 15485 30243
rect 15485 30209 15519 30243
rect 15519 30209 15528 30243
rect 15476 30200 15528 30209
rect 15660 30200 15712 30252
rect 15936 30243 15988 30252
rect 15936 30209 15945 30243
rect 15945 30209 15979 30243
rect 15979 30209 15988 30243
rect 15936 30200 15988 30209
rect 16212 30268 16264 30320
rect 16948 30311 17000 30320
rect 16948 30277 16957 30311
rect 16957 30277 16991 30311
rect 16991 30277 17000 30311
rect 16948 30268 17000 30277
rect 18604 30268 18656 30320
rect 20720 30336 20772 30388
rect 22008 30336 22060 30388
rect 14188 30132 14240 30184
rect 14280 30064 14332 30116
rect 15200 30132 15252 30184
rect 16212 30132 16264 30184
rect 16488 30132 16540 30184
rect 17132 30200 17184 30252
rect 17500 30200 17552 30252
rect 17592 30243 17644 30252
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 17132 30064 17184 30116
rect 14004 29996 14056 30048
rect 17224 30039 17276 30048
rect 17224 30005 17233 30039
rect 17233 30005 17267 30039
rect 17267 30005 17276 30039
rect 17224 29996 17276 30005
rect 17684 29996 17736 30048
rect 17960 30200 18012 30252
rect 20352 30268 20404 30320
rect 20444 30268 20496 30320
rect 22928 30336 22980 30388
rect 23480 30336 23532 30388
rect 23940 30336 23992 30388
rect 25136 30336 25188 30388
rect 21088 30200 21140 30252
rect 19064 30064 19116 30116
rect 19156 30064 19208 30116
rect 19524 30064 19576 30116
rect 18328 29996 18380 30048
rect 18880 30039 18932 30048
rect 18880 30005 18889 30039
rect 18889 30005 18923 30039
rect 18923 30005 18932 30039
rect 18880 29996 18932 30005
rect 19340 29996 19392 30048
rect 19800 30175 19852 30184
rect 19800 30141 19809 30175
rect 19809 30141 19843 30175
rect 19843 30141 19852 30175
rect 19800 30132 19852 30141
rect 20812 30132 20864 30184
rect 21364 30200 21416 30252
rect 21640 30132 21692 30184
rect 20996 30064 21048 30116
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 22376 30132 22428 30184
rect 23296 30243 23348 30252
rect 23296 30209 23305 30243
rect 23305 30209 23339 30243
rect 23339 30209 23348 30243
rect 23296 30200 23348 30209
rect 24584 30268 24636 30320
rect 23664 30200 23716 30252
rect 23480 30132 23532 30184
rect 23848 30175 23900 30184
rect 23848 30141 23857 30175
rect 23857 30141 23891 30175
rect 23891 30141 23900 30175
rect 23848 30132 23900 30141
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 24768 30200 24820 30252
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 25412 30200 25464 30252
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 25596 30243 25648 30252
rect 25596 30209 25605 30243
rect 25605 30209 25639 30243
rect 25639 30209 25648 30243
rect 25596 30200 25648 30209
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 26516 30243 26568 30252
rect 26516 30209 26525 30243
rect 26525 30209 26559 30243
rect 26559 30209 26568 30243
rect 26516 30200 26568 30209
rect 26792 30200 26844 30252
rect 27712 30336 27764 30388
rect 28172 30336 28224 30388
rect 28816 30336 28868 30388
rect 29276 30336 29328 30388
rect 27436 30200 27488 30252
rect 28080 30268 28132 30320
rect 28540 30268 28592 30320
rect 30288 30336 30340 30388
rect 30748 30336 30800 30388
rect 33508 30379 33560 30388
rect 33508 30345 33517 30379
rect 33517 30345 33551 30379
rect 33551 30345 33560 30379
rect 33508 30336 33560 30345
rect 24124 30132 24176 30184
rect 22192 30064 22244 30116
rect 23296 30064 23348 30116
rect 25688 30132 25740 30184
rect 28356 30132 28408 30184
rect 28816 30200 28868 30252
rect 28908 30200 28960 30252
rect 29184 30243 29236 30252
rect 29184 30209 29193 30243
rect 29193 30209 29227 30243
rect 29227 30209 29236 30243
rect 29184 30200 29236 30209
rect 29460 30243 29512 30252
rect 29460 30209 29469 30243
rect 29469 30209 29503 30243
rect 29503 30209 29512 30243
rect 29460 30200 29512 30209
rect 30196 30311 30248 30320
rect 30196 30277 30205 30311
rect 30205 30277 30239 30311
rect 30239 30277 30248 30311
rect 30196 30268 30248 30277
rect 30472 30268 30524 30320
rect 31024 30268 31076 30320
rect 20076 29996 20128 30048
rect 22652 29996 22704 30048
rect 23480 30039 23532 30048
rect 23480 30005 23489 30039
rect 23489 30005 23523 30039
rect 23523 30005 23532 30039
rect 23480 29996 23532 30005
rect 23664 30039 23716 30048
rect 23664 30005 23673 30039
rect 23673 30005 23707 30039
rect 23707 30005 23716 30039
rect 23664 29996 23716 30005
rect 23756 30039 23808 30048
rect 23756 30005 23765 30039
rect 23765 30005 23799 30039
rect 23799 30005 23808 30039
rect 23756 29996 23808 30005
rect 23848 29996 23900 30048
rect 24308 29996 24360 30048
rect 25412 30107 25464 30116
rect 25412 30073 25421 30107
rect 25421 30073 25455 30107
rect 25455 30073 25464 30107
rect 25412 30064 25464 30073
rect 25780 30064 25832 30116
rect 26240 30107 26292 30116
rect 26240 30073 26249 30107
rect 26249 30073 26283 30107
rect 26283 30073 26292 30107
rect 26240 30064 26292 30073
rect 26884 30064 26936 30116
rect 25964 29996 26016 30048
rect 26056 29996 26108 30048
rect 26700 29996 26752 30048
rect 27068 29996 27120 30048
rect 27620 29996 27672 30048
rect 28448 29996 28500 30048
rect 28632 29996 28684 30048
rect 28724 29996 28776 30048
rect 31944 30268 31996 30320
rect 30472 30132 30524 30184
rect 31392 30243 31444 30252
rect 31392 30209 31401 30243
rect 31401 30209 31435 30243
rect 31435 30209 31444 30243
rect 31392 30200 31444 30209
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 31760 30243 31812 30252
rect 31760 30209 31769 30243
rect 31769 30209 31803 30243
rect 31803 30209 31812 30243
rect 31760 30200 31812 30209
rect 32220 30200 32272 30252
rect 30932 30132 30984 30184
rect 32036 30132 32088 30184
rect 30472 29996 30524 30048
rect 30564 30039 30616 30048
rect 30564 30005 30573 30039
rect 30573 30005 30607 30039
rect 30607 30005 30616 30039
rect 30564 29996 30616 30005
rect 30656 29996 30708 30048
rect 31944 30039 31996 30048
rect 31944 30005 31953 30039
rect 31953 30005 31987 30039
rect 31987 30005 31996 30039
rect 31944 29996 31996 30005
rect 32312 29996 32364 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2504 29792 2556 29844
rect 3240 29792 3292 29844
rect 3424 29792 3476 29844
rect 1584 29724 1636 29776
rect 2964 29724 3016 29776
rect 1216 29656 1268 29708
rect 2688 29656 2740 29708
rect 2044 29588 2096 29640
rect 2412 29588 2464 29640
rect 3516 29656 3568 29708
rect 3976 29656 4028 29708
rect 1860 29452 1912 29504
rect 2780 29452 2832 29504
rect 3332 29631 3384 29640
rect 3332 29597 3341 29631
rect 3341 29597 3375 29631
rect 3375 29597 3384 29631
rect 3332 29588 3384 29597
rect 3424 29631 3476 29640
rect 3424 29597 3433 29631
rect 3433 29597 3467 29631
rect 3467 29597 3476 29631
rect 3424 29588 3476 29597
rect 4712 29835 4764 29844
rect 4712 29801 4721 29835
rect 4721 29801 4755 29835
rect 4755 29801 4764 29835
rect 4712 29792 4764 29801
rect 5172 29792 5224 29844
rect 6184 29792 6236 29844
rect 4712 29588 4764 29640
rect 3976 29452 4028 29504
rect 4896 29452 4948 29504
rect 5264 29631 5316 29640
rect 5264 29597 5273 29631
rect 5273 29597 5307 29631
rect 5307 29597 5316 29631
rect 5264 29588 5316 29597
rect 6460 29724 6512 29776
rect 6828 29792 6880 29844
rect 8208 29835 8260 29844
rect 8208 29801 8217 29835
rect 8217 29801 8251 29835
rect 8251 29801 8260 29835
rect 8208 29792 8260 29801
rect 8576 29835 8628 29844
rect 8576 29801 8585 29835
rect 8585 29801 8619 29835
rect 8619 29801 8628 29835
rect 8576 29792 8628 29801
rect 8668 29792 8720 29844
rect 9220 29792 9272 29844
rect 10508 29792 10560 29844
rect 11612 29792 11664 29844
rect 11888 29792 11940 29844
rect 12440 29835 12492 29844
rect 12440 29801 12449 29835
rect 12449 29801 12483 29835
rect 12483 29801 12492 29835
rect 12440 29792 12492 29801
rect 14004 29792 14056 29844
rect 16212 29792 16264 29844
rect 17224 29792 17276 29844
rect 19064 29792 19116 29844
rect 21088 29792 21140 29844
rect 22192 29792 22244 29844
rect 22744 29792 22796 29844
rect 23664 29792 23716 29844
rect 25136 29792 25188 29844
rect 25228 29792 25280 29844
rect 25780 29792 25832 29844
rect 26792 29792 26844 29844
rect 27436 29792 27488 29844
rect 27712 29835 27764 29844
rect 27712 29801 27721 29835
rect 27721 29801 27755 29835
rect 27755 29801 27764 29835
rect 27712 29792 27764 29801
rect 27804 29835 27856 29844
rect 27804 29801 27813 29835
rect 27813 29801 27847 29835
rect 27847 29801 27856 29835
rect 27804 29792 27856 29801
rect 28264 29792 28316 29844
rect 28816 29792 28868 29844
rect 29092 29792 29144 29844
rect 30564 29792 30616 29844
rect 5080 29520 5132 29572
rect 6828 29631 6880 29640
rect 6828 29597 6837 29631
rect 6837 29597 6871 29631
rect 6871 29597 6880 29631
rect 6828 29588 6880 29597
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 7012 29520 7064 29572
rect 6460 29452 6512 29504
rect 7840 29588 7892 29640
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 11244 29656 11296 29708
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 9956 29588 10008 29640
rect 10784 29588 10836 29640
rect 12256 29656 12308 29708
rect 12808 29724 12860 29776
rect 12716 29656 12768 29708
rect 13360 29699 13412 29708
rect 13360 29665 13369 29699
rect 13369 29665 13403 29699
rect 13403 29665 13412 29699
rect 13360 29656 13412 29665
rect 11152 29520 11204 29572
rect 10232 29452 10284 29504
rect 10324 29495 10376 29504
rect 10324 29461 10333 29495
rect 10333 29461 10367 29495
rect 10367 29461 10376 29495
rect 10324 29452 10376 29461
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 11980 29631 12032 29640
rect 11980 29597 11989 29631
rect 11989 29597 12023 29631
rect 12023 29597 12032 29631
rect 11980 29588 12032 29597
rect 12992 29588 13044 29640
rect 13176 29631 13228 29640
rect 13176 29597 13185 29631
rect 13185 29597 13219 29631
rect 13219 29597 13228 29631
rect 14464 29656 14516 29708
rect 14648 29656 14700 29708
rect 14832 29656 14884 29708
rect 13176 29588 13228 29597
rect 12164 29563 12216 29572
rect 12164 29529 12173 29563
rect 12173 29529 12207 29563
rect 12207 29529 12216 29563
rect 12164 29520 12216 29529
rect 12348 29520 12400 29572
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14924 29631 14976 29640
rect 14924 29597 14933 29631
rect 14933 29597 14967 29631
rect 14967 29597 14976 29631
rect 15476 29724 15528 29776
rect 14924 29588 14976 29597
rect 12716 29495 12768 29504
rect 12716 29461 12725 29495
rect 12725 29461 12759 29495
rect 12759 29461 12768 29495
rect 12716 29452 12768 29461
rect 13544 29452 13596 29504
rect 15568 29631 15620 29640
rect 15568 29597 15575 29631
rect 15575 29597 15620 29631
rect 15568 29588 15620 29597
rect 15844 29631 15896 29640
rect 15844 29597 15858 29631
rect 15858 29597 15892 29631
rect 15892 29597 15896 29631
rect 16764 29656 16816 29708
rect 20536 29656 20588 29708
rect 15844 29588 15896 29597
rect 16120 29520 16172 29572
rect 16488 29452 16540 29504
rect 17592 29588 17644 29640
rect 17776 29520 17828 29572
rect 18512 29520 18564 29572
rect 19800 29588 19852 29640
rect 18328 29452 18380 29504
rect 20812 29520 20864 29572
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 21180 29631 21232 29640
rect 21180 29597 21189 29631
rect 21189 29597 21223 29631
rect 21223 29597 21232 29631
rect 21180 29588 21232 29597
rect 22468 29724 22520 29776
rect 22284 29656 22336 29708
rect 24952 29724 25004 29776
rect 26700 29724 26752 29776
rect 31852 29792 31904 29844
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 22744 29631 22796 29640
rect 22744 29597 22753 29631
rect 22753 29597 22787 29631
rect 22787 29597 22796 29631
rect 22744 29588 22796 29597
rect 23112 29699 23164 29708
rect 23112 29665 23121 29699
rect 23121 29665 23155 29699
rect 23155 29665 23164 29699
rect 23112 29656 23164 29665
rect 22928 29631 22980 29640
rect 22928 29597 22937 29631
rect 22937 29597 22971 29631
rect 22971 29597 22980 29631
rect 22928 29588 22980 29597
rect 23572 29656 23624 29708
rect 20904 29452 20956 29504
rect 22468 29452 22520 29504
rect 22560 29495 22612 29504
rect 22560 29461 22569 29495
rect 22569 29461 22603 29495
rect 22603 29461 22612 29495
rect 22560 29452 22612 29461
rect 23112 29452 23164 29504
rect 23480 29588 23532 29640
rect 24584 29631 24636 29640
rect 24584 29597 24593 29631
rect 24593 29597 24627 29631
rect 24627 29597 24636 29631
rect 24584 29588 24636 29597
rect 24768 29588 24820 29640
rect 23572 29563 23624 29572
rect 23572 29529 23581 29563
rect 23581 29529 23615 29563
rect 23615 29529 23624 29563
rect 23572 29520 23624 29529
rect 23664 29563 23716 29572
rect 23664 29529 23673 29563
rect 23673 29529 23707 29563
rect 23707 29529 23716 29563
rect 23664 29520 23716 29529
rect 25228 29631 25280 29640
rect 25228 29597 25237 29631
rect 25237 29597 25271 29631
rect 25271 29597 25280 29631
rect 25228 29588 25280 29597
rect 27436 29656 27488 29708
rect 25136 29520 25188 29572
rect 26332 29520 26384 29572
rect 26516 29520 26568 29572
rect 26884 29563 26936 29572
rect 26884 29529 26893 29563
rect 26893 29529 26927 29563
rect 26927 29529 26936 29563
rect 26884 29520 26936 29529
rect 24124 29452 24176 29504
rect 24860 29452 24912 29504
rect 25688 29452 25740 29504
rect 26056 29452 26108 29504
rect 27252 29588 27304 29640
rect 27436 29520 27488 29572
rect 28448 29588 28500 29640
rect 28632 29588 28684 29640
rect 29552 29588 29604 29640
rect 30656 29656 30708 29708
rect 32220 29724 32272 29776
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 30288 29588 30340 29597
rect 30472 29631 30524 29640
rect 30472 29597 30481 29631
rect 30481 29597 30515 29631
rect 30515 29597 30524 29631
rect 30472 29588 30524 29597
rect 31116 29588 31168 29640
rect 31392 29631 31444 29640
rect 31392 29597 31401 29631
rect 31401 29597 31435 29631
rect 31435 29597 31444 29631
rect 31392 29588 31444 29597
rect 29092 29520 29144 29572
rect 30012 29520 30064 29572
rect 30564 29520 30616 29572
rect 30840 29520 30892 29572
rect 31300 29563 31352 29572
rect 31300 29529 31309 29563
rect 31309 29529 31343 29563
rect 31343 29529 31352 29563
rect 31300 29520 31352 29529
rect 32036 29520 32088 29572
rect 36268 29563 36320 29572
rect 36268 29529 36277 29563
rect 36277 29529 36311 29563
rect 36311 29529 36320 29563
rect 36268 29520 36320 29529
rect 30288 29452 30340 29504
rect 31484 29452 31536 29504
rect 31576 29495 31628 29504
rect 31576 29461 31585 29495
rect 31585 29461 31619 29495
rect 31619 29461 31628 29495
rect 31576 29452 31628 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1860 29223 1912 29232
rect 1860 29189 1869 29223
rect 1869 29189 1903 29223
rect 1903 29189 1912 29223
rect 1860 29180 1912 29189
rect 2688 29248 2740 29300
rect 3608 29291 3660 29300
rect 3608 29257 3617 29291
rect 3617 29257 3651 29291
rect 3651 29257 3660 29291
rect 3608 29248 3660 29257
rect 4068 29248 4120 29300
rect 4620 29248 4672 29300
rect 5080 29248 5132 29300
rect 5264 29248 5316 29300
rect 3332 29180 3384 29232
rect 2504 29044 2556 29096
rect 2596 29044 2648 29096
rect 1492 28976 1544 29028
rect 2320 28976 2372 29028
rect 3056 29155 3108 29164
rect 3056 29121 3065 29155
rect 3065 29121 3099 29155
rect 3099 29121 3108 29155
rect 3056 29112 3108 29121
rect 6644 29180 6696 29232
rect 3240 29044 3292 29096
rect 3424 29044 3476 29096
rect 4528 29155 4580 29164
rect 4528 29121 4537 29155
rect 4537 29121 4571 29155
rect 4571 29121 4580 29155
rect 4528 29112 4580 29121
rect 4712 29155 4764 29164
rect 4712 29121 4721 29155
rect 4721 29121 4755 29155
rect 4755 29121 4764 29155
rect 4712 29112 4764 29121
rect 4988 29155 5040 29164
rect 4988 29121 4997 29155
rect 4997 29121 5031 29155
rect 5031 29121 5040 29155
rect 4988 29112 5040 29121
rect 1768 28908 1820 28960
rect 2228 28951 2280 28960
rect 2228 28917 2237 28951
rect 2237 28917 2271 28951
rect 2271 28917 2280 28951
rect 2228 28908 2280 28917
rect 2412 28908 2464 28960
rect 3148 28976 3200 29028
rect 5448 29112 5500 29164
rect 7012 29248 7064 29300
rect 7012 29155 7064 29164
rect 7012 29121 7021 29155
rect 7021 29121 7055 29155
rect 7055 29121 7064 29155
rect 7012 29112 7064 29121
rect 7840 29248 7892 29300
rect 8116 29291 8168 29300
rect 8116 29257 8125 29291
rect 8125 29257 8159 29291
rect 8159 29257 8168 29291
rect 8116 29248 8168 29257
rect 9312 29248 9364 29300
rect 9496 29248 9548 29300
rect 7288 29112 7340 29164
rect 7564 29155 7616 29164
rect 7564 29121 7573 29155
rect 7573 29121 7607 29155
rect 7607 29121 7616 29155
rect 7564 29112 7616 29121
rect 8392 29180 8444 29232
rect 10324 29248 10376 29300
rect 11244 29248 11296 29300
rect 11612 29248 11664 29300
rect 12164 29248 12216 29300
rect 12532 29248 12584 29300
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 13084 29248 13136 29300
rect 16948 29248 17000 29300
rect 18144 29248 18196 29300
rect 18512 29291 18564 29300
rect 18512 29257 18521 29291
rect 18521 29257 18555 29291
rect 18555 29257 18564 29291
rect 18512 29248 18564 29257
rect 18880 29248 18932 29300
rect 19248 29248 19300 29300
rect 19616 29248 19668 29300
rect 8944 29044 8996 29096
rect 9220 29155 9272 29164
rect 9220 29121 9229 29155
rect 9229 29121 9263 29155
rect 9263 29121 9272 29155
rect 9220 29112 9272 29121
rect 9496 29155 9548 29164
rect 9496 29121 9524 29155
rect 9524 29121 9548 29155
rect 10416 29223 10468 29232
rect 10416 29189 10425 29223
rect 10425 29189 10459 29223
rect 10459 29189 10468 29223
rect 10416 29180 10468 29189
rect 10508 29180 10560 29232
rect 9496 29112 9548 29121
rect 9312 29087 9364 29096
rect 9312 29053 9321 29087
rect 9321 29053 9355 29087
rect 9355 29053 9364 29087
rect 9312 29044 9364 29053
rect 9772 29155 9824 29164
rect 9772 29121 9781 29155
rect 9781 29121 9815 29155
rect 9815 29121 9824 29155
rect 9772 29112 9824 29121
rect 10876 29155 10928 29164
rect 10876 29121 10885 29155
rect 10885 29121 10919 29155
rect 10919 29121 10928 29155
rect 10876 29112 10928 29121
rect 9128 28976 9180 29028
rect 2780 28908 2832 28960
rect 3332 28908 3384 28960
rect 3424 28951 3476 28960
rect 3424 28917 3433 28951
rect 3433 28917 3467 28951
rect 3467 28917 3476 28951
rect 3424 28908 3476 28917
rect 4804 28908 4856 28960
rect 5816 28908 5868 28960
rect 7012 28908 7064 28960
rect 8300 28908 8352 28960
rect 11336 29180 11388 29232
rect 11060 29155 11112 29164
rect 11060 29121 11069 29155
rect 11069 29121 11103 29155
rect 11103 29121 11112 29155
rect 11060 29112 11112 29121
rect 11152 29155 11204 29164
rect 11152 29121 11161 29155
rect 11161 29121 11195 29155
rect 11195 29121 11204 29155
rect 11152 29112 11204 29121
rect 11520 29112 11572 29164
rect 12900 29180 12952 29232
rect 11980 29112 12032 29164
rect 12808 29155 12860 29164
rect 12532 29087 12584 29096
rect 12532 29053 12541 29087
rect 12541 29053 12575 29087
rect 12575 29053 12584 29087
rect 12532 29044 12584 29053
rect 12808 29121 12814 29155
rect 12814 29121 12848 29155
rect 12848 29121 12860 29155
rect 12808 29112 12860 29121
rect 15936 29180 15988 29232
rect 13452 29112 13504 29164
rect 13636 29155 13688 29164
rect 13636 29121 13645 29155
rect 13645 29121 13679 29155
rect 13679 29121 13688 29155
rect 13636 29112 13688 29121
rect 13268 29087 13320 29096
rect 13268 29053 13277 29087
rect 13277 29053 13311 29087
rect 13311 29053 13320 29087
rect 13268 29044 13320 29053
rect 13728 29044 13780 29096
rect 10600 28908 10652 28960
rect 11060 28908 11112 28960
rect 11612 28908 11664 28960
rect 12072 28908 12124 28960
rect 12348 28951 12400 28960
rect 12348 28917 12357 28951
rect 12357 28917 12391 28951
rect 12391 28917 12400 28951
rect 12348 28908 12400 28917
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 14740 29112 14792 29164
rect 14924 29112 14976 29164
rect 15568 29112 15620 29164
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 17040 29223 17092 29232
rect 17040 29189 17049 29223
rect 17049 29189 17083 29223
rect 17083 29189 17092 29223
rect 17040 29180 17092 29189
rect 18420 29180 18472 29232
rect 20720 29248 20772 29300
rect 20812 29291 20864 29300
rect 20812 29257 20821 29291
rect 20821 29257 20855 29291
rect 20855 29257 20864 29291
rect 20812 29248 20864 29257
rect 20996 29248 21048 29300
rect 17408 29112 17460 29164
rect 17500 29112 17552 29164
rect 18144 29112 18196 29164
rect 14832 29044 14884 29096
rect 14740 28976 14792 29028
rect 15844 29087 15896 29096
rect 15844 29053 15853 29087
rect 15853 29053 15887 29087
rect 15887 29053 15896 29087
rect 15844 29044 15896 29053
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 17776 29044 17828 29096
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 19340 29044 19392 29096
rect 19984 29112 20036 29164
rect 19616 29044 19668 29096
rect 20536 29112 20588 29164
rect 21180 29248 21232 29300
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 21180 29112 21232 29121
rect 22744 29248 22796 29300
rect 23664 29248 23716 29300
rect 23756 29248 23808 29300
rect 23848 29248 23900 29300
rect 24400 29248 24452 29300
rect 23296 29180 23348 29232
rect 21456 29155 21508 29164
rect 21456 29121 21475 29155
rect 21475 29121 21508 29155
rect 21456 29112 21508 29121
rect 21732 29112 21784 29164
rect 22744 29112 22796 29164
rect 23020 29155 23072 29164
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23204 29155 23256 29164
rect 23204 29121 23213 29155
rect 23213 29121 23247 29155
rect 23247 29121 23256 29155
rect 23204 29112 23256 29121
rect 23664 29155 23716 29164
rect 23664 29121 23673 29155
rect 23673 29121 23707 29155
rect 23707 29121 23716 29155
rect 23664 29112 23716 29121
rect 22928 29087 22980 29096
rect 22928 29053 22937 29087
rect 22937 29053 22971 29087
rect 22971 29053 22980 29087
rect 22928 29044 22980 29053
rect 24216 29180 24268 29232
rect 24308 29112 24360 29164
rect 24952 29180 25004 29232
rect 25228 29248 25280 29300
rect 25504 29248 25556 29300
rect 26976 29291 27028 29300
rect 26976 29257 26985 29291
rect 26985 29257 27019 29291
rect 27019 29257 27028 29291
rect 26976 29248 27028 29257
rect 24584 29155 24636 29164
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 24676 29155 24728 29164
rect 24676 29121 24685 29155
rect 24685 29121 24719 29155
rect 24719 29121 24728 29155
rect 24676 29112 24728 29121
rect 25044 29155 25096 29164
rect 25044 29121 25053 29155
rect 25053 29121 25087 29155
rect 25087 29121 25096 29155
rect 27068 29180 27120 29232
rect 25044 29112 25096 29121
rect 24768 29044 24820 29096
rect 25412 29155 25464 29164
rect 25412 29121 25422 29155
rect 25422 29121 25456 29155
rect 25456 29121 25464 29155
rect 25412 29112 25464 29121
rect 25688 29112 25740 29164
rect 26424 29112 26476 29164
rect 27528 29248 27580 29300
rect 27712 29248 27764 29300
rect 28724 29248 28776 29300
rect 27436 29180 27488 29232
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27528 29112 27580 29164
rect 27896 29180 27948 29232
rect 26240 29044 26292 29096
rect 28540 29180 28592 29232
rect 29092 29248 29144 29300
rect 29184 29248 29236 29300
rect 29092 29112 29144 29164
rect 29368 29155 29420 29164
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 29460 29155 29512 29164
rect 29460 29121 29469 29155
rect 29469 29121 29503 29155
rect 29503 29121 29512 29155
rect 29460 29112 29512 29121
rect 29552 29112 29604 29164
rect 30380 29248 30432 29300
rect 31576 29248 31628 29300
rect 33232 29248 33284 29300
rect 30840 29223 30892 29232
rect 30840 29189 30849 29223
rect 30849 29189 30883 29223
rect 30883 29189 30892 29223
rect 30840 29180 30892 29189
rect 12532 28908 12584 28960
rect 12992 28908 13044 28960
rect 13452 28951 13504 28960
rect 13452 28917 13461 28951
rect 13461 28917 13495 28951
rect 13495 28917 13504 28951
rect 13452 28908 13504 28917
rect 13544 28908 13596 28960
rect 17684 28908 17736 28960
rect 19064 28908 19116 28960
rect 19156 28908 19208 28960
rect 20536 28908 20588 28960
rect 22652 28908 22704 28960
rect 24400 28908 24452 28960
rect 27896 28976 27948 29028
rect 28080 28976 28132 29028
rect 28540 29019 28592 29028
rect 28540 28985 28549 29019
rect 28549 28985 28583 29019
rect 28583 28985 28592 29019
rect 28540 28976 28592 28985
rect 28632 28976 28684 29028
rect 29276 29044 29328 29096
rect 30288 29155 30340 29164
rect 30288 29121 30297 29155
rect 30297 29121 30331 29155
rect 30331 29121 30340 29155
rect 30288 29112 30340 29121
rect 30564 29112 30616 29164
rect 31024 29155 31076 29164
rect 31024 29121 31033 29155
rect 31033 29121 31067 29155
rect 31067 29121 31076 29155
rect 31024 29112 31076 29121
rect 31116 29112 31168 29164
rect 30104 29087 30156 29096
rect 30104 29053 30113 29087
rect 30113 29053 30147 29087
rect 30147 29053 30156 29087
rect 30104 29044 30156 29053
rect 31392 29112 31444 29164
rect 31668 29180 31720 29232
rect 33416 29112 33468 29164
rect 29644 28976 29696 29028
rect 30656 28976 30708 29028
rect 33048 29044 33100 29096
rect 33692 28976 33744 29028
rect 34060 28976 34112 29028
rect 28908 28908 28960 28960
rect 30564 28908 30616 28960
rect 33508 28908 33560 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2504 28704 2556 28756
rect 3424 28704 3476 28756
rect 3700 28704 3752 28756
rect 3976 28747 4028 28756
rect 3976 28713 3985 28747
rect 3985 28713 4019 28747
rect 4019 28713 4028 28747
rect 3976 28704 4028 28713
rect 5080 28704 5132 28756
rect 5448 28704 5500 28756
rect 5632 28704 5684 28756
rect 7196 28704 7248 28756
rect 7840 28747 7892 28756
rect 7840 28713 7849 28747
rect 7849 28713 7883 28747
rect 7883 28713 7892 28747
rect 7840 28704 7892 28713
rect 9312 28704 9364 28756
rect 9956 28747 10008 28756
rect 9956 28713 9965 28747
rect 9965 28713 9999 28747
rect 9999 28713 10008 28747
rect 9956 28704 10008 28713
rect 10324 28704 10376 28756
rect 11152 28704 11204 28756
rect 11520 28704 11572 28756
rect 11980 28704 12032 28756
rect 12348 28704 12400 28756
rect 12716 28704 12768 28756
rect 13268 28704 13320 28756
rect 13360 28747 13412 28756
rect 13360 28713 13369 28747
rect 13369 28713 13403 28747
rect 13403 28713 13412 28747
rect 13360 28704 13412 28713
rect 14188 28704 14240 28756
rect 14832 28704 14884 28756
rect 17316 28704 17368 28756
rect 1216 28568 1268 28620
rect 3792 28568 3844 28620
rect 4344 28568 4396 28620
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 2596 28500 2648 28552
rect 3056 28543 3108 28552
rect 3056 28509 3065 28543
rect 3065 28509 3099 28543
rect 3099 28509 3108 28543
rect 3056 28500 3108 28509
rect 1860 28364 1912 28416
rect 3240 28407 3292 28416
rect 3240 28373 3249 28407
rect 3249 28373 3283 28407
rect 3283 28373 3292 28407
rect 3240 28364 3292 28373
rect 3424 28432 3476 28484
rect 3792 28475 3844 28484
rect 3792 28441 3801 28475
rect 3801 28441 3835 28475
rect 3835 28441 3844 28475
rect 3792 28432 3844 28441
rect 4436 28475 4488 28484
rect 4436 28441 4445 28475
rect 4445 28441 4479 28475
rect 4479 28441 4488 28475
rect 4436 28432 4488 28441
rect 4896 28432 4948 28484
rect 5264 28475 5316 28484
rect 5264 28441 5273 28475
rect 5273 28441 5307 28475
rect 5307 28441 5316 28475
rect 5264 28432 5316 28441
rect 5448 28543 5500 28552
rect 5448 28509 5457 28543
rect 5457 28509 5491 28543
rect 5491 28509 5500 28543
rect 5448 28500 5500 28509
rect 5540 28543 5592 28552
rect 5540 28509 5549 28543
rect 5549 28509 5583 28543
rect 5583 28509 5592 28543
rect 5816 28636 5868 28688
rect 6368 28568 6420 28620
rect 6552 28568 6604 28620
rect 6736 28568 6788 28620
rect 5540 28500 5592 28509
rect 5816 28500 5868 28552
rect 10508 28636 10560 28688
rect 8300 28611 8352 28620
rect 8300 28577 8309 28611
rect 8309 28577 8343 28611
rect 8343 28577 8352 28611
rect 8300 28568 8352 28577
rect 8668 28568 8720 28620
rect 9588 28568 9640 28620
rect 12164 28568 12216 28620
rect 6092 28432 6144 28484
rect 6736 28432 6788 28484
rect 7196 28432 7248 28484
rect 4160 28407 4212 28416
rect 4160 28373 4169 28407
rect 4169 28373 4203 28407
rect 4203 28373 4212 28407
rect 4160 28364 4212 28373
rect 4988 28364 5040 28416
rect 5080 28364 5132 28416
rect 5172 28407 5224 28416
rect 5172 28373 5181 28407
rect 5181 28373 5215 28407
rect 5215 28373 5224 28407
rect 5172 28364 5224 28373
rect 5356 28407 5408 28416
rect 5356 28373 5371 28407
rect 5371 28373 5405 28407
rect 5405 28373 5408 28407
rect 5356 28364 5408 28373
rect 5632 28364 5684 28416
rect 7564 28364 7616 28416
rect 9220 28500 9272 28552
rect 8944 28432 8996 28484
rect 9680 28432 9732 28484
rect 10784 28500 10836 28552
rect 15844 28636 15896 28688
rect 12624 28568 12676 28620
rect 13452 28611 13504 28620
rect 13452 28577 13461 28611
rect 13461 28577 13495 28611
rect 13495 28577 13504 28611
rect 13452 28568 13504 28577
rect 11244 28432 11296 28484
rect 11888 28432 11940 28484
rect 12532 28432 12584 28484
rect 11612 28364 11664 28416
rect 11796 28407 11848 28416
rect 11796 28373 11805 28407
rect 11805 28373 11839 28407
rect 11839 28373 11848 28407
rect 11796 28364 11848 28373
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 13452 28432 13504 28484
rect 13728 28543 13780 28552
rect 13728 28509 13737 28543
rect 13737 28509 13771 28543
rect 13771 28509 13780 28543
rect 13728 28500 13780 28509
rect 16764 28500 16816 28552
rect 17316 28500 17368 28552
rect 17960 28704 18012 28756
rect 17868 28636 17920 28688
rect 20168 28704 20220 28756
rect 18604 28636 18656 28688
rect 18972 28636 19024 28688
rect 19800 28679 19852 28688
rect 19800 28645 19809 28679
rect 19809 28645 19843 28679
rect 19843 28645 19852 28679
rect 19800 28636 19852 28645
rect 19892 28636 19944 28688
rect 23204 28747 23256 28756
rect 23204 28713 23213 28747
rect 23213 28713 23247 28747
rect 23247 28713 23256 28747
rect 23204 28704 23256 28713
rect 23664 28704 23716 28756
rect 24124 28704 24176 28756
rect 24400 28704 24452 28756
rect 26424 28747 26476 28756
rect 26424 28713 26433 28747
rect 26433 28713 26467 28747
rect 26467 28713 26476 28747
rect 26424 28704 26476 28713
rect 26884 28704 26936 28756
rect 27160 28704 27212 28756
rect 27528 28704 27580 28756
rect 14372 28432 14424 28484
rect 16488 28432 16540 28484
rect 18604 28500 18656 28552
rect 18972 28500 19024 28552
rect 19064 28500 19116 28552
rect 19156 28500 19208 28552
rect 20812 28568 20864 28620
rect 14096 28364 14148 28416
rect 15292 28364 15344 28416
rect 15936 28407 15988 28416
rect 15936 28373 15945 28407
rect 15945 28373 15979 28407
rect 15979 28373 15988 28407
rect 15936 28364 15988 28373
rect 16948 28364 17000 28416
rect 17500 28364 17552 28416
rect 18144 28432 18196 28484
rect 20076 28543 20128 28552
rect 20076 28509 20085 28543
rect 20085 28509 20119 28543
rect 20119 28509 20128 28543
rect 20076 28500 20128 28509
rect 20168 28543 20220 28552
rect 20168 28509 20177 28543
rect 20177 28509 20211 28543
rect 20211 28509 20220 28543
rect 20168 28500 20220 28509
rect 20352 28500 20404 28552
rect 26608 28636 26660 28688
rect 27344 28636 27396 28688
rect 26240 28568 26292 28620
rect 26884 28611 26936 28620
rect 26884 28577 26893 28611
rect 26893 28577 26927 28611
rect 26927 28577 26936 28611
rect 26884 28568 26936 28577
rect 19156 28364 19208 28416
rect 19423 28364 19475 28416
rect 20444 28407 20496 28416
rect 20444 28373 20453 28407
rect 20453 28373 20487 28407
rect 20487 28373 20496 28407
rect 20444 28364 20496 28373
rect 20904 28364 20956 28416
rect 25688 28432 25740 28484
rect 26700 28500 26752 28552
rect 27436 28568 27488 28620
rect 28724 28704 28776 28756
rect 28816 28704 28868 28756
rect 28264 28636 28316 28688
rect 29000 28636 29052 28688
rect 31116 28704 31168 28756
rect 32956 28704 33008 28756
rect 33416 28747 33468 28756
rect 33416 28713 33425 28747
rect 33425 28713 33459 28747
rect 33459 28713 33468 28747
rect 33416 28704 33468 28713
rect 43536 28704 43588 28756
rect 42156 28679 42208 28688
rect 42156 28645 42165 28679
rect 42165 28645 42199 28679
rect 42199 28645 42208 28679
rect 42156 28636 42208 28645
rect 28540 28568 28592 28620
rect 29184 28568 29236 28620
rect 29736 28568 29788 28620
rect 26240 28475 26292 28484
rect 26240 28441 26249 28475
rect 26249 28441 26283 28475
rect 26283 28441 26292 28475
rect 26240 28432 26292 28441
rect 26332 28432 26384 28484
rect 27712 28500 27764 28552
rect 28264 28432 28316 28484
rect 28724 28543 28776 28552
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 28724 28500 28776 28509
rect 29092 28500 29144 28552
rect 32036 28611 32088 28620
rect 32036 28577 32045 28611
rect 32045 28577 32079 28611
rect 32079 28577 32088 28611
rect 32036 28568 32088 28577
rect 33048 28568 33100 28620
rect 30288 28500 30340 28552
rect 31024 28500 31076 28552
rect 28540 28432 28592 28484
rect 30380 28432 30432 28484
rect 30748 28475 30800 28484
rect 30748 28441 30757 28475
rect 30757 28441 30791 28475
rect 30791 28441 30800 28475
rect 30748 28432 30800 28441
rect 31392 28543 31444 28552
rect 31392 28509 31401 28543
rect 31401 28509 31435 28543
rect 31435 28509 31444 28543
rect 31392 28500 31444 28509
rect 33508 28543 33560 28552
rect 33508 28509 33517 28543
rect 33517 28509 33551 28543
rect 33551 28509 33560 28543
rect 33508 28500 33560 28509
rect 41880 28500 41932 28552
rect 42340 28543 42392 28552
rect 42340 28509 42349 28543
rect 42349 28509 42383 28543
rect 42383 28509 42392 28543
rect 42340 28500 42392 28509
rect 42800 28500 42852 28552
rect 32128 28432 32180 28484
rect 33968 28432 34020 28484
rect 36268 28432 36320 28484
rect 42984 28432 43036 28484
rect 21916 28364 21968 28416
rect 24308 28364 24360 28416
rect 25044 28407 25096 28416
rect 25044 28373 25053 28407
rect 25053 28373 25087 28407
rect 25087 28373 25096 28407
rect 25044 28364 25096 28373
rect 26148 28407 26200 28416
rect 26148 28373 26157 28407
rect 26157 28373 26191 28407
rect 26191 28373 26200 28407
rect 26148 28364 26200 28373
rect 26424 28407 26476 28416
rect 26424 28373 26449 28407
rect 26449 28373 26476 28407
rect 26424 28364 26476 28373
rect 26608 28407 26660 28416
rect 26608 28373 26617 28407
rect 26617 28373 26651 28407
rect 26651 28373 26660 28407
rect 26608 28364 26660 28373
rect 27252 28364 27304 28416
rect 27528 28364 27580 28416
rect 28632 28364 28684 28416
rect 33232 28364 33284 28416
rect 33508 28364 33560 28416
rect 41880 28407 41932 28416
rect 41880 28373 41889 28407
rect 41889 28373 41923 28407
rect 41923 28373 41932 28407
rect 41880 28364 41932 28373
rect 43260 28364 43312 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 1768 28160 1820 28212
rect 1860 28203 1912 28212
rect 1860 28169 1869 28203
rect 1869 28169 1903 28203
rect 1903 28169 1912 28203
rect 1860 28160 1912 28169
rect 2412 28160 2464 28212
rect 3792 28160 3844 28212
rect 4068 28160 4120 28212
rect 4344 28203 4396 28212
rect 4344 28169 4353 28203
rect 4353 28169 4387 28203
rect 4387 28169 4396 28203
rect 4344 28160 4396 28169
rect 4712 28160 4764 28212
rect 5172 28160 5224 28212
rect 5448 28160 5500 28212
rect 6736 28160 6788 28212
rect 9128 28160 9180 28212
rect 9220 28160 9272 28212
rect 10600 28203 10652 28212
rect 10600 28169 10609 28203
rect 10609 28169 10643 28203
rect 10643 28169 10652 28203
rect 10600 28160 10652 28169
rect 10784 28160 10836 28212
rect 12992 28160 13044 28212
rect 13084 28160 13136 28212
rect 13176 28160 13228 28212
rect 3056 28135 3108 28144
rect 3056 28101 3065 28135
rect 3065 28101 3099 28135
rect 3099 28101 3108 28135
rect 3056 28092 3108 28101
rect 1860 28024 1912 28076
rect 3240 28092 3292 28144
rect 3516 28067 3568 28076
rect 3516 28033 3525 28067
rect 3525 28033 3559 28067
rect 3559 28033 3568 28067
rect 3516 28024 3568 28033
rect 2136 27956 2188 28008
rect 2504 27999 2556 28008
rect 2504 27965 2513 27999
rect 2513 27965 2547 27999
rect 2547 27965 2556 27999
rect 2504 27956 2556 27965
rect 3884 27888 3936 27940
rect 4528 27888 4580 27940
rect 4620 27888 4672 27940
rect 4804 27956 4856 28008
rect 5356 28024 5408 28076
rect 5632 28024 5684 28076
rect 6092 28092 6144 28144
rect 5540 27956 5592 28008
rect 7104 28092 7156 28144
rect 6644 28067 6696 28076
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 6828 28024 6880 28076
rect 7196 28024 7248 28076
rect 8300 28024 8352 28076
rect 10508 28135 10560 28144
rect 10508 28101 10517 28135
rect 10517 28101 10551 28135
rect 10551 28101 10560 28135
rect 10508 28092 10560 28101
rect 6184 27888 6236 27940
rect 2688 27863 2740 27872
rect 2688 27829 2697 27863
rect 2697 27829 2731 27863
rect 2731 27829 2740 27863
rect 2688 27820 2740 27829
rect 3148 27820 3200 27872
rect 5264 27820 5316 27872
rect 5448 27820 5500 27872
rect 8024 27956 8076 28008
rect 9312 27956 9364 28008
rect 8208 27888 8260 27940
rect 6828 27820 6880 27872
rect 7564 27820 7616 27872
rect 7932 27820 7984 27872
rect 8760 27863 8812 27872
rect 8760 27829 8769 27863
rect 8769 27829 8803 27863
rect 8803 27829 8812 27863
rect 8760 27820 8812 27829
rect 8944 27888 8996 27940
rect 9496 27888 9548 27940
rect 9864 28067 9916 28076
rect 9864 28033 9873 28067
rect 9873 28033 9907 28067
rect 9907 28033 9916 28067
rect 9864 28024 9916 28033
rect 10324 27956 10376 28008
rect 10416 27956 10468 28008
rect 11060 27999 11112 28008
rect 11060 27965 11069 27999
rect 11069 27965 11103 27999
rect 11103 27965 11112 27999
rect 11060 27956 11112 27965
rect 11244 28092 11296 28144
rect 11336 28024 11388 28076
rect 11888 28092 11940 28144
rect 13360 28160 13412 28212
rect 13820 28160 13872 28212
rect 14188 28160 14240 28212
rect 15016 28203 15068 28212
rect 15016 28169 15025 28203
rect 15025 28169 15059 28203
rect 15059 28169 15068 28203
rect 15016 28160 15068 28169
rect 15384 28160 15436 28212
rect 15936 28160 15988 28212
rect 16764 28160 16816 28212
rect 13084 28067 13136 28076
rect 13084 28033 13112 28067
rect 13112 28033 13136 28067
rect 13084 28024 13136 28033
rect 12072 27956 12124 28008
rect 12992 27956 13044 28008
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 13728 28092 13780 28144
rect 15292 28092 15344 28144
rect 16396 28092 16448 28144
rect 13820 28067 13872 28076
rect 13820 28033 13829 28067
rect 13829 28033 13863 28067
rect 13863 28033 13872 28067
rect 13820 28024 13872 28033
rect 16488 28024 16540 28076
rect 9680 27888 9732 27940
rect 10232 27888 10284 27940
rect 11612 27931 11664 27940
rect 11612 27897 11621 27931
rect 11621 27897 11655 27931
rect 11655 27897 11664 27931
rect 11612 27888 11664 27897
rect 12348 27888 12400 27940
rect 12440 27888 12492 27940
rect 14188 27956 14240 28008
rect 14648 27956 14700 28008
rect 15568 27999 15620 28008
rect 15568 27965 15577 27999
rect 15577 27965 15611 27999
rect 15611 27965 15620 27999
rect 15568 27956 15620 27965
rect 16764 27956 16816 28008
rect 18420 28092 18472 28144
rect 17592 28067 17644 28076
rect 17592 28033 17601 28067
rect 17601 28033 17635 28067
rect 17635 28033 17644 28067
rect 17592 28024 17644 28033
rect 17684 27956 17736 28008
rect 19340 28024 19392 28076
rect 19800 28092 19852 28144
rect 24308 28203 24360 28212
rect 24308 28169 24317 28203
rect 24317 28169 24351 28203
rect 24351 28169 24360 28203
rect 24308 28160 24360 28169
rect 24400 28160 24452 28212
rect 26240 28160 26292 28212
rect 27712 28160 27764 28212
rect 20444 28024 20496 28076
rect 20904 28092 20956 28144
rect 13636 27888 13688 27940
rect 15200 27888 15252 27940
rect 12164 27820 12216 27872
rect 13544 27820 13596 27872
rect 14372 27863 14424 27872
rect 14372 27829 14381 27863
rect 14381 27829 14415 27863
rect 14415 27829 14424 27863
rect 14372 27820 14424 27829
rect 15016 27820 15068 27872
rect 16212 27863 16264 27872
rect 16212 27829 16221 27863
rect 16221 27829 16255 27863
rect 16255 27829 16264 27863
rect 16212 27820 16264 27829
rect 17040 27888 17092 27940
rect 17592 27820 17644 27872
rect 17776 27820 17828 27872
rect 18972 27956 19024 28008
rect 21916 28067 21968 28076
rect 21916 28033 21925 28067
rect 21925 28033 21959 28067
rect 21959 28033 21968 28067
rect 21916 28024 21968 28033
rect 22468 28024 22520 28076
rect 22652 28024 22704 28076
rect 27804 28092 27856 28144
rect 30748 28160 30800 28212
rect 32128 28160 32180 28212
rect 33968 28203 34020 28212
rect 33968 28169 33977 28203
rect 33977 28169 34011 28203
rect 34011 28169 34020 28203
rect 33968 28160 34020 28169
rect 25044 28024 25096 28076
rect 25872 28024 25924 28076
rect 26792 28024 26844 28076
rect 27252 28024 27304 28076
rect 27528 28024 27580 28076
rect 27620 28067 27672 28076
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 27712 28067 27764 28076
rect 27712 28033 27721 28067
rect 27721 28033 27755 28067
rect 27755 28033 27764 28067
rect 27712 28024 27764 28033
rect 28080 28024 28132 28076
rect 28632 28024 28684 28076
rect 29276 28092 29328 28144
rect 18420 27820 18472 27872
rect 20720 27820 20772 27872
rect 20812 27820 20864 27872
rect 21088 27863 21140 27872
rect 21088 27829 21097 27863
rect 21097 27829 21131 27863
rect 21131 27829 21140 27863
rect 21088 27820 21140 27829
rect 21272 27820 21324 27872
rect 26240 27888 26292 27940
rect 23664 27820 23716 27872
rect 25688 27820 25740 27872
rect 26332 27820 26384 27872
rect 26700 27820 26752 27872
rect 27068 27820 27120 27872
rect 27344 27888 27396 27940
rect 27528 27888 27580 27940
rect 30656 28024 30708 28076
rect 28356 27888 28408 27940
rect 28540 27888 28592 27940
rect 30380 27956 30432 28008
rect 30104 27863 30156 27872
rect 30104 27829 30113 27863
rect 30113 27829 30147 27863
rect 30147 27829 30156 27863
rect 30104 27820 30156 27829
rect 30196 27820 30248 27872
rect 32128 28067 32180 28076
rect 32128 28033 32137 28067
rect 32137 28033 32171 28067
rect 32171 28033 32180 28067
rect 32128 28024 32180 28033
rect 33508 28024 33560 28076
rect 33600 28067 33652 28076
rect 33600 28033 33609 28067
rect 33609 28033 33643 28067
rect 33643 28033 33652 28067
rect 33600 28024 33652 28033
rect 33692 28024 33744 28076
rect 36268 28024 36320 28076
rect 41880 28160 41932 28212
rect 42340 28160 42392 28212
rect 42800 28092 42852 28144
rect 42984 28135 43036 28144
rect 42984 28101 43002 28135
rect 43002 28101 43036 28135
rect 42984 28092 43036 28101
rect 43812 28024 43864 28076
rect 43260 27820 43312 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3792 27616 3844 27668
rect 4160 27616 4212 27668
rect 2044 27548 2096 27600
rect 3332 27548 3384 27600
rect 5080 27616 5132 27668
rect 1216 27480 1268 27532
rect 3148 27412 3200 27464
rect 4344 27480 4396 27532
rect 5356 27548 5408 27600
rect 5632 27616 5684 27668
rect 6184 27548 6236 27600
rect 6368 27591 6420 27600
rect 6368 27557 6377 27591
rect 6377 27557 6411 27591
rect 6411 27557 6420 27591
rect 6368 27548 6420 27557
rect 7104 27659 7156 27668
rect 7104 27625 7113 27659
rect 7113 27625 7147 27659
rect 7147 27625 7156 27659
rect 7104 27616 7156 27625
rect 8300 27616 8352 27668
rect 8760 27616 8812 27668
rect 9864 27616 9916 27668
rect 10324 27659 10376 27668
rect 10324 27625 10333 27659
rect 10333 27625 10367 27659
rect 10367 27625 10376 27659
rect 10324 27616 10376 27625
rect 11152 27616 11204 27668
rect 11796 27616 11848 27668
rect 12348 27616 12400 27668
rect 13176 27616 13228 27668
rect 16948 27616 17000 27668
rect 17960 27616 18012 27668
rect 18972 27659 19024 27668
rect 18972 27625 18981 27659
rect 18981 27625 19015 27659
rect 19015 27625 19024 27659
rect 18972 27616 19024 27625
rect 19340 27616 19392 27668
rect 20076 27616 20128 27668
rect 20352 27616 20404 27668
rect 21732 27616 21784 27668
rect 3700 27412 3752 27464
rect 3884 27412 3936 27464
rect 4712 27412 4764 27464
rect 4988 27455 5040 27464
rect 4988 27421 4997 27455
rect 4997 27421 5031 27455
rect 5031 27421 5040 27455
rect 4988 27412 5040 27421
rect 4344 27387 4396 27396
rect 4344 27353 4353 27387
rect 4353 27353 4387 27387
rect 4387 27353 4396 27387
rect 4344 27344 4396 27353
rect 4436 27344 4488 27396
rect 1584 27276 1636 27328
rect 2504 27276 2556 27328
rect 4252 27276 4304 27328
rect 4804 27344 4856 27396
rect 5264 27412 5316 27464
rect 5632 27412 5684 27464
rect 5540 27344 5592 27396
rect 7288 27412 7340 27464
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 7564 27412 7616 27421
rect 8208 27548 8260 27600
rect 8392 27591 8444 27600
rect 8392 27557 8401 27591
rect 8401 27557 8435 27591
rect 8435 27557 8444 27591
rect 8392 27548 8444 27557
rect 9220 27548 9272 27600
rect 7932 27412 7984 27464
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 5632 27319 5684 27328
rect 5632 27285 5641 27319
rect 5641 27285 5675 27319
rect 5675 27285 5684 27319
rect 5632 27276 5684 27285
rect 6000 27319 6052 27328
rect 6000 27285 6009 27319
rect 6009 27285 6043 27319
rect 6043 27285 6052 27319
rect 6000 27276 6052 27285
rect 6092 27276 6144 27328
rect 6828 27276 6880 27328
rect 7196 27276 7248 27328
rect 7748 27276 7800 27328
rect 8576 27455 8628 27464
rect 8576 27421 8585 27455
rect 8585 27421 8619 27455
rect 8619 27421 8628 27455
rect 8576 27412 8628 27421
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 9220 27412 9272 27421
rect 9220 27276 9272 27328
rect 9588 27412 9640 27464
rect 10232 27523 10284 27532
rect 10232 27489 10241 27523
rect 10241 27489 10275 27523
rect 10275 27489 10284 27523
rect 10232 27480 10284 27489
rect 10140 27455 10192 27464
rect 10140 27421 10149 27455
rect 10149 27421 10183 27455
rect 10183 27421 10192 27455
rect 10140 27412 10192 27421
rect 12164 27548 12216 27600
rect 12808 27548 12860 27600
rect 12900 27548 12952 27600
rect 13728 27591 13780 27600
rect 13728 27557 13737 27591
rect 13737 27557 13771 27591
rect 13771 27557 13780 27591
rect 13728 27548 13780 27557
rect 15016 27591 15068 27600
rect 10416 27344 10468 27396
rect 10692 27344 10744 27396
rect 9680 27276 9732 27328
rect 11060 27412 11112 27464
rect 11244 27412 11296 27464
rect 15016 27557 15025 27591
rect 15025 27557 15059 27591
rect 15059 27557 15068 27591
rect 15016 27548 15068 27557
rect 20996 27548 21048 27600
rect 21180 27548 21232 27600
rect 14004 27480 14056 27532
rect 19432 27480 19484 27532
rect 20720 27480 20772 27532
rect 23388 27548 23440 27600
rect 24492 27548 24544 27600
rect 23572 27480 23624 27532
rect 12624 27455 12676 27464
rect 12624 27421 12633 27455
rect 12633 27421 12667 27455
rect 12667 27421 12676 27455
rect 12624 27412 12676 27421
rect 13176 27455 13228 27464
rect 13176 27421 13185 27455
rect 13185 27421 13219 27455
rect 13219 27421 13228 27455
rect 13176 27412 13228 27421
rect 13268 27412 13320 27464
rect 14280 27412 14332 27464
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 14740 27344 14792 27396
rect 14924 27412 14976 27464
rect 17224 27455 17276 27464
rect 17224 27421 17233 27455
rect 17233 27421 17267 27455
rect 17267 27421 17276 27455
rect 17224 27412 17276 27421
rect 17868 27412 17920 27464
rect 11336 27276 11388 27328
rect 11428 27276 11480 27328
rect 13268 27276 13320 27328
rect 15292 27276 15344 27328
rect 16212 27344 16264 27396
rect 18052 27344 18104 27396
rect 20076 27455 20128 27464
rect 20076 27421 20085 27455
rect 20085 27421 20119 27455
rect 20119 27421 20128 27455
rect 20076 27412 20128 27421
rect 21088 27412 21140 27464
rect 21272 27412 21324 27464
rect 23756 27412 23808 27464
rect 22192 27387 22244 27396
rect 22192 27353 22201 27387
rect 22201 27353 22235 27387
rect 22235 27353 22244 27387
rect 22192 27344 22244 27353
rect 22928 27344 22980 27396
rect 24032 27412 24084 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 26332 27548 26384 27600
rect 27344 27616 27396 27668
rect 28080 27616 28132 27668
rect 28724 27659 28776 27668
rect 28724 27625 28733 27659
rect 28733 27625 28767 27659
rect 28767 27625 28776 27659
rect 28724 27616 28776 27625
rect 25320 27480 25372 27532
rect 25596 27412 25648 27464
rect 26056 27412 26108 27464
rect 17408 27276 17460 27328
rect 19248 27319 19300 27328
rect 19248 27285 19257 27319
rect 19257 27285 19291 27319
rect 19291 27285 19300 27319
rect 19248 27276 19300 27285
rect 19432 27276 19484 27328
rect 20720 27319 20772 27328
rect 20720 27285 20729 27319
rect 20729 27285 20763 27319
rect 20763 27285 20772 27319
rect 20720 27276 20772 27285
rect 21640 27276 21692 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 25596 27276 25648 27328
rect 26056 27319 26108 27328
rect 26056 27285 26065 27319
rect 26065 27285 26099 27319
rect 26099 27285 26108 27319
rect 26056 27276 26108 27285
rect 26424 27480 26476 27532
rect 26516 27412 26568 27464
rect 26792 27455 26844 27464
rect 26792 27421 26801 27455
rect 26801 27421 26835 27455
rect 26835 27421 26844 27455
rect 26792 27412 26844 27421
rect 28724 27480 28776 27532
rect 26424 27387 26476 27396
rect 26424 27353 26433 27387
rect 26433 27353 26467 27387
rect 26467 27353 26476 27387
rect 26424 27344 26476 27353
rect 27344 27455 27396 27464
rect 27344 27421 27353 27455
rect 27353 27421 27387 27455
rect 27387 27421 27396 27455
rect 27344 27412 27396 27421
rect 27252 27344 27304 27396
rect 27528 27412 27580 27464
rect 28080 27412 28132 27464
rect 28172 27412 28224 27464
rect 29828 27548 29880 27600
rect 30196 27616 30248 27668
rect 31024 27616 31076 27668
rect 30564 27548 30616 27600
rect 29000 27455 29052 27464
rect 29000 27421 29009 27455
rect 29009 27421 29043 27455
rect 29043 27421 29052 27455
rect 29000 27412 29052 27421
rect 30288 27455 30340 27464
rect 30288 27421 30297 27455
rect 30297 27421 30331 27455
rect 30331 27421 30340 27455
rect 30288 27412 30340 27421
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30748 27412 30800 27464
rect 30932 27455 30984 27464
rect 30932 27421 30941 27455
rect 30941 27421 30975 27455
rect 30975 27421 30984 27455
rect 30932 27412 30984 27421
rect 31208 27616 31260 27668
rect 34060 27659 34112 27668
rect 34060 27625 34069 27659
rect 34069 27625 34103 27659
rect 34103 27625 34112 27659
rect 34060 27616 34112 27625
rect 31760 27548 31812 27600
rect 33048 27548 33100 27600
rect 27160 27319 27212 27328
rect 27160 27285 27169 27319
rect 27169 27285 27203 27319
rect 27203 27285 27212 27319
rect 27160 27276 27212 27285
rect 27896 27344 27948 27396
rect 29368 27344 29420 27396
rect 29828 27344 29880 27396
rect 31484 27412 31536 27464
rect 31944 27455 31996 27464
rect 31944 27421 31953 27455
rect 31953 27421 31987 27455
rect 31987 27421 31996 27455
rect 31944 27412 31996 27421
rect 32680 27412 32732 27464
rect 33232 27480 33284 27532
rect 28172 27319 28224 27328
rect 28172 27285 28181 27319
rect 28181 27285 28215 27319
rect 28215 27285 28224 27319
rect 28172 27276 28224 27285
rect 29736 27319 29788 27328
rect 29736 27285 29745 27319
rect 29745 27285 29779 27319
rect 29779 27285 29788 27319
rect 29736 27276 29788 27285
rect 31024 27276 31076 27328
rect 32220 27276 32272 27328
rect 32588 27344 32640 27396
rect 32956 27387 33008 27396
rect 32956 27353 32965 27387
rect 32965 27353 32999 27387
rect 32999 27353 33008 27387
rect 32956 27344 33008 27353
rect 34060 27344 34112 27396
rect 33784 27319 33836 27328
rect 33784 27285 33793 27319
rect 33793 27285 33827 27319
rect 33827 27285 33836 27319
rect 33784 27276 33836 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2872 27072 2924 27124
rect 3424 27115 3476 27124
rect 3424 27081 3433 27115
rect 3433 27081 3467 27115
rect 3467 27081 3476 27115
rect 3424 27072 3476 27081
rect 3424 26936 3476 26988
rect 4160 27072 4212 27124
rect 3792 26979 3844 26988
rect 3792 26945 3801 26979
rect 3801 26945 3835 26979
rect 3835 26945 3844 26979
rect 3792 26936 3844 26945
rect 4436 27004 4488 27056
rect 4068 26936 4120 26988
rect 4804 27072 4856 27124
rect 4988 27072 5040 27124
rect 4712 27004 4764 27056
rect 6092 27072 6144 27124
rect 6276 27072 6328 27124
rect 8208 27072 8260 27124
rect 8300 27115 8352 27124
rect 8300 27081 8309 27115
rect 8309 27081 8343 27115
rect 8343 27081 8352 27115
rect 8300 27072 8352 27081
rect 8576 27115 8628 27124
rect 8576 27081 8585 27115
rect 8585 27081 8619 27115
rect 8619 27081 8628 27115
rect 8576 27072 8628 27081
rect 8944 27072 8996 27124
rect 9128 27072 9180 27124
rect 9496 27072 9548 27124
rect 10140 27072 10192 27124
rect 10692 27072 10744 27124
rect 11244 27072 11296 27124
rect 11520 27072 11572 27124
rect 1860 26911 1912 26920
rect 1860 26877 1869 26911
rect 1869 26877 1903 26911
rect 1903 26877 1912 26911
rect 1860 26868 1912 26877
rect 3516 26868 3568 26920
rect 4344 26868 4396 26920
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 7656 27004 7708 27056
rect 5172 26936 5224 26988
rect 5264 26979 5316 26988
rect 5264 26945 5273 26979
rect 5273 26945 5307 26979
rect 5307 26945 5316 26979
rect 5264 26936 5316 26945
rect 5540 26979 5592 26988
rect 5540 26945 5549 26979
rect 5549 26945 5583 26979
rect 5583 26945 5592 26979
rect 5540 26936 5592 26945
rect 5724 26979 5776 26988
rect 5724 26945 5731 26979
rect 5731 26945 5776 26979
rect 5724 26936 5776 26945
rect 5908 26979 5960 26988
rect 5908 26945 5917 26979
rect 5917 26945 5951 26979
rect 5951 26945 5960 26979
rect 5908 26936 5960 26945
rect 4988 26868 5040 26920
rect 5448 26868 5500 26920
rect 6368 26979 6420 26988
rect 6368 26945 6377 26979
rect 6377 26945 6411 26979
rect 6411 26945 6420 26979
rect 6368 26936 6420 26945
rect 6460 26979 6512 26988
rect 6460 26945 6470 26979
rect 6470 26945 6504 26979
rect 6504 26945 6512 26979
rect 6460 26936 6512 26945
rect 6736 26979 6788 26988
rect 6736 26945 6745 26979
rect 6745 26945 6779 26979
rect 6779 26945 6788 26979
rect 6736 26936 6788 26945
rect 6828 26936 6880 26988
rect 7564 26936 7616 26988
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 7288 26868 7340 26920
rect 8024 26868 8076 26920
rect 4804 26800 4856 26852
rect 5172 26800 5224 26852
rect 8392 26936 8444 26988
rect 8668 26936 8720 26988
rect 8760 26979 8812 26988
rect 8760 26945 8769 26979
rect 8769 26945 8803 26979
rect 8803 26945 8812 26979
rect 8760 26936 8812 26945
rect 8852 26936 8904 26988
rect 9220 27047 9272 27056
rect 9220 27013 9229 27047
rect 9229 27013 9263 27047
rect 9263 27013 9272 27047
rect 9220 27004 9272 27013
rect 8300 26868 8352 26920
rect 11428 27004 11480 27056
rect 5448 26732 5500 26784
rect 6184 26732 6236 26784
rect 6460 26732 6512 26784
rect 7012 26775 7064 26784
rect 7012 26741 7021 26775
rect 7021 26741 7055 26775
rect 7055 26741 7064 26775
rect 7012 26732 7064 26741
rect 7472 26775 7524 26784
rect 7472 26741 7481 26775
rect 7481 26741 7515 26775
rect 7515 26741 7524 26775
rect 7472 26732 7524 26741
rect 8760 26800 8812 26852
rect 9312 26800 9364 26852
rect 10600 26936 10652 26988
rect 11152 26936 11204 26988
rect 11336 26868 11388 26920
rect 9680 26732 9732 26784
rect 11704 26979 11756 26988
rect 11704 26945 11713 26979
rect 11713 26945 11747 26979
rect 11747 26945 11756 26979
rect 11704 26936 11756 26945
rect 12808 27072 12860 27124
rect 13176 27072 13228 27124
rect 13544 27072 13596 27124
rect 14464 27072 14516 27124
rect 15568 27072 15620 27124
rect 17132 27072 17184 27124
rect 18052 27115 18104 27124
rect 18052 27081 18061 27115
rect 18061 27081 18095 27115
rect 18095 27081 18104 27115
rect 18052 27072 18104 27081
rect 18328 27072 18380 27124
rect 18604 27072 18656 27124
rect 20628 27072 20680 27124
rect 20720 27072 20772 27124
rect 22928 27072 22980 27124
rect 26516 27072 26568 27124
rect 11980 26979 12032 26988
rect 11980 26945 11989 26979
rect 11989 26945 12023 26979
rect 12023 26945 12032 26979
rect 11980 26936 12032 26945
rect 11612 26868 11664 26920
rect 12164 26979 12216 26988
rect 12164 26945 12178 26979
rect 12178 26945 12212 26979
rect 12212 26945 12216 26979
rect 12164 26936 12216 26945
rect 12900 26979 12952 26988
rect 12900 26945 12909 26979
rect 12909 26945 12943 26979
rect 12943 26945 12952 26979
rect 12900 26936 12952 26945
rect 12992 26936 13044 26988
rect 12624 26868 12676 26920
rect 15384 27004 15436 27056
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 13636 26868 13688 26920
rect 14556 26979 14608 26988
rect 14556 26945 14565 26979
rect 14565 26945 14599 26979
rect 14599 26945 14608 26979
rect 14556 26936 14608 26945
rect 14280 26868 14332 26920
rect 15200 26936 15252 26988
rect 14740 26868 14792 26920
rect 15016 26868 15068 26920
rect 17224 27004 17276 27056
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 18420 26979 18472 26988
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18420 26936 18472 26945
rect 16764 26868 16816 26920
rect 17224 26868 17276 26920
rect 18604 26911 18656 26920
rect 18604 26877 18613 26911
rect 18613 26877 18647 26911
rect 18647 26877 18656 26911
rect 18604 26868 18656 26877
rect 20352 26936 20404 26988
rect 20904 26936 20956 26988
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 22284 26979 22336 26988
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 22652 26936 22704 26988
rect 17684 26800 17736 26852
rect 20536 26868 20588 26920
rect 20812 26868 20864 26920
rect 21180 26868 21232 26920
rect 23296 26868 23348 26920
rect 13820 26732 13872 26784
rect 15108 26732 15160 26784
rect 17316 26732 17368 26784
rect 17868 26732 17920 26784
rect 17960 26775 18012 26784
rect 17960 26741 17969 26775
rect 17969 26741 18003 26775
rect 18003 26741 18012 26775
rect 17960 26732 18012 26741
rect 18788 26732 18840 26784
rect 19432 26732 19484 26784
rect 19892 26732 19944 26784
rect 23480 26979 23532 26988
rect 23480 26945 23489 26979
rect 23489 26945 23523 26979
rect 23523 26945 23532 26979
rect 23480 26936 23532 26945
rect 25228 27004 25280 27056
rect 26332 27004 26384 27056
rect 27160 27072 27212 27124
rect 27620 27072 27672 27124
rect 27988 27072 28040 27124
rect 28080 27072 28132 27124
rect 29460 27072 29512 27124
rect 30012 27072 30064 27124
rect 30932 27072 30984 27124
rect 31116 27072 31168 27124
rect 24952 26936 25004 26988
rect 25044 26979 25096 26988
rect 25044 26945 25053 26979
rect 25053 26945 25087 26979
rect 25087 26945 25096 26979
rect 25044 26936 25096 26945
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 26148 26936 26200 26988
rect 24400 26911 24452 26920
rect 24400 26877 24409 26911
rect 24409 26877 24443 26911
rect 24443 26877 24452 26911
rect 24400 26868 24452 26877
rect 24492 26868 24544 26920
rect 25320 26868 25372 26920
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 27620 26936 27672 26988
rect 27344 26868 27396 26920
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 27896 26936 27948 26945
rect 27988 26936 28040 26988
rect 28356 26936 28408 26988
rect 28816 26979 28868 26988
rect 28816 26945 28819 26979
rect 28819 26945 28853 26979
rect 28853 26945 28868 26979
rect 28816 26936 28868 26945
rect 31852 27004 31904 27056
rect 33784 27072 33836 27124
rect 34060 27072 34112 27124
rect 20536 26775 20588 26784
rect 20536 26741 20545 26775
rect 20545 26741 20579 26775
rect 20579 26741 20588 26775
rect 20536 26732 20588 26741
rect 20720 26732 20772 26784
rect 22192 26732 22244 26784
rect 26516 26800 26568 26852
rect 25688 26775 25740 26784
rect 25688 26741 25697 26775
rect 25697 26741 25731 26775
rect 25731 26741 25740 26775
rect 25688 26732 25740 26741
rect 26792 26775 26844 26784
rect 26792 26741 26801 26775
rect 26801 26741 26835 26775
rect 26835 26741 26844 26775
rect 26792 26732 26844 26741
rect 27436 26732 27488 26784
rect 28356 26800 28408 26852
rect 29736 26843 29788 26852
rect 29736 26809 29745 26843
rect 29745 26809 29779 26843
rect 29779 26809 29788 26843
rect 30196 26868 30248 26920
rect 30748 26936 30800 26988
rect 30840 26979 30892 26988
rect 30840 26945 30849 26979
rect 30849 26945 30883 26979
rect 30883 26945 30892 26979
rect 30840 26936 30892 26945
rect 30932 26979 30984 26988
rect 30932 26945 30941 26979
rect 30941 26945 30975 26979
rect 30975 26945 30984 26979
rect 30932 26936 30984 26945
rect 31024 26979 31076 26988
rect 31024 26945 31033 26979
rect 31033 26945 31067 26979
rect 31067 26945 31076 26979
rect 31024 26936 31076 26945
rect 31208 26979 31260 26988
rect 31208 26945 31217 26979
rect 31217 26945 31251 26979
rect 31251 26945 31260 26979
rect 31208 26936 31260 26945
rect 31300 26979 31352 26988
rect 31300 26945 31309 26979
rect 31309 26945 31343 26979
rect 31343 26945 31352 26979
rect 31300 26936 31352 26945
rect 31944 26936 31996 26988
rect 32128 26979 32180 26988
rect 32128 26945 32137 26979
rect 32137 26945 32171 26979
rect 32171 26945 32180 26979
rect 32128 26936 32180 26945
rect 32220 26936 32272 26988
rect 33876 26868 33928 26920
rect 29736 26800 29788 26809
rect 31852 26800 31904 26852
rect 27712 26775 27764 26784
rect 27712 26741 27721 26775
rect 27721 26741 27755 26775
rect 27755 26741 27764 26775
rect 27712 26732 27764 26741
rect 28080 26775 28132 26784
rect 28080 26741 28089 26775
rect 28089 26741 28123 26775
rect 28123 26741 28132 26775
rect 28080 26732 28132 26741
rect 28632 26775 28684 26784
rect 28632 26741 28641 26775
rect 28641 26741 28675 26775
rect 28675 26741 28684 26775
rect 28632 26732 28684 26741
rect 28908 26732 28960 26784
rect 29460 26732 29512 26784
rect 29828 26732 29880 26784
rect 30380 26732 30432 26784
rect 30564 26775 30616 26784
rect 30564 26741 30573 26775
rect 30573 26741 30607 26775
rect 30607 26741 30616 26775
rect 30564 26732 30616 26741
rect 30656 26732 30708 26784
rect 31484 26732 31536 26784
rect 32036 26732 32088 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4804 26528 4856 26580
rect 5632 26528 5684 26580
rect 7748 26528 7800 26580
rect 8208 26528 8260 26580
rect 1584 26460 1636 26512
rect 4436 26460 4488 26512
rect 4988 26460 5040 26512
rect 5172 26460 5224 26512
rect 4344 26392 4396 26444
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 3884 26324 3936 26376
rect 5080 26324 5132 26376
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 5908 26460 5960 26512
rect 6460 26460 6512 26512
rect 7564 26460 7616 26512
rect 11244 26528 11296 26580
rect 12992 26528 13044 26580
rect 16120 26528 16172 26580
rect 17684 26528 17736 26580
rect 17776 26528 17828 26580
rect 17960 26528 18012 26580
rect 2780 26256 2832 26308
rect 3792 26256 3844 26308
rect 3976 26256 4028 26308
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 6828 26324 6880 26376
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 7380 26367 7432 26376
rect 7380 26333 7390 26367
rect 7390 26333 7424 26367
rect 7424 26333 7432 26367
rect 8300 26435 8352 26444
rect 8300 26401 8309 26435
rect 8309 26401 8343 26435
rect 8343 26401 8352 26435
rect 8300 26392 8352 26401
rect 8392 26392 8444 26444
rect 7380 26324 7432 26333
rect 8208 26324 8260 26376
rect 5632 26256 5684 26308
rect 3700 26188 3752 26240
rect 5172 26188 5224 26240
rect 5540 26188 5592 26240
rect 5816 26188 5868 26240
rect 6000 26188 6052 26240
rect 7564 26299 7616 26308
rect 7564 26265 7573 26299
rect 7573 26265 7607 26299
rect 7607 26265 7616 26299
rect 7564 26256 7616 26265
rect 8116 26256 8168 26308
rect 9220 26367 9272 26376
rect 9220 26333 9229 26367
rect 9229 26333 9263 26367
rect 9263 26333 9272 26367
rect 9220 26324 9272 26333
rect 9404 26324 9456 26376
rect 8852 26256 8904 26308
rect 9036 26256 9088 26308
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 10876 26392 10928 26444
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 11244 26392 11296 26444
rect 11520 26392 11572 26444
rect 10968 26324 11020 26376
rect 11796 26324 11848 26376
rect 12532 26324 12584 26376
rect 14004 26392 14056 26444
rect 14372 26392 14424 26444
rect 15752 26460 15804 26512
rect 13728 26324 13780 26376
rect 13820 26367 13872 26376
rect 13820 26333 13829 26367
rect 13829 26333 13863 26367
rect 13863 26333 13872 26367
rect 13820 26324 13872 26333
rect 12348 26256 12400 26308
rect 12440 26256 12492 26308
rect 14556 26299 14608 26308
rect 14556 26265 14565 26299
rect 14565 26265 14599 26299
rect 14599 26265 14608 26299
rect 14556 26256 14608 26265
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 15384 26324 15436 26376
rect 15660 26392 15712 26444
rect 16948 26460 17000 26512
rect 15936 26324 15988 26376
rect 16396 26324 16448 26376
rect 16488 26324 16540 26376
rect 16672 26324 16724 26376
rect 16764 26324 16816 26376
rect 7104 26188 7156 26240
rect 7748 26188 7800 26240
rect 10324 26188 10376 26240
rect 10508 26188 10560 26240
rect 11060 26188 11112 26240
rect 14464 26188 14516 26240
rect 15108 26231 15160 26240
rect 15108 26197 15117 26231
rect 15117 26197 15151 26231
rect 15151 26197 15160 26231
rect 15108 26188 15160 26197
rect 15844 26188 15896 26240
rect 16948 26299 17000 26308
rect 16948 26265 16957 26299
rect 16957 26265 16991 26299
rect 16991 26265 17000 26299
rect 16948 26256 17000 26265
rect 17316 26256 17368 26308
rect 18788 26460 18840 26512
rect 20076 26528 20128 26580
rect 20628 26528 20680 26580
rect 22284 26528 22336 26580
rect 23480 26571 23532 26580
rect 23480 26537 23489 26571
rect 23489 26537 23523 26571
rect 23523 26537 23532 26571
rect 23480 26528 23532 26537
rect 23756 26528 23808 26580
rect 24584 26528 24636 26580
rect 25044 26528 25096 26580
rect 25872 26528 25924 26580
rect 26056 26528 26108 26580
rect 26240 26571 26292 26580
rect 26240 26537 26249 26571
rect 26249 26537 26283 26571
rect 26283 26537 26292 26571
rect 26240 26528 26292 26537
rect 26884 26528 26936 26580
rect 27620 26528 27672 26580
rect 28448 26528 28500 26580
rect 20812 26460 20864 26512
rect 17776 26367 17828 26376
rect 17776 26333 17785 26367
rect 17785 26333 17819 26367
rect 17819 26333 17828 26367
rect 17776 26324 17828 26333
rect 18236 26324 18288 26376
rect 18420 26392 18472 26444
rect 18880 26435 18932 26444
rect 18880 26401 18889 26435
rect 18889 26401 18923 26435
rect 18923 26401 18932 26435
rect 18880 26392 18932 26401
rect 19156 26392 19208 26444
rect 16396 26231 16448 26240
rect 16396 26197 16405 26231
rect 16405 26197 16439 26231
rect 16439 26197 16448 26231
rect 16396 26188 16448 26197
rect 16672 26231 16724 26240
rect 16672 26197 16681 26231
rect 16681 26197 16715 26231
rect 16715 26197 16724 26231
rect 16672 26188 16724 26197
rect 17224 26188 17276 26240
rect 21180 26435 21232 26444
rect 21180 26401 21189 26435
rect 21189 26401 21223 26435
rect 21223 26401 21232 26435
rect 21180 26392 21232 26401
rect 21364 26392 21416 26444
rect 21732 26435 21784 26444
rect 21732 26401 21741 26435
rect 21741 26401 21775 26435
rect 21775 26401 21784 26435
rect 21732 26392 21784 26401
rect 19965 26367 20017 26376
rect 19965 26333 19974 26367
rect 19974 26333 20008 26367
rect 20008 26333 20017 26367
rect 19965 26324 20017 26333
rect 20076 26367 20128 26376
rect 20076 26333 20085 26367
rect 20085 26333 20119 26367
rect 20119 26333 20128 26367
rect 20076 26324 20128 26333
rect 20352 26324 20404 26376
rect 20628 26324 20680 26376
rect 21548 26367 21600 26376
rect 21548 26333 21557 26367
rect 21557 26333 21591 26367
rect 21591 26333 21600 26367
rect 21548 26324 21600 26333
rect 20720 26256 20772 26308
rect 20996 26256 21048 26308
rect 22008 26367 22060 26376
rect 22008 26333 22017 26367
rect 22017 26333 22051 26367
rect 22051 26333 22060 26367
rect 22008 26324 22060 26333
rect 22652 26324 22704 26376
rect 23296 26324 23348 26376
rect 23756 26367 23808 26376
rect 23756 26333 23763 26367
rect 23763 26333 23808 26367
rect 23756 26324 23808 26333
rect 25412 26392 25464 26444
rect 25504 26392 25556 26444
rect 20444 26188 20496 26240
rect 20536 26231 20588 26240
rect 20536 26197 20545 26231
rect 20545 26197 20579 26231
rect 20579 26197 20588 26231
rect 20536 26188 20588 26197
rect 21088 26188 21140 26240
rect 23480 26256 23532 26308
rect 23940 26299 23992 26308
rect 23940 26265 23949 26299
rect 23949 26265 23983 26299
rect 23983 26265 23992 26299
rect 23940 26256 23992 26265
rect 25320 26324 25372 26376
rect 25780 26367 25832 26376
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 25780 26324 25832 26333
rect 24308 26256 24360 26308
rect 25964 26392 26016 26444
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 26424 26324 26476 26376
rect 27252 26324 27304 26376
rect 27620 26435 27672 26444
rect 27620 26401 27629 26435
rect 27629 26401 27663 26435
rect 27663 26401 27672 26435
rect 27620 26392 27672 26401
rect 27804 26367 27856 26370
rect 27804 26333 27813 26367
rect 27813 26333 27847 26367
rect 27847 26333 27856 26367
rect 27804 26318 27856 26333
rect 28908 26528 28960 26580
rect 28724 26460 28776 26512
rect 30748 26571 30800 26580
rect 30748 26537 30757 26571
rect 30757 26537 30791 26571
rect 30791 26537 30800 26571
rect 30748 26528 30800 26537
rect 31116 26528 31168 26580
rect 31300 26528 31352 26580
rect 33876 26571 33928 26580
rect 33876 26537 33885 26571
rect 33885 26537 33919 26571
rect 33919 26537 33928 26571
rect 33876 26528 33928 26537
rect 32772 26460 32824 26512
rect 28908 26392 28960 26444
rect 29552 26392 29604 26444
rect 30380 26392 30432 26444
rect 28448 26256 28500 26308
rect 26424 26188 26476 26240
rect 26792 26188 26844 26240
rect 27252 26231 27304 26240
rect 27252 26197 27261 26231
rect 27261 26197 27295 26231
rect 27295 26197 27304 26231
rect 27252 26188 27304 26197
rect 27988 26188 28040 26240
rect 28540 26231 28592 26240
rect 28540 26197 28549 26231
rect 28549 26197 28583 26231
rect 28583 26197 28592 26231
rect 28540 26188 28592 26197
rect 28724 26188 28776 26240
rect 29000 26231 29052 26240
rect 29000 26197 29009 26231
rect 29009 26197 29043 26231
rect 29043 26197 29052 26231
rect 29000 26188 29052 26197
rect 29092 26188 29144 26240
rect 29552 26231 29604 26240
rect 29552 26197 29561 26231
rect 29561 26197 29595 26231
rect 29595 26197 29604 26231
rect 29552 26188 29604 26197
rect 29828 26367 29880 26376
rect 29828 26333 29837 26367
rect 29837 26333 29871 26367
rect 29871 26333 29880 26367
rect 29828 26324 29880 26333
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 30196 26367 30248 26376
rect 30196 26333 30205 26367
rect 30205 26333 30239 26367
rect 30239 26333 30248 26367
rect 30196 26324 30248 26333
rect 30288 26299 30340 26308
rect 30288 26265 30297 26299
rect 30297 26265 30331 26299
rect 30331 26265 30340 26299
rect 30288 26256 30340 26265
rect 30656 26367 30708 26376
rect 30656 26333 30665 26367
rect 30665 26333 30699 26367
rect 30699 26333 30708 26367
rect 30656 26324 30708 26333
rect 30932 26324 30984 26376
rect 31208 26324 31260 26376
rect 32036 26299 32088 26308
rect 32036 26265 32070 26299
rect 32070 26265 32088 26299
rect 32036 26256 32088 26265
rect 32128 26256 32180 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3240 25848 3292 25900
rect 3884 25984 3936 26036
rect 4896 25984 4948 26036
rect 5080 25984 5132 26036
rect 3700 25959 3752 25968
rect 3700 25925 3709 25959
rect 3709 25925 3743 25959
rect 3743 25925 3752 25959
rect 3700 25916 3752 25925
rect 3884 25848 3936 25900
rect 1400 25823 1452 25832
rect 1400 25789 1409 25823
rect 1409 25789 1443 25823
rect 1443 25789 1452 25823
rect 1400 25780 1452 25789
rect 4344 25848 4396 25900
rect 5172 25916 5224 25968
rect 5816 25984 5868 26036
rect 6736 25984 6788 26036
rect 4712 25891 4764 25900
rect 4712 25857 4721 25891
rect 4721 25857 4755 25891
rect 4755 25857 4764 25891
rect 4712 25848 4764 25857
rect 4988 25848 5040 25900
rect 5080 25891 5132 25900
rect 5080 25857 5089 25891
rect 5089 25857 5123 25891
rect 5123 25857 5132 25891
rect 5080 25848 5132 25857
rect 5264 25891 5316 25900
rect 5264 25857 5273 25891
rect 5273 25857 5307 25891
rect 5307 25857 5316 25891
rect 5264 25848 5316 25857
rect 3976 25644 4028 25696
rect 4620 25780 4672 25832
rect 5632 25848 5684 25900
rect 5724 25848 5776 25900
rect 6552 25848 6604 25900
rect 7932 25916 7984 25968
rect 6368 25780 6420 25832
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 7012 25848 7064 25857
rect 7104 25891 7156 25900
rect 7104 25857 7113 25891
rect 7113 25857 7147 25891
rect 7147 25857 7156 25891
rect 7104 25848 7156 25857
rect 8484 25916 8536 25968
rect 9036 26027 9088 26036
rect 9036 25993 9045 26027
rect 9045 25993 9079 26027
rect 9079 25993 9088 26027
rect 9036 25984 9088 25993
rect 9496 26027 9548 26036
rect 9496 25993 9505 26027
rect 9505 25993 9539 26027
rect 9539 25993 9548 26027
rect 9496 25984 9548 25993
rect 10048 25984 10100 26036
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 10692 25916 10744 25968
rect 10968 25959 11020 25968
rect 10968 25925 10977 25959
rect 10977 25925 11011 25959
rect 11011 25925 11020 25959
rect 10968 25916 11020 25925
rect 11060 25959 11112 25968
rect 11060 25925 11069 25959
rect 11069 25925 11103 25959
rect 11103 25925 11112 25959
rect 11060 25916 11112 25925
rect 8300 25848 8352 25900
rect 9036 25848 9088 25900
rect 8024 25780 8076 25832
rect 8208 25780 8260 25832
rect 10508 25848 10560 25900
rect 10876 25848 10928 25900
rect 11612 25984 11664 26036
rect 12440 25984 12492 26036
rect 13452 26027 13504 26036
rect 13452 25993 13461 26027
rect 13461 25993 13495 26027
rect 13495 25993 13504 26027
rect 13452 25984 13504 25993
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 14372 25984 14424 26036
rect 15292 25984 15344 26036
rect 15660 25984 15712 26036
rect 16488 25984 16540 26036
rect 16672 25984 16724 26036
rect 19984 25984 20036 26036
rect 20076 25984 20128 26036
rect 11520 25959 11572 25968
rect 11520 25925 11529 25959
rect 11529 25925 11563 25959
rect 11563 25925 11572 25959
rect 11520 25916 11572 25925
rect 12164 25780 12216 25832
rect 16396 25916 16448 25968
rect 13636 25891 13688 25900
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 5080 25644 5132 25696
rect 5632 25644 5684 25696
rect 6644 25687 6696 25696
rect 6644 25653 6653 25687
rect 6653 25653 6687 25687
rect 6687 25653 6696 25687
rect 6644 25644 6696 25653
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 7288 25644 7340 25653
rect 7748 25644 7800 25696
rect 8484 25712 8536 25764
rect 8760 25712 8812 25764
rect 11336 25712 11388 25764
rect 8576 25644 8628 25696
rect 9312 25644 9364 25696
rect 11060 25644 11112 25696
rect 11980 25644 12032 25696
rect 12808 25780 12860 25832
rect 14188 25848 14240 25900
rect 15476 25848 15528 25900
rect 15660 25848 15712 25900
rect 15844 25891 15896 25900
rect 15844 25857 15853 25891
rect 15853 25857 15887 25891
rect 15887 25857 15896 25891
rect 15844 25848 15896 25857
rect 17960 25916 18012 25968
rect 20536 25984 20588 26036
rect 21640 26027 21692 26036
rect 21640 25993 21649 26027
rect 21649 25993 21683 26027
rect 21683 25993 21692 26027
rect 21640 25984 21692 25993
rect 23388 25984 23440 26036
rect 16580 25848 16632 25900
rect 18604 25848 18656 25900
rect 19064 25848 19116 25900
rect 12532 25712 12584 25764
rect 13268 25755 13320 25764
rect 13268 25721 13277 25755
rect 13277 25721 13311 25755
rect 13311 25721 13320 25755
rect 13268 25712 13320 25721
rect 16396 25780 16448 25832
rect 16488 25780 16540 25832
rect 20720 25891 20772 25900
rect 20720 25857 20729 25891
rect 20729 25857 20763 25891
rect 20763 25857 20772 25891
rect 20720 25848 20772 25857
rect 20812 25823 20864 25832
rect 20812 25789 20821 25823
rect 20821 25789 20855 25823
rect 20855 25789 20864 25823
rect 20812 25780 20864 25789
rect 20996 25848 21048 25900
rect 24400 25959 24452 25968
rect 24400 25925 24409 25959
rect 24409 25925 24443 25959
rect 24443 25925 24452 25959
rect 24400 25916 24452 25925
rect 21640 25780 21692 25832
rect 22468 25891 22520 25900
rect 22468 25857 22477 25891
rect 22477 25857 22511 25891
rect 22511 25857 22520 25891
rect 22468 25848 22520 25857
rect 22928 25891 22980 25900
rect 22928 25857 22937 25891
rect 22937 25857 22971 25891
rect 22971 25857 22980 25891
rect 22928 25848 22980 25857
rect 23204 25848 23256 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 23664 25891 23716 25900
rect 23664 25857 23673 25891
rect 23673 25857 23707 25891
rect 23707 25857 23716 25891
rect 23664 25848 23716 25857
rect 24216 25891 24268 25900
rect 24216 25857 24225 25891
rect 24225 25857 24259 25891
rect 24259 25857 24268 25891
rect 24216 25848 24268 25857
rect 25780 25916 25832 25968
rect 25964 25916 26016 25968
rect 27896 25984 27948 26036
rect 27988 25984 28040 26036
rect 28816 25984 28868 26036
rect 29552 25984 29604 26036
rect 27344 25916 27396 25968
rect 27712 25959 27764 25968
rect 27712 25925 27721 25959
rect 27721 25925 27755 25959
rect 27755 25925 27764 25959
rect 27712 25916 27764 25925
rect 29460 25916 29512 25968
rect 32588 25984 32640 26036
rect 23480 25780 23532 25832
rect 24124 25780 24176 25832
rect 24308 25780 24360 25832
rect 25596 25848 25648 25900
rect 24860 25780 24912 25832
rect 25228 25823 25280 25832
rect 25228 25789 25237 25823
rect 25237 25789 25271 25823
rect 25271 25789 25280 25823
rect 25228 25780 25280 25789
rect 26056 25780 26108 25832
rect 14464 25644 14516 25696
rect 15292 25687 15344 25696
rect 15292 25653 15301 25687
rect 15301 25653 15335 25687
rect 15335 25653 15344 25687
rect 15292 25644 15344 25653
rect 15660 25712 15712 25764
rect 15752 25755 15804 25764
rect 15752 25721 15761 25755
rect 15761 25721 15795 25755
rect 15795 25721 15804 25755
rect 15752 25712 15804 25721
rect 15936 25755 15988 25764
rect 15936 25721 15945 25755
rect 15945 25721 15979 25755
rect 15979 25721 15988 25755
rect 15936 25712 15988 25721
rect 16672 25712 16724 25764
rect 18236 25712 18288 25764
rect 19248 25712 19300 25764
rect 22376 25712 22428 25764
rect 26240 25891 26292 25900
rect 26240 25857 26249 25891
rect 26249 25857 26283 25891
rect 26283 25857 26292 25891
rect 26240 25848 26292 25857
rect 28172 25848 28224 25900
rect 31852 25916 31904 25968
rect 28448 25780 28500 25832
rect 28908 25823 28960 25832
rect 28908 25789 28917 25823
rect 28917 25789 28951 25823
rect 28951 25789 28960 25823
rect 28908 25780 28960 25789
rect 30104 25848 30156 25900
rect 32128 25891 32180 25900
rect 32128 25857 32137 25891
rect 32137 25857 32171 25891
rect 32171 25857 32180 25891
rect 32128 25848 32180 25857
rect 31116 25823 31168 25832
rect 31116 25789 31125 25823
rect 31125 25789 31159 25823
rect 31159 25789 31168 25823
rect 31116 25780 31168 25789
rect 16212 25644 16264 25696
rect 17500 25644 17552 25696
rect 18512 25644 18564 25696
rect 19156 25687 19208 25696
rect 19156 25653 19165 25687
rect 19165 25653 19199 25687
rect 19199 25653 19208 25687
rect 19156 25644 19208 25653
rect 19892 25644 19944 25696
rect 20628 25644 20680 25696
rect 21088 25644 21140 25696
rect 21456 25644 21508 25696
rect 23388 25644 23440 25696
rect 27712 25712 27764 25764
rect 28264 25712 28316 25764
rect 26792 25644 26844 25696
rect 27620 25644 27672 25696
rect 28724 25712 28776 25764
rect 29092 25712 29144 25764
rect 29184 25712 29236 25764
rect 29552 25712 29604 25764
rect 30932 25755 30984 25764
rect 30932 25721 30941 25755
rect 30941 25721 30975 25755
rect 30975 25721 30984 25755
rect 30932 25712 30984 25721
rect 30840 25644 30892 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3240 25483 3292 25492
rect 3240 25449 3249 25483
rect 3249 25449 3283 25483
rect 3283 25449 3292 25483
rect 3240 25440 3292 25449
rect 3700 25440 3752 25492
rect 5264 25440 5316 25492
rect 5448 25440 5500 25492
rect 6184 25440 6236 25492
rect 3332 25372 3384 25424
rect 3884 25372 3936 25424
rect 2688 25304 2740 25356
rect 4712 25304 4764 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 2044 25236 2096 25288
rect 1768 25168 1820 25220
rect 1492 25100 1544 25152
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 3976 25236 4028 25288
rect 5172 25236 5224 25288
rect 4988 25211 5040 25220
rect 4988 25177 4997 25211
rect 4997 25177 5031 25211
rect 5031 25177 5040 25211
rect 5632 25236 5684 25288
rect 5724 25279 5776 25288
rect 5724 25245 5733 25279
rect 5733 25245 5767 25279
rect 5767 25245 5776 25279
rect 5724 25236 5776 25245
rect 5816 25279 5868 25288
rect 5816 25245 5826 25279
rect 5826 25245 5860 25279
rect 5860 25245 5868 25279
rect 5816 25236 5868 25245
rect 6000 25279 6052 25288
rect 6000 25245 6009 25279
rect 6009 25245 6043 25279
rect 6043 25245 6052 25279
rect 6000 25236 6052 25245
rect 6828 25304 6880 25356
rect 7196 25415 7248 25424
rect 7196 25381 7205 25415
rect 7205 25381 7239 25415
rect 7239 25381 7248 25415
rect 7196 25372 7248 25381
rect 7380 25372 7432 25424
rect 6460 25279 6512 25288
rect 6460 25245 6469 25279
rect 6469 25245 6503 25279
rect 6503 25245 6512 25279
rect 6460 25236 6512 25245
rect 6552 25279 6604 25288
rect 6552 25245 6562 25279
rect 6562 25245 6596 25279
rect 6596 25245 6604 25279
rect 6552 25236 6604 25245
rect 6736 25279 6788 25288
rect 6736 25245 6745 25279
rect 6745 25245 6779 25279
rect 6779 25245 6788 25279
rect 6736 25236 6788 25245
rect 7104 25236 7156 25288
rect 8484 25440 8536 25492
rect 8760 25440 8812 25492
rect 11520 25440 11572 25492
rect 11980 25483 12032 25492
rect 11980 25449 11989 25483
rect 11989 25449 12023 25483
rect 12023 25449 12032 25483
rect 11980 25440 12032 25449
rect 14280 25440 14332 25492
rect 14740 25440 14792 25492
rect 8300 25372 8352 25424
rect 10232 25372 10284 25424
rect 4988 25168 5040 25177
rect 3424 25100 3476 25152
rect 4068 25100 4120 25152
rect 4896 25100 4948 25152
rect 5264 25100 5316 25152
rect 5540 25100 5592 25152
rect 6460 25100 6512 25152
rect 6736 25100 6788 25152
rect 8208 25236 8260 25288
rect 8576 25236 8628 25288
rect 7932 25168 7984 25220
rect 8392 25211 8444 25220
rect 8392 25177 8401 25211
rect 8401 25177 8435 25211
rect 8435 25177 8444 25211
rect 8392 25168 8444 25177
rect 8668 25168 8720 25220
rect 9220 25279 9272 25288
rect 9220 25245 9229 25279
rect 9229 25245 9263 25279
rect 9263 25245 9272 25279
rect 9220 25236 9272 25245
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9496 25236 9548 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 10324 25236 10376 25288
rect 7472 25100 7524 25152
rect 7656 25100 7708 25152
rect 8208 25100 8260 25152
rect 10140 25211 10192 25220
rect 10140 25177 10149 25211
rect 10149 25177 10183 25211
rect 10183 25177 10192 25211
rect 10140 25168 10192 25177
rect 10416 25100 10468 25152
rect 10600 25236 10652 25288
rect 11060 25236 11112 25288
rect 11152 25279 11204 25288
rect 11152 25245 11161 25279
rect 11161 25245 11195 25279
rect 11195 25245 11204 25279
rect 11152 25236 11204 25245
rect 11520 25236 11572 25288
rect 11612 25279 11664 25288
rect 11612 25245 11621 25279
rect 11621 25245 11655 25279
rect 11655 25245 11664 25279
rect 11612 25236 11664 25245
rect 10600 25100 10652 25152
rect 10968 25168 11020 25220
rect 11980 25236 12032 25288
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 14372 25372 14424 25424
rect 13728 25236 13780 25288
rect 11152 25100 11204 25152
rect 13544 25168 13596 25220
rect 14188 25236 14240 25288
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 14648 25236 14700 25288
rect 14004 25168 14056 25220
rect 14740 25168 14792 25220
rect 15384 25372 15436 25424
rect 16212 25440 16264 25492
rect 16304 25483 16356 25492
rect 16304 25449 16313 25483
rect 16313 25449 16347 25483
rect 16347 25449 16356 25483
rect 16304 25440 16356 25449
rect 16580 25483 16632 25492
rect 16580 25449 16589 25483
rect 16589 25449 16623 25483
rect 16623 25449 16632 25483
rect 16580 25440 16632 25449
rect 17132 25440 17184 25492
rect 17500 25483 17552 25492
rect 17500 25449 17509 25483
rect 17509 25449 17543 25483
rect 17543 25449 17552 25483
rect 17500 25440 17552 25449
rect 17776 25440 17828 25492
rect 18420 25440 18472 25492
rect 19524 25440 19576 25492
rect 16028 25347 16080 25356
rect 16028 25313 16037 25347
rect 16037 25313 16071 25347
rect 16071 25313 16080 25347
rect 16028 25304 16080 25313
rect 16856 25372 16908 25424
rect 15292 25236 15344 25288
rect 15936 25236 15988 25288
rect 16304 25236 16356 25288
rect 16672 25347 16724 25356
rect 16672 25313 16681 25347
rect 16681 25313 16715 25347
rect 16715 25313 16724 25347
rect 16672 25304 16724 25313
rect 17500 25304 17552 25356
rect 18236 25372 18288 25424
rect 18972 25372 19024 25424
rect 17408 25236 17460 25288
rect 18512 25236 18564 25288
rect 19340 25236 19392 25288
rect 20168 25483 20220 25492
rect 20168 25449 20177 25483
rect 20177 25449 20211 25483
rect 20211 25449 20220 25483
rect 20168 25440 20220 25449
rect 20352 25440 20404 25492
rect 20536 25440 20588 25492
rect 19892 25372 19944 25424
rect 21272 25483 21324 25492
rect 21272 25449 21281 25483
rect 21281 25449 21315 25483
rect 21315 25449 21324 25483
rect 21272 25440 21324 25449
rect 22008 25440 22060 25492
rect 22928 25483 22980 25492
rect 22928 25449 22937 25483
rect 22937 25449 22971 25483
rect 22971 25449 22980 25483
rect 22928 25440 22980 25449
rect 19984 25236 20036 25288
rect 20168 25236 20220 25288
rect 17040 25168 17092 25220
rect 17592 25168 17644 25220
rect 20444 25236 20496 25288
rect 23020 25372 23072 25424
rect 24676 25440 24728 25492
rect 25136 25440 25188 25492
rect 22836 25304 22888 25356
rect 20812 25236 20864 25288
rect 20996 25236 21048 25288
rect 21640 25236 21692 25288
rect 12900 25100 12952 25152
rect 15384 25100 15436 25152
rect 15844 25100 15896 25152
rect 16764 25100 16816 25152
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 17316 25100 17368 25152
rect 17500 25143 17552 25152
rect 17500 25109 17518 25143
rect 17518 25109 17552 25143
rect 20720 25168 20772 25220
rect 21456 25168 21508 25220
rect 17500 25100 17552 25109
rect 19800 25100 19852 25152
rect 20076 25100 20128 25152
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 22192 25279 22244 25288
rect 22192 25245 22201 25279
rect 22201 25245 22235 25279
rect 22235 25245 22244 25279
rect 22192 25236 22244 25245
rect 22376 25279 22428 25288
rect 22376 25245 22385 25279
rect 22385 25245 22419 25279
rect 22419 25245 22428 25279
rect 22376 25236 22428 25245
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 23204 25279 23256 25288
rect 23204 25245 23213 25279
rect 23213 25245 23247 25279
rect 23247 25245 23256 25279
rect 23204 25236 23256 25245
rect 24492 25372 24544 25424
rect 25412 25372 25464 25424
rect 29644 25483 29696 25492
rect 29644 25449 29653 25483
rect 29653 25449 29687 25483
rect 29687 25449 29696 25483
rect 29644 25440 29696 25449
rect 31116 25440 31168 25492
rect 32496 25483 32548 25492
rect 32496 25449 32505 25483
rect 32505 25449 32539 25483
rect 32539 25449 32548 25483
rect 32496 25440 32548 25449
rect 32956 25440 33008 25492
rect 43260 25440 43312 25492
rect 29460 25372 29512 25424
rect 29552 25372 29604 25424
rect 23940 25236 23992 25288
rect 24032 25279 24084 25288
rect 24032 25245 24041 25279
rect 24041 25245 24075 25279
rect 24075 25245 24084 25279
rect 24032 25236 24084 25245
rect 22100 25100 22152 25152
rect 22836 25143 22888 25152
rect 22836 25109 22845 25143
rect 22845 25109 22879 25143
rect 22879 25109 22888 25143
rect 22836 25100 22888 25109
rect 23296 25100 23348 25152
rect 23572 25143 23624 25152
rect 23572 25109 23581 25143
rect 23581 25109 23615 25143
rect 23615 25109 23624 25143
rect 23572 25100 23624 25109
rect 24400 25211 24452 25220
rect 24400 25177 24409 25211
rect 24409 25177 24443 25211
rect 24443 25177 24452 25211
rect 24400 25168 24452 25177
rect 24584 25236 24636 25288
rect 24860 25304 24912 25356
rect 26516 25304 26568 25356
rect 27988 25347 28040 25356
rect 27988 25313 27997 25347
rect 27997 25313 28031 25347
rect 28031 25313 28040 25347
rect 27988 25304 28040 25313
rect 28908 25304 28960 25356
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 27344 25236 27396 25288
rect 32680 25347 32732 25356
rect 32680 25313 32689 25347
rect 32689 25313 32723 25347
rect 32723 25313 32732 25347
rect 32680 25304 32732 25313
rect 25320 25168 25372 25220
rect 29092 25242 29101 25266
rect 29101 25242 29135 25266
rect 29135 25242 29144 25266
rect 29092 25214 29144 25242
rect 29276 25236 29328 25288
rect 29736 25236 29788 25288
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 31576 25236 31628 25288
rect 27252 25100 27304 25152
rect 30196 25168 30248 25220
rect 30564 25168 30616 25220
rect 29092 25100 29144 25152
rect 31760 25100 31812 25152
rect 32220 25100 32272 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1768 24939 1820 24948
rect 1768 24905 1777 24939
rect 1777 24905 1811 24939
rect 1811 24905 1820 24939
rect 1768 24896 1820 24905
rect 5172 24896 5224 24948
rect 5356 24939 5408 24948
rect 5356 24905 5365 24939
rect 5365 24905 5399 24939
rect 5399 24905 5408 24939
rect 5356 24896 5408 24905
rect 5448 24896 5500 24948
rect 6736 24896 6788 24948
rect 8668 24896 8720 24948
rect 9036 24939 9088 24948
rect 9036 24905 9045 24939
rect 9045 24905 9079 24939
rect 9079 24905 9088 24939
rect 9036 24896 9088 24905
rect 9864 24896 9916 24948
rect 2044 24828 2096 24880
rect 5080 24871 5132 24880
rect 1492 24692 1544 24744
rect 5080 24837 5089 24871
rect 5089 24837 5123 24871
rect 5123 24837 5132 24871
rect 5080 24828 5132 24837
rect 3608 24760 3660 24812
rect 3700 24760 3752 24812
rect 4620 24760 4672 24812
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 4804 24760 4856 24769
rect 2596 24624 2648 24676
rect 4528 24692 4580 24744
rect 5264 24760 5316 24812
rect 5908 24871 5960 24880
rect 5908 24837 5917 24871
rect 5917 24837 5951 24871
rect 5951 24837 5960 24871
rect 5908 24828 5960 24837
rect 5540 24803 5592 24812
rect 5540 24769 5549 24803
rect 5549 24769 5583 24803
rect 5583 24769 5592 24803
rect 5540 24760 5592 24769
rect 6920 24828 6972 24880
rect 7656 24828 7708 24880
rect 6276 24760 6328 24812
rect 5540 24624 5592 24676
rect 5908 24692 5960 24744
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 7196 24803 7248 24812
rect 7196 24769 7203 24803
rect 7203 24769 7248 24803
rect 7196 24760 7248 24769
rect 7932 24760 7984 24812
rect 7748 24692 7800 24744
rect 8208 24760 8260 24812
rect 9680 24828 9732 24880
rect 10968 24896 11020 24948
rect 11244 24896 11296 24948
rect 11704 24896 11756 24948
rect 12072 24896 12124 24948
rect 12624 24896 12676 24948
rect 13636 24896 13688 24948
rect 14280 24896 14332 24948
rect 15936 24896 15988 24948
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8803 24803
rect 8803 24769 8812 24803
rect 8760 24760 8812 24769
rect 9036 24760 9088 24812
rect 9128 24803 9180 24812
rect 9128 24769 9137 24803
rect 9137 24769 9171 24803
rect 9171 24769 9180 24803
rect 9128 24760 9180 24769
rect 9312 24760 9364 24812
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 9864 24760 9916 24812
rect 10876 24760 10928 24812
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 10968 24760 11020 24769
rect 11152 24692 11204 24744
rect 11336 24803 11388 24812
rect 11336 24769 11345 24803
rect 11345 24769 11379 24803
rect 11379 24769 11388 24803
rect 11336 24760 11388 24769
rect 11704 24760 11756 24812
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 10508 24624 10560 24676
rect 14188 24828 14240 24880
rect 15384 24828 15436 24880
rect 16212 24896 16264 24948
rect 16304 24896 16356 24948
rect 12256 24760 12308 24812
rect 13176 24803 13228 24812
rect 13176 24769 13185 24803
rect 13185 24769 13219 24803
rect 13219 24769 13228 24803
rect 13176 24760 13228 24769
rect 13452 24760 13504 24812
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 13912 24760 13964 24812
rect 14464 24760 14516 24812
rect 14280 24692 14332 24744
rect 14188 24624 14240 24676
rect 15292 24624 15344 24676
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 19248 24896 19300 24948
rect 16396 24828 16448 24880
rect 16764 24760 16816 24812
rect 16856 24760 16908 24812
rect 17316 24760 17368 24812
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 16580 24692 16632 24744
rect 17592 24692 17644 24744
rect 2872 24556 2924 24608
rect 4712 24599 4764 24608
rect 4712 24565 4721 24599
rect 4721 24565 4755 24599
rect 4755 24565 4764 24599
rect 4712 24556 4764 24565
rect 6276 24556 6328 24608
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 7564 24556 7616 24608
rect 7932 24556 7984 24608
rect 9312 24556 9364 24608
rect 9772 24599 9824 24608
rect 9772 24565 9781 24599
rect 9781 24565 9815 24599
rect 9815 24565 9824 24599
rect 9772 24556 9824 24565
rect 9864 24556 9916 24608
rect 10692 24556 10744 24608
rect 11888 24556 11940 24608
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 13452 24556 13504 24608
rect 15752 24599 15804 24608
rect 15752 24565 15761 24599
rect 15761 24565 15795 24599
rect 15795 24565 15804 24599
rect 15752 24556 15804 24565
rect 16764 24667 16816 24676
rect 16764 24633 16773 24667
rect 16773 24633 16807 24667
rect 16807 24633 16816 24667
rect 16764 24624 16816 24633
rect 17500 24599 17552 24608
rect 17500 24565 17509 24599
rect 17509 24565 17543 24599
rect 17543 24565 17552 24599
rect 17500 24556 17552 24565
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 18328 24760 18380 24812
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 18604 24692 18656 24744
rect 19248 24760 19300 24812
rect 20812 24896 20864 24948
rect 21548 24896 21600 24948
rect 22744 24896 22796 24948
rect 20996 24828 21048 24880
rect 19064 24692 19116 24744
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 20076 24760 20128 24812
rect 19432 24624 19484 24676
rect 19800 24692 19852 24744
rect 20352 24760 20404 24812
rect 20536 24760 20588 24812
rect 20812 24803 20864 24812
rect 20812 24769 20821 24803
rect 20821 24769 20855 24803
rect 20855 24769 20864 24803
rect 20812 24760 20864 24769
rect 21364 24828 21416 24880
rect 21824 24871 21876 24880
rect 21456 24803 21508 24812
rect 21456 24769 21465 24803
rect 21465 24769 21499 24803
rect 21499 24769 21508 24803
rect 21456 24760 21508 24769
rect 21824 24837 21833 24871
rect 21833 24837 21867 24871
rect 21867 24837 21876 24871
rect 21824 24828 21876 24837
rect 22376 24828 22428 24880
rect 21916 24760 21968 24812
rect 23112 24828 23164 24880
rect 24492 24896 24544 24948
rect 24584 24896 24636 24948
rect 27528 24896 27580 24948
rect 18144 24556 18196 24608
rect 18880 24556 18932 24608
rect 20260 24667 20312 24676
rect 20260 24633 20269 24667
rect 20269 24633 20303 24667
rect 20303 24633 20312 24667
rect 20260 24624 20312 24633
rect 19892 24599 19944 24608
rect 19892 24565 19901 24599
rect 19901 24565 19935 24599
rect 19935 24565 19944 24599
rect 19892 24556 19944 24565
rect 20168 24556 20220 24608
rect 21364 24692 21416 24744
rect 20444 24667 20496 24676
rect 20444 24633 20453 24667
rect 20453 24633 20487 24667
rect 20487 24633 20496 24667
rect 20444 24624 20496 24633
rect 20628 24624 20680 24676
rect 20904 24624 20956 24676
rect 22836 24760 22888 24812
rect 23572 24760 23624 24812
rect 23756 24760 23808 24812
rect 24124 24871 24176 24880
rect 24124 24837 24159 24871
rect 24159 24837 24176 24871
rect 24124 24828 24176 24837
rect 24400 24760 24452 24812
rect 23204 24692 23256 24744
rect 24676 24871 24728 24880
rect 24676 24837 24685 24871
rect 24685 24837 24719 24871
rect 24719 24837 24728 24871
rect 24676 24828 24728 24837
rect 25044 24828 25096 24880
rect 25320 24828 25372 24880
rect 25596 24828 25648 24880
rect 27160 24828 27212 24880
rect 28264 24896 28316 24948
rect 28816 24896 28868 24948
rect 30104 24896 30156 24948
rect 32680 24896 32732 24948
rect 24584 24803 24636 24812
rect 24584 24769 24593 24803
rect 24593 24769 24627 24803
rect 24627 24769 24636 24803
rect 24584 24760 24636 24769
rect 25504 24760 25556 24812
rect 26332 24760 26384 24812
rect 27344 24760 27396 24812
rect 24492 24624 24544 24676
rect 24584 24624 24636 24676
rect 24860 24624 24912 24676
rect 25136 24692 25188 24744
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 28724 24828 28776 24880
rect 28172 24803 28224 24812
rect 28172 24769 28181 24803
rect 28181 24769 28215 24803
rect 28215 24769 28224 24803
rect 28172 24760 28224 24769
rect 28264 24760 28316 24812
rect 33876 24896 33928 24948
rect 21088 24556 21140 24608
rect 22376 24556 22428 24608
rect 22836 24599 22888 24608
rect 22836 24565 22845 24599
rect 22845 24565 22879 24599
rect 22879 24565 22888 24599
rect 22836 24556 22888 24565
rect 23020 24556 23072 24608
rect 23572 24599 23624 24608
rect 23572 24565 23581 24599
rect 23581 24565 23615 24599
rect 23615 24565 23624 24599
rect 23572 24556 23624 24565
rect 24308 24556 24360 24608
rect 24952 24556 25004 24608
rect 25320 24556 25372 24608
rect 25872 24556 25924 24608
rect 26608 24556 26660 24608
rect 27804 24556 27856 24608
rect 28448 24735 28500 24744
rect 28448 24701 28457 24735
rect 28457 24701 28491 24735
rect 28491 24701 28500 24735
rect 28448 24692 28500 24701
rect 28908 24760 28960 24812
rect 32220 24760 32272 24812
rect 32956 24760 33008 24812
rect 33600 24803 33652 24812
rect 33600 24769 33609 24803
rect 33609 24769 33643 24803
rect 33643 24769 33652 24803
rect 33600 24760 33652 24769
rect 36452 24760 36504 24812
rect 29092 24735 29144 24744
rect 29092 24701 29101 24735
rect 29101 24701 29135 24735
rect 29135 24701 29144 24735
rect 29092 24692 29144 24701
rect 28172 24624 28224 24676
rect 28264 24556 28316 24608
rect 28632 24624 28684 24676
rect 29000 24624 29052 24676
rect 28724 24599 28776 24608
rect 28724 24565 28733 24599
rect 28733 24565 28767 24599
rect 28767 24565 28776 24599
rect 28724 24556 28776 24565
rect 32404 24692 32456 24744
rect 31944 24599 31996 24608
rect 31944 24565 31953 24599
rect 31953 24565 31987 24599
rect 31987 24565 31996 24599
rect 31944 24556 31996 24565
rect 33784 24599 33836 24608
rect 33784 24565 33793 24599
rect 33793 24565 33827 24599
rect 33827 24565 33836 24599
rect 33784 24556 33836 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3056 24352 3108 24404
rect 3608 24352 3660 24404
rect 3884 24352 3936 24404
rect 4528 24284 4580 24336
rect 4988 24352 5040 24404
rect 1216 24216 1268 24268
rect 2780 24216 2832 24268
rect 3516 24259 3568 24268
rect 3516 24225 3525 24259
rect 3525 24225 3559 24259
rect 3559 24225 3568 24259
rect 3516 24216 3568 24225
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 3884 24148 3936 24200
rect 4068 24148 4120 24200
rect 4712 24216 4764 24268
rect 4988 24148 5040 24200
rect 5080 24148 5132 24200
rect 5264 24148 5316 24200
rect 6920 24352 6972 24404
rect 7012 24352 7064 24404
rect 9128 24352 9180 24404
rect 3056 24080 3108 24132
rect 4068 24012 4120 24064
rect 5356 24123 5408 24132
rect 5356 24089 5365 24123
rect 5365 24089 5399 24123
rect 5399 24089 5408 24123
rect 5356 24080 5408 24089
rect 5632 24012 5684 24064
rect 5908 24148 5960 24200
rect 6092 24191 6144 24200
rect 6092 24157 6102 24191
rect 6102 24157 6136 24191
rect 6136 24157 6144 24191
rect 6092 24148 6144 24157
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 6828 24284 6880 24336
rect 7932 24284 7984 24336
rect 8668 24284 8720 24336
rect 6644 24148 6696 24200
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 6828 24080 6880 24132
rect 6920 24080 6972 24132
rect 7104 24012 7156 24064
rect 7932 24191 7984 24200
rect 7932 24157 7941 24191
rect 7941 24157 7975 24191
rect 7975 24157 7984 24191
rect 7932 24148 7984 24157
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 8208 24191 8260 24200
rect 8208 24157 8218 24191
rect 8218 24157 8252 24191
rect 8252 24157 8260 24191
rect 8208 24148 8260 24157
rect 7380 24123 7432 24132
rect 7380 24089 7389 24123
rect 7389 24089 7423 24123
rect 7423 24089 7432 24123
rect 7380 24080 7432 24089
rect 8392 24123 8444 24132
rect 8392 24089 8401 24123
rect 8401 24089 8435 24123
rect 8435 24089 8444 24123
rect 8392 24080 8444 24089
rect 8484 24123 8536 24132
rect 8484 24089 8493 24123
rect 8493 24089 8527 24123
rect 8527 24089 8536 24123
rect 8484 24080 8536 24089
rect 8760 24080 8812 24132
rect 7564 24012 7616 24064
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 9036 24191 9088 24200
rect 9036 24157 9046 24191
rect 9046 24157 9080 24191
rect 9080 24157 9088 24191
rect 10232 24284 10284 24336
rect 10508 24327 10560 24336
rect 10508 24293 10517 24327
rect 10517 24293 10551 24327
rect 10551 24293 10560 24327
rect 10508 24284 10560 24293
rect 9312 24216 9364 24268
rect 11336 24352 11388 24404
rect 11612 24352 11664 24404
rect 11980 24352 12032 24404
rect 13728 24352 13780 24404
rect 14096 24352 14148 24404
rect 15476 24352 15528 24404
rect 16580 24352 16632 24404
rect 17960 24352 18012 24404
rect 18788 24352 18840 24404
rect 9036 24148 9088 24157
rect 9680 24148 9732 24200
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 10968 24191 11020 24200
rect 10968 24157 10977 24191
rect 10977 24157 11011 24191
rect 11011 24157 11020 24191
rect 10968 24148 11020 24157
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 11244 24148 11296 24200
rect 11888 24216 11940 24268
rect 11612 24191 11664 24200
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 12716 24259 12768 24268
rect 12716 24225 12725 24259
rect 12725 24225 12759 24259
rect 12759 24225 12768 24259
rect 12716 24216 12768 24225
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 13360 24284 13412 24336
rect 13820 24216 13872 24268
rect 9312 24123 9364 24132
rect 9312 24089 9321 24123
rect 9321 24089 9355 24123
rect 9355 24089 9364 24123
rect 9312 24080 9364 24089
rect 9496 24012 9548 24064
rect 12072 24080 12124 24132
rect 13728 24191 13780 24200
rect 13728 24157 13737 24191
rect 13737 24157 13771 24191
rect 13771 24157 13780 24191
rect 13728 24148 13780 24157
rect 13912 24148 13964 24200
rect 13452 24080 13504 24132
rect 14372 24284 14424 24336
rect 14096 24216 14148 24268
rect 15384 24284 15436 24336
rect 15568 24284 15620 24336
rect 16672 24284 16724 24336
rect 17224 24284 17276 24336
rect 17316 24284 17368 24336
rect 18052 24216 18104 24268
rect 18512 24284 18564 24336
rect 19892 24352 19944 24404
rect 18972 24284 19024 24336
rect 20076 24284 20128 24336
rect 20168 24284 20220 24336
rect 21640 24352 21692 24404
rect 21732 24352 21784 24404
rect 20260 24216 20312 24268
rect 14188 24012 14240 24064
rect 14556 24080 14608 24132
rect 15292 24080 15344 24132
rect 15660 24148 15712 24200
rect 16120 24191 16172 24200
rect 16120 24157 16129 24191
rect 16129 24157 16163 24191
rect 16163 24157 16172 24191
rect 16120 24148 16172 24157
rect 16488 24191 16540 24200
rect 16488 24157 16497 24191
rect 16497 24157 16531 24191
rect 16531 24157 16540 24191
rect 16488 24148 16540 24157
rect 16948 24148 17000 24200
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 17960 24148 18012 24200
rect 17316 24080 17368 24132
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 18880 24148 18932 24200
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 19708 24148 19760 24200
rect 19800 24148 19852 24200
rect 15568 24012 15620 24064
rect 15936 24055 15988 24064
rect 15936 24021 15945 24055
rect 15945 24021 15979 24055
rect 15979 24021 15988 24055
rect 15936 24012 15988 24021
rect 16304 24012 16356 24064
rect 17776 24012 17828 24064
rect 18328 24012 18380 24064
rect 19984 24080 20036 24132
rect 20444 24080 20496 24132
rect 19800 24012 19852 24064
rect 20076 24012 20128 24064
rect 20168 24012 20220 24064
rect 20812 24148 20864 24200
rect 21088 24148 21140 24200
rect 21180 24148 21232 24200
rect 21548 24148 21600 24200
rect 22100 24191 22152 24200
rect 22100 24157 22109 24191
rect 22109 24157 22143 24191
rect 22143 24157 22152 24191
rect 22100 24148 22152 24157
rect 23204 24352 23256 24404
rect 24032 24352 24084 24404
rect 24768 24352 24820 24404
rect 25044 24352 25096 24404
rect 25412 24352 25464 24404
rect 26332 24352 26384 24404
rect 27160 24352 27212 24404
rect 27528 24352 27580 24404
rect 27712 24352 27764 24404
rect 29000 24352 29052 24404
rect 30196 24352 30248 24404
rect 23756 24284 23808 24336
rect 23296 24216 23348 24268
rect 23480 24259 23532 24268
rect 23480 24225 23489 24259
rect 23489 24225 23523 24259
rect 23523 24225 23532 24259
rect 23480 24216 23532 24225
rect 22376 24191 22428 24200
rect 22376 24157 22385 24191
rect 22385 24157 22419 24191
rect 22419 24157 22428 24191
rect 22376 24148 22428 24157
rect 24032 24148 24084 24200
rect 25504 24216 25556 24268
rect 24768 24191 24820 24200
rect 24768 24157 24777 24191
rect 24777 24157 24811 24191
rect 24811 24157 24820 24191
rect 24768 24148 24820 24157
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 25596 24148 25648 24200
rect 25872 24216 25924 24268
rect 23388 24123 23440 24132
rect 23388 24089 23397 24123
rect 23397 24089 23431 24123
rect 23431 24089 23440 24123
rect 23388 24080 23440 24089
rect 24308 24080 24360 24132
rect 20904 24012 20956 24064
rect 20996 24012 21048 24064
rect 21456 24012 21508 24064
rect 23480 24012 23532 24064
rect 24124 24012 24176 24064
rect 24400 24055 24452 24064
rect 24400 24021 24409 24055
rect 24409 24021 24443 24055
rect 24443 24021 24452 24055
rect 24400 24012 24452 24021
rect 24584 24080 24636 24132
rect 25872 24123 25924 24132
rect 25872 24089 25881 24123
rect 25881 24089 25915 24123
rect 25915 24089 25924 24123
rect 25872 24080 25924 24089
rect 26148 24148 26200 24200
rect 26700 24284 26752 24336
rect 26884 24216 26936 24268
rect 27804 24284 27856 24336
rect 28724 24284 28776 24336
rect 25228 24012 25280 24064
rect 25688 24012 25740 24064
rect 26148 24012 26200 24064
rect 26286 24012 26338 24064
rect 26976 24080 27028 24132
rect 27804 24191 27856 24200
rect 27804 24157 27813 24191
rect 27813 24157 27847 24191
rect 27847 24157 27856 24191
rect 27804 24148 27856 24157
rect 31944 24352 31996 24404
rect 33784 24352 33836 24404
rect 32128 24216 32180 24268
rect 27528 24080 27580 24132
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 27160 24012 27212 24064
rect 27896 24080 27948 24132
rect 29092 24080 29144 24132
rect 29460 24080 29512 24132
rect 27988 24055 28040 24064
rect 27988 24021 27997 24055
rect 27997 24021 28031 24055
rect 28031 24021 28040 24055
rect 27988 24012 28040 24021
rect 32312 24055 32364 24064
rect 32312 24021 32321 24055
rect 32321 24021 32355 24055
rect 32355 24021 32364 24055
rect 32312 24012 32364 24021
rect 33784 24055 33836 24064
rect 33784 24021 33793 24055
rect 33793 24021 33827 24055
rect 33827 24021 33836 24055
rect 33784 24012 33836 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4068 23808 4120 23860
rect 4712 23808 4764 23860
rect 5540 23851 5592 23860
rect 5540 23817 5549 23851
rect 5549 23817 5583 23851
rect 5583 23817 5592 23851
rect 5540 23808 5592 23817
rect 5724 23808 5776 23860
rect 6828 23808 6880 23860
rect 7656 23808 7708 23860
rect 8668 23808 8720 23860
rect 8944 23808 8996 23860
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 9864 23808 9916 23860
rect 13084 23808 13136 23860
rect 13452 23808 13504 23860
rect 14004 23808 14056 23860
rect 2136 23672 2188 23724
rect 3148 23672 3200 23724
rect 3332 23672 3384 23724
rect 3792 23672 3844 23724
rect 1768 23604 1820 23656
rect 2044 23647 2096 23656
rect 2044 23613 2053 23647
rect 2053 23613 2087 23647
rect 2087 23613 2096 23647
rect 2044 23604 2096 23613
rect 4160 23647 4212 23656
rect 3240 23536 3292 23588
rect 4160 23613 4169 23647
rect 4169 23613 4203 23647
rect 4203 23613 4212 23647
rect 4160 23604 4212 23613
rect 5080 23672 5132 23724
rect 5172 23672 5224 23724
rect 4804 23604 4856 23656
rect 5816 23672 5868 23724
rect 6000 23672 6052 23724
rect 7012 23740 7064 23792
rect 6736 23672 6788 23724
rect 9496 23740 9548 23792
rect 11980 23740 12032 23792
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 11244 23672 11296 23724
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 11888 23672 11940 23724
rect 12624 23715 12676 23724
rect 12624 23681 12633 23715
rect 12633 23681 12667 23715
rect 12667 23681 12676 23715
rect 12624 23672 12676 23681
rect 12992 23672 13044 23724
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 7288 23604 7340 23656
rect 7472 23604 7524 23656
rect 7840 23604 7892 23656
rect 9036 23604 9088 23656
rect 9220 23604 9272 23656
rect 10508 23604 10560 23656
rect 5264 23536 5316 23588
rect 9128 23536 9180 23588
rect 10876 23536 10928 23588
rect 3332 23468 3384 23520
rect 4068 23468 4120 23520
rect 5172 23468 5224 23520
rect 5632 23468 5684 23520
rect 5816 23511 5868 23520
rect 5816 23477 5825 23511
rect 5825 23477 5859 23511
rect 5859 23477 5868 23511
rect 5816 23468 5868 23477
rect 6828 23468 6880 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 7840 23511 7892 23520
rect 7840 23477 7849 23511
rect 7849 23477 7883 23511
rect 7883 23477 7892 23511
rect 7840 23468 7892 23477
rect 8208 23511 8260 23520
rect 8208 23477 8217 23511
rect 8217 23477 8251 23511
rect 8251 23477 8260 23511
rect 8208 23468 8260 23477
rect 9956 23468 10008 23520
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 10692 23468 10744 23520
rect 11612 23468 11664 23520
rect 12256 23536 12308 23588
rect 14188 23672 14240 23724
rect 14740 23808 14792 23860
rect 15200 23851 15252 23860
rect 15200 23817 15209 23851
rect 15209 23817 15243 23851
rect 15243 23817 15252 23851
rect 15200 23808 15252 23817
rect 14556 23740 14608 23792
rect 14832 23740 14884 23792
rect 15292 23715 15344 23724
rect 15292 23681 15301 23715
rect 15301 23681 15335 23715
rect 15335 23681 15344 23715
rect 15292 23672 15344 23681
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 14280 23604 14332 23656
rect 15016 23604 15068 23656
rect 15200 23604 15252 23656
rect 17500 23740 17552 23792
rect 17960 23740 18012 23792
rect 19800 23808 19852 23860
rect 16764 23672 16816 23724
rect 17776 23672 17828 23724
rect 18512 23740 18564 23792
rect 20628 23808 20680 23860
rect 20720 23808 20772 23860
rect 21088 23808 21140 23860
rect 21272 23808 21324 23860
rect 21364 23808 21416 23860
rect 18972 23715 19024 23724
rect 18972 23681 18989 23715
rect 18989 23681 19024 23715
rect 18972 23672 19024 23681
rect 19248 23672 19300 23724
rect 19340 23715 19392 23724
rect 19340 23681 19349 23715
rect 19349 23681 19383 23715
rect 19383 23681 19392 23715
rect 19340 23672 19392 23681
rect 17132 23536 17184 23588
rect 17592 23604 17644 23656
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 18144 23536 18196 23588
rect 18420 23536 18472 23588
rect 12624 23468 12676 23520
rect 14004 23468 14056 23520
rect 15568 23468 15620 23520
rect 16304 23468 16356 23520
rect 16764 23511 16816 23520
rect 16764 23477 16773 23511
rect 16773 23477 16807 23511
rect 16807 23477 16816 23511
rect 16764 23468 16816 23477
rect 18052 23511 18104 23520
rect 18052 23477 18061 23511
rect 18061 23477 18095 23511
rect 18095 23477 18104 23511
rect 18052 23468 18104 23477
rect 18880 23511 18932 23520
rect 18880 23477 18889 23511
rect 18889 23477 18923 23511
rect 18923 23477 18932 23511
rect 18880 23468 18932 23477
rect 19524 23579 19576 23588
rect 19524 23545 19533 23579
rect 19533 23545 19567 23579
rect 19567 23545 19576 23579
rect 20076 23740 20128 23792
rect 21640 23808 21692 23860
rect 22008 23808 22060 23860
rect 20444 23715 20496 23724
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 20444 23672 20496 23681
rect 20536 23672 20588 23724
rect 20720 23672 20772 23724
rect 19984 23604 20036 23656
rect 20996 23604 21048 23656
rect 21456 23672 21508 23724
rect 22100 23740 22152 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 23020 23740 23072 23792
rect 23296 23783 23348 23792
rect 23296 23749 23305 23783
rect 23305 23749 23339 23783
rect 23339 23749 23348 23783
rect 23296 23740 23348 23749
rect 23388 23783 23440 23792
rect 23388 23749 23397 23783
rect 23397 23749 23431 23783
rect 23431 23749 23440 23783
rect 23388 23740 23440 23749
rect 23756 23808 23808 23860
rect 25320 23808 25372 23860
rect 25504 23851 25556 23860
rect 25504 23817 25513 23851
rect 25513 23817 25547 23851
rect 25547 23817 25556 23851
rect 25504 23808 25556 23817
rect 25872 23808 25924 23860
rect 22560 23672 22612 23724
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 23572 23672 23624 23724
rect 25044 23740 25096 23792
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 24124 23715 24176 23724
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 24768 23672 24820 23724
rect 24860 23672 24912 23724
rect 19524 23536 19576 23545
rect 20076 23536 20128 23588
rect 20260 23536 20312 23588
rect 21364 23536 21416 23588
rect 21640 23536 21692 23588
rect 22284 23536 22336 23588
rect 22468 23536 22520 23588
rect 25044 23536 25096 23588
rect 20352 23468 20404 23520
rect 21272 23468 21324 23520
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 27896 23808 27948 23860
rect 29000 23808 29052 23860
rect 30012 23808 30064 23860
rect 25964 23783 26016 23792
rect 25964 23749 25973 23783
rect 25973 23749 26007 23783
rect 26007 23749 26016 23783
rect 25964 23740 26016 23749
rect 27068 23740 27120 23792
rect 27436 23740 27488 23792
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27620 23715 27672 23724
rect 27620 23681 27629 23715
rect 27629 23681 27663 23715
rect 27663 23681 27672 23715
rect 27620 23672 27672 23681
rect 27896 23715 27948 23724
rect 27896 23681 27905 23715
rect 27905 23681 27939 23715
rect 27939 23681 27948 23715
rect 27896 23672 27948 23681
rect 29552 23740 29604 23792
rect 31668 23783 31720 23792
rect 31668 23749 31677 23783
rect 31677 23749 31711 23783
rect 31711 23749 31720 23783
rect 31668 23740 31720 23749
rect 25964 23536 26016 23588
rect 26056 23536 26108 23588
rect 27804 23604 27856 23656
rect 32312 23672 32364 23724
rect 33784 23808 33836 23860
rect 29460 23647 29512 23656
rect 29460 23613 29469 23647
rect 29469 23613 29503 23647
rect 29503 23613 29512 23647
rect 29460 23604 29512 23613
rect 23756 23468 23808 23520
rect 25136 23468 25188 23520
rect 25320 23511 25372 23520
rect 25320 23477 25329 23511
rect 25329 23477 25363 23511
rect 25363 23477 25372 23511
rect 25320 23468 25372 23477
rect 25780 23468 25832 23520
rect 27528 23511 27580 23520
rect 27528 23477 27537 23511
rect 27537 23477 27571 23511
rect 27571 23477 27580 23511
rect 27528 23468 27580 23477
rect 28172 23511 28224 23520
rect 28172 23477 28181 23511
rect 28181 23477 28215 23511
rect 28215 23477 28224 23511
rect 28172 23468 28224 23477
rect 33140 23511 33192 23520
rect 33140 23477 33149 23511
rect 33149 23477 33183 23511
rect 33183 23477 33192 23511
rect 33140 23468 33192 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2872 23307 2924 23316
rect 2872 23273 2881 23307
rect 2881 23273 2915 23307
rect 2915 23273 2924 23307
rect 2872 23264 2924 23273
rect 3332 23264 3384 23316
rect 7104 23264 7156 23316
rect 7196 23264 7248 23316
rect 7932 23264 7984 23316
rect 1216 23128 1268 23180
rect 6368 23239 6420 23248
rect 6368 23205 6377 23239
rect 6377 23205 6411 23239
rect 6411 23205 6420 23239
rect 6368 23196 6420 23205
rect 6736 23196 6788 23248
rect 3608 23128 3660 23180
rect 3240 23103 3292 23112
rect 3240 23069 3249 23103
rect 3249 23069 3283 23103
rect 3283 23069 3292 23103
rect 3240 23060 3292 23069
rect 2136 22992 2188 23044
rect 4068 23060 4120 23112
rect 4620 23128 4672 23180
rect 3792 23035 3844 23044
rect 3792 23001 3801 23035
rect 3801 23001 3835 23035
rect 3835 23001 3844 23035
rect 3792 22992 3844 23001
rect 4712 23103 4764 23112
rect 4712 23069 4726 23103
rect 4726 23069 4760 23103
rect 4760 23069 4764 23103
rect 4712 23060 4764 23069
rect 1584 22924 1636 22976
rect 3056 22924 3108 22976
rect 3240 22924 3292 22976
rect 3516 22924 3568 22976
rect 4620 23035 4672 23044
rect 4620 23001 4629 23035
rect 4629 23001 4663 23035
rect 4663 23001 4672 23035
rect 4620 22992 4672 23001
rect 4252 22924 4304 22976
rect 5908 23128 5960 23180
rect 8668 23196 8720 23248
rect 8852 23264 8904 23316
rect 9680 23264 9732 23316
rect 10876 23264 10928 23316
rect 11336 23264 11388 23316
rect 10692 23196 10744 23248
rect 5816 23103 5868 23112
rect 5816 23069 5826 23103
rect 5826 23069 5860 23103
rect 5860 23069 5868 23103
rect 5816 23060 5868 23069
rect 5172 22924 5224 22976
rect 5356 22924 5408 22976
rect 5632 22992 5684 23044
rect 6736 23060 6788 23112
rect 7104 23060 7156 23112
rect 7380 23103 7432 23112
rect 7380 23069 7394 23103
rect 7394 23069 7428 23103
rect 7428 23069 7432 23103
rect 7380 23060 7432 23069
rect 10600 23060 10652 23112
rect 10324 22992 10376 23044
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11428 23128 11480 23180
rect 11888 23196 11940 23248
rect 11060 23060 11112 23069
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 14832 23264 14884 23316
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 17040 23307 17092 23316
rect 17040 23273 17049 23307
rect 17049 23273 17083 23307
rect 17083 23273 17092 23307
rect 17040 23264 17092 23273
rect 12440 23060 12492 23112
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 13084 23060 13136 23112
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 14740 23196 14792 23248
rect 17224 23264 17276 23316
rect 17316 23196 17368 23248
rect 18328 23264 18380 23316
rect 18972 23264 19024 23316
rect 19248 23264 19300 23316
rect 19892 23307 19944 23316
rect 19892 23273 19901 23307
rect 19901 23273 19935 23307
rect 19935 23273 19944 23307
rect 19892 23264 19944 23273
rect 20076 23264 20128 23316
rect 21364 23264 21416 23316
rect 15108 23060 15160 23112
rect 16764 23060 16816 23112
rect 17776 23103 17828 23112
rect 17776 23069 17785 23103
rect 17785 23069 17819 23103
rect 17819 23069 17828 23103
rect 17776 23060 17828 23069
rect 6368 22924 6420 22976
rect 6552 22924 6604 22976
rect 6920 22924 6972 22976
rect 7564 22967 7616 22976
rect 7564 22933 7573 22967
rect 7573 22933 7607 22967
rect 7607 22933 7616 22967
rect 7564 22924 7616 22933
rect 7656 22924 7708 22976
rect 8116 22924 8168 22976
rect 8208 22924 8260 22976
rect 10784 22924 10836 22976
rect 11060 22924 11112 22976
rect 12072 22924 12124 22976
rect 12256 23035 12308 23044
rect 12256 23001 12262 23035
rect 12262 23001 12296 23035
rect 12296 23001 12308 23035
rect 12256 22992 12308 23001
rect 12532 22967 12584 22976
rect 12532 22933 12541 22967
rect 12541 22933 12575 22967
rect 12575 22933 12584 22967
rect 12532 22924 12584 22933
rect 12808 23035 12860 23044
rect 12808 23001 12817 23035
rect 12817 23001 12851 23035
rect 12851 23001 12860 23035
rect 12808 22992 12860 23001
rect 12900 23035 12952 23044
rect 12900 23001 12909 23035
rect 12909 23001 12943 23035
rect 12943 23001 12952 23035
rect 12900 22992 12952 23001
rect 13360 22992 13412 23044
rect 14004 22992 14056 23044
rect 16580 23035 16632 23044
rect 16580 23001 16589 23035
rect 16589 23001 16623 23035
rect 16623 23001 16632 23035
rect 16580 22992 16632 23001
rect 17040 22992 17092 23044
rect 19616 23196 19668 23248
rect 20444 23196 20496 23248
rect 20720 23196 20772 23248
rect 18420 23103 18472 23112
rect 18420 23069 18441 23103
rect 18441 23069 18472 23103
rect 18420 23060 18472 23069
rect 18328 23035 18380 23044
rect 18328 23001 18337 23035
rect 18337 23001 18371 23035
rect 18371 23001 18380 23035
rect 18328 22992 18380 23001
rect 18788 23103 18840 23112
rect 18788 23069 18797 23103
rect 18797 23069 18831 23103
rect 18831 23069 18840 23103
rect 18788 23060 18840 23069
rect 19340 23103 19392 23112
rect 19340 23069 19349 23103
rect 19349 23069 19383 23103
rect 19383 23069 19392 23103
rect 19340 23060 19392 23069
rect 19892 23060 19944 23112
rect 20168 23103 20220 23112
rect 20168 23069 20177 23103
rect 20177 23069 20211 23103
rect 20211 23069 20220 23103
rect 20168 23060 20220 23069
rect 20536 23060 20588 23112
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 20904 23060 20956 23112
rect 21548 23196 21600 23248
rect 21916 23264 21968 23316
rect 22928 23264 22980 23316
rect 23296 23264 23348 23316
rect 23940 23264 23992 23316
rect 25136 23307 25188 23316
rect 25136 23273 25145 23307
rect 25145 23273 25179 23307
rect 25179 23273 25188 23307
rect 25136 23264 25188 23273
rect 27344 23264 27396 23316
rect 28080 23264 28132 23316
rect 32404 23264 32456 23316
rect 33140 23264 33192 23316
rect 33600 23264 33652 23316
rect 21180 23060 21232 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 22284 23128 22336 23180
rect 21916 23060 21968 23112
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 25412 23196 25464 23248
rect 26056 23128 26108 23180
rect 15200 22924 15252 22976
rect 15568 22924 15620 22976
rect 17316 22924 17368 22976
rect 17500 22924 17552 22976
rect 18052 22924 18104 22976
rect 20536 22924 20588 22976
rect 21272 22924 21324 22976
rect 21732 22924 21784 22976
rect 22008 22924 22060 22976
rect 23480 23060 23532 23112
rect 25688 23060 25740 23112
rect 23112 22924 23164 22976
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 23572 22924 23624 22976
rect 24124 22992 24176 23044
rect 24768 22992 24820 23044
rect 24860 23035 24912 23044
rect 24860 23001 24869 23035
rect 24869 23001 24903 23035
rect 24903 23001 24912 23035
rect 24860 22992 24912 23001
rect 24952 22992 25004 23044
rect 25872 23103 25924 23112
rect 25872 23069 25882 23103
rect 25882 23069 25916 23103
rect 25916 23069 25924 23103
rect 25872 23060 25924 23069
rect 26424 23060 26476 23112
rect 26608 23060 26660 23112
rect 26700 23103 26752 23112
rect 26700 23069 26709 23103
rect 26709 23069 26743 23103
rect 26743 23069 26752 23103
rect 26700 23060 26752 23069
rect 26976 23060 27028 23112
rect 27436 23060 27488 23112
rect 27804 23060 27856 23112
rect 28540 23128 28592 23180
rect 32312 23128 32364 23180
rect 28264 23060 28316 23112
rect 25136 22924 25188 22976
rect 26240 22924 26292 22976
rect 26424 22967 26476 22976
rect 26424 22933 26433 22967
rect 26433 22933 26467 22967
rect 26467 22933 26476 22967
rect 26424 22924 26476 22933
rect 27160 22924 27212 22976
rect 27712 22924 27764 22976
rect 28356 22924 28408 22976
rect 28448 22924 28500 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3148 22720 3200 22772
rect 3884 22720 3936 22772
rect 3976 22652 4028 22704
rect 3884 22584 3936 22636
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 3700 22559 3752 22568
rect 3700 22525 3709 22559
rect 3709 22525 3743 22559
rect 3743 22525 3752 22559
rect 3700 22516 3752 22525
rect 6552 22720 6604 22772
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 5080 22584 5132 22636
rect 5540 22627 5592 22636
rect 5540 22593 5549 22627
rect 5549 22593 5583 22627
rect 5583 22593 5592 22627
rect 5540 22584 5592 22593
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 5724 22584 5776 22636
rect 5908 22627 5960 22636
rect 5908 22593 5917 22627
rect 5917 22593 5951 22627
rect 5951 22593 5960 22627
rect 5908 22584 5960 22593
rect 6276 22584 6328 22636
rect 6644 22652 6696 22704
rect 7196 22695 7248 22704
rect 7196 22661 7205 22695
rect 7205 22661 7239 22695
rect 7239 22661 7248 22695
rect 7196 22652 7248 22661
rect 6828 22584 6880 22636
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 7104 22584 7156 22636
rect 6644 22516 6696 22568
rect 7380 22584 7432 22636
rect 7932 22695 7984 22704
rect 7932 22661 7941 22695
rect 7941 22661 7975 22695
rect 7975 22661 7984 22695
rect 7932 22652 7984 22661
rect 8024 22695 8076 22704
rect 8024 22661 8033 22695
rect 8033 22661 8067 22695
rect 8067 22661 8076 22695
rect 8024 22652 8076 22661
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 10048 22652 10100 22704
rect 10324 22763 10376 22772
rect 10324 22729 10333 22763
rect 10333 22729 10367 22763
rect 10367 22729 10376 22763
rect 10324 22720 10376 22729
rect 10876 22720 10928 22772
rect 11060 22720 11112 22772
rect 12348 22720 12400 22772
rect 13268 22720 13320 22772
rect 13820 22720 13872 22772
rect 15108 22720 15160 22772
rect 15384 22720 15436 22772
rect 15844 22720 15896 22772
rect 16120 22720 16172 22772
rect 18052 22720 18104 22772
rect 19064 22720 19116 22772
rect 19248 22720 19300 22772
rect 19524 22720 19576 22772
rect 20168 22720 20220 22772
rect 8484 22584 8536 22636
rect 8852 22584 8904 22636
rect 3148 22448 3200 22500
rect 4068 22448 4120 22500
rect 1768 22380 1820 22432
rect 2412 22380 2464 22432
rect 4896 22380 4948 22432
rect 5448 22448 5500 22500
rect 6000 22448 6052 22500
rect 6828 22491 6880 22500
rect 6828 22457 6837 22491
rect 6837 22457 6871 22491
rect 6871 22457 6880 22491
rect 6828 22448 6880 22457
rect 7840 22448 7892 22500
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9128 22584 9180 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9496 22584 9548 22636
rect 11244 22652 11296 22704
rect 12808 22652 12860 22704
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 10232 22448 10284 22500
rect 10600 22448 10652 22500
rect 6092 22380 6144 22432
rect 6736 22380 6788 22432
rect 7012 22380 7064 22432
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 8300 22423 8352 22432
rect 8300 22389 8309 22423
rect 8309 22389 8343 22423
rect 8343 22389 8352 22423
rect 8300 22380 8352 22389
rect 9128 22380 9180 22432
rect 9680 22380 9732 22432
rect 9956 22380 10008 22432
rect 10324 22380 10376 22432
rect 11152 22584 11204 22636
rect 10968 22516 11020 22568
rect 11612 22516 11664 22568
rect 12348 22448 12400 22500
rect 12716 22559 12768 22568
rect 12716 22525 12725 22559
rect 12725 22525 12759 22559
rect 12759 22525 12768 22559
rect 12716 22516 12768 22525
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 17960 22652 18012 22704
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 15016 22584 15068 22636
rect 13636 22516 13688 22568
rect 15384 22516 15436 22568
rect 15568 22584 15620 22636
rect 16396 22584 16448 22636
rect 17224 22584 17276 22636
rect 17684 22584 17736 22636
rect 19616 22652 19668 22704
rect 16764 22516 16816 22568
rect 17316 22516 17368 22568
rect 18420 22584 18472 22636
rect 18512 22516 18564 22568
rect 13084 22448 13136 22500
rect 13360 22448 13412 22500
rect 11612 22380 11664 22432
rect 11796 22380 11848 22432
rect 16672 22448 16724 22500
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 19340 22584 19392 22636
rect 19432 22627 19484 22636
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 19524 22584 19576 22636
rect 19892 22584 19944 22636
rect 20720 22720 20772 22772
rect 21088 22720 21140 22772
rect 21456 22720 21508 22772
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 23480 22763 23532 22772
rect 23480 22729 23489 22763
rect 23489 22729 23523 22763
rect 23523 22729 23532 22763
rect 23480 22720 23532 22729
rect 24400 22720 24452 22772
rect 24584 22720 24636 22772
rect 20352 22627 20404 22636
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 20444 22584 20496 22636
rect 20628 22584 20680 22636
rect 21364 22652 21416 22704
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 21088 22584 21140 22593
rect 21180 22584 21232 22636
rect 21364 22516 21416 22568
rect 13912 22380 13964 22432
rect 14832 22380 14884 22432
rect 15476 22380 15528 22432
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 16580 22380 16632 22432
rect 17132 22380 17184 22432
rect 17592 22380 17644 22432
rect 17960 22380 18012 22432
rect 18420 22380 18472 22432
rect 18696 22423 18748 22432
rect 18696 22389 18705 22423
rect 18705 22389 18739 22423
rect 18739 22389 18748 22423
rect 18696 22380 18748 22389
rect 18788 22380 18840 22432
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 20904 22448 20956 22500
rect 21088 22491 21140 22500
rect 21088 22457 21097 22491
rect 21097 22457 21131 22491
rect 21131 22457 21140 22491
rect 21916 22652 21968 22704
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 21824 22516 21876 22568
rect 22284 22516 22336 22568
rect 22560 22584 22612 22636
rect 22744 22627 22796 22636
rect 22744 22593 22753 22627
rect 22753 22593 22787 22627
rect 22787 22593 22796 22627
rect 22744 22584 22796 22593
rect 21088 22448 21140 22457
rect 20260 22380 20312 22432
rect 20536 22380 20588 22432
rect 20720 22380 20772 22432
rect 22192 22448 22244 22500
rect 22928 22584 22980 22636
rect 23756 22584 23808 22636
rect 25136 22652 25188 22704
rect 26884 22652 26936 22704
rect 27436 22720 27488 22772
rect 27712 22652 27764 22704
rect 27896 22695 27948 22704
rect 27896 22661 27905 22695
rect 27905 22661 27939 22695
rect 27939 22661 27948 22695
rect 27896 22652 27948 22661
rect 21640 22380 21692 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 22652 22380 22704 22432
rect 23296 22516 23348 22568
rect 23480 22516 23532 22568
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 24492 22584 24544 22636
rect 24768 22627 24820 22636
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 23572 22448 23624 22500
rect 26240 22584 26292 22636
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 28080 22652 28132 22704
rect 28540 22763 28592 22772
rect 28540 22729 28549 22763
rect 28549 22729 28583 22763
rect 28583 22729 28592 22763
rect 28540 22720 28592 22729
rect 26608 22516 26660 22568
rect 28264 22627 28316 22636
rect 28264 22593 28273 22627
rect 28273 22593 28307 22627
rect 28307 22593 28316 22627
rect 28264 22584 28316 22593
rect 28356 22584 28408 22636
rect 28632 22584 28684 22636
rect 25872 22448 25924 22500
rect 24860 22380 24912 22432
rect 24952 22423 25004 22432
rect 24952 22389 24961 22423
rect 24961 22389 24995 22423
rect 24995 22389 25004 22423
rect 24952 22380 25004 22389
rect 25780 22423 25832 22432
rect 25780 22389 25789 22423
rect 25789 22389 25823 22423
rect 25823 22389 25832 22423
rect 25780 22380 25832 22389
rect 27988 22448 28040 22500
rect 26148 22380 26200 22432
rect 27436 22380 27488 22432
rect 27620 22380 27672 22432
rect 27896 22380 27948 22432
rect 28448 22380 28500 22432
rect 28632 22380 28684 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2872 22176 2924 22228
rect 1216 22040 1268 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 3700 22108 3752 22160
rect 3424 22040 3476 22092
rect 4712 22176 4764 22228
rect 5356 22219 5408 22228
rect 5356 22185 5365 22219
rect 5365 22185 5399 22219
rect 5399 22185 5408 22219
rect 5356 22176 5408 22185
rect 5632 22176 5684 22228
rect 4620 22108 4672 22160
rect 7932 22176 7984 22228
rect 8116 22176 8168 22228
rect 9404 22176 9456 22228
rect 9772 22176 9824 22228
rect 11152 22176 11204 22228
rect 11520 22176 11572 22228
rect 12348 22176 12400 22228
rect 5908 22108 5960 22160
rect 4344 22040 4396 22092
rect 5264 22040 5316 22092
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5356 21972 5408 22024
rect 5724 22040 5776 22092
rect 6276 22040 6328 22092
rect 6000 21972 6052 22024
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6460 22040 6512 22092
rect 6736 22151 6788 22160
rect 6736 22117 6745 22151
rect 6745 22117 6779 22151
rect 6779 22117 6788 22151
rect 6736 22108 6788 22117
rect 7104 22108 7156 22160
rect 8852 22108 8904 22160
rect 4436 21904 4488 21956
rect 4988 21947 5040 21956
rect 4988 21913 4997 21947
rect 4997 21913 5031 21947
rect 5031 21913 5040 21947
rect 4988 21904 5040 21913
rect 5264 21904 5316 21956
rect 5448 21836 5500 21888
rect 5816 21836 5868 21888
rect 6184 21836 6236 21888
rect 7380 21972 7432 22024
rect 8024 22040 8076 22092
rect 8300 22040 8352 22092
rect 9128 22040 9180 22092
rect 9496 22040 9548 22092
rect 6828 21947 6880 21956
rect 6828 21913 6837 21947
rect 6837 21913 6871 21947
rect 6871 21913 6880 21947
rect 6828 21904 6880 21913
rect 7104 21904 7156 21956
rect 7564 21947 7616 21956
rect 7564 21913 7573 21947
rect 7573 21913 7607 21947
rect 7607 21913 7616 21947
rect 7564 21904 7616 21913
rect 8392 21972 8444 22024
rect 8484 21972 8536 22024
rect 7932 21904 7984 21956
rect 8116 21947 8168 21956
rect 8116 21913 8125 21947
rect 8125 21913 8159 21947
rect 8159 21913 8168 21947
rect 8116 21904 8168 21913
rect 8668 21972 8720 22024
rect 9036 21972 9088 22024
rect 9404 22015 9456 22024
rect 9404 21981 9414 22015
rect 9414 21981 9448 22015
rect 9448 21981 9456 22015
rect 9956 22151 10008 22160
rect 9956 22117 9965 22151
rect 9965 22117 9999 22151
rect 9999 22117 10008 22151
rect 9956 22108 10008 22117
rect 10968 22108 11020 22160
rect 10600 22040 10652 22092
rect 11244 22040 11296 22092
rect 11796 22040 11848 22092
rect 11980 22108 12032 22160
rect 9404 21972 9456 21981
rect 6920 21836 6972 21888
rect 7840 21836 7892 21888
rect 8208 21836 8260 21888
rect 8852 21836 8904 21888
rect 9496 21904 9548 21956
rect 9404 21836 9456 21888
rect 9680 21836 9732 21888
rect 10140 21904 10192 21956
rect 10600 21947 10652 21956
rect 10600 21913 10609 21947
rect 10609 21913 10643 21947
rect 10643 21913 10652 21947
rect 10600 21904 10652 21913
rect 10416 21836 10468 21888
rect 10508 21836 10560 21888
rect 11428 21972 11480 22024
rect 11888 21972 11940 22024
rect 12348 22040 12400 22092
rect 13176 22108 13228 22160
rect 13452 22108 13504 22160
rect 12440 21972 12492 22024
rect 11520 21947 11572 21956
rect 11520 21913 11529 21947
rect 11529 21913 11563 21947
rect 11563 21913 11572 21947
rect 11520 21904 11572 21913
rect 11796 21904 11848 21956
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 13360 22015 13412 22024
rect 13360 21981 13370 22015
rect 13370 21981 13404 22015
rect 13404 21981 13412 22015
rect 13360 21972 13412 21981
rect 13544 22015 13596 22024
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 13912 22176 13964 22228
rect 14280 22176 14332 22228
rect 14648 22176 14700 22228
rect 16488 22176 16540 22228
rect 16580 22176 16632 22228
rect 16948 22176 17000 22228
rect 13728 22108 13780 22160
rect 15292 22108 15344 22160
rect 17316 22151 17368 22160
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 14648 21972 14700 22024
rect 14924 22015 14976 22024
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 15016 21972 15068 22024
rect 16304 22040 16356 22092
rect 17316 22117 17325 22151
rect 17325 22117 17359 22151
rect 17359 22117 17368 22151
rect 17316 22108 17368 22117
rect 18236 22176 18288 22228
rect 17684 22083 17736 22092
rect 17684 22049 17693 22083
rect 17693 22049 17727 22083
rect 17727 22049 17736 22083
rect 17684 22040 17736 22049
rect 12256 21836 12308 21888
rect 12624 21879 12676 21888
rect 12624 21845 12633 21879
rect 12633 21845 12667 21879
rect 12667 21845 12676 21879
rect 12624 21836 12676 21845
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 14004 21836 14056 21888
rect 14556 21836 14608 21888
rect 15292 21904 15344 21956
rect 16580 21972 16632 22024
rect 15752 21836 15804 21888
rect 15936 21836 15988 21888
rect 16396 21836 16448 21888
rect 16948 21904 17000 21956
rect 17408 21972 17460 22024
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 18420 21972 18472 22024
rect 19524 22176 19576 22228
rect 19984 22176 20036 22228
rect 19340 22040 19392 22092
rect 19432 22040 19484 22092
rect 19800 22040 19852 22092
rect 17500 21904 17552 21956
rect 17684 21904 17736 21956
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 19064 21972 19116 22024
rect 20444 22108 20496 22160
rect 20812 22108 20864 22160
rect 20996 22176 21048 22228
rect 21640 22176 21692 22228
rect 24216 22219 24268 22228
rect 24216 22185 24225 22219
rect 24225 22185 24259 22219
rect 24259 22185 24268 22219
rect 24216 22176 24268 22185
rect 24400 22176 24452 22228
rect 21364 22108 21416 22160
rect 20720 22040 20772 22092
rect 19156 21904 19208 21956
rect 20260 22015 20312 22024
rect 20260 21981 20269 22015
rect 20269 21981 20303 22015
rect 20303 21981 20312 22015
rect 20260 21972 20312 21981
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 21180 22040 21232 22092
rect 21732 22040 21784 22092
rect 22192 22040 22244 22092
rect 21272 21972 21324 22024
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 18052 21836 18104 21888
rect 19616 21836 19668 21888
rect 21088 21904 21140 21956
rect 22560 21972 22612 22024
rect 22744 21972 22796 22024
rect 23112 21972 23164 22024
rect 23756 22040 23808 22092
rect 24584 22108 24636 22160
rect 24676 22108 24728 22160
rect 23664 21972 23716 22024
rect 23388 21947 23440 21956
rect 23388 21913 23397 21947
rect 23397 21913 23431 21947
rect 23431 21913 23440 21947
rect 23388 21904 23440 21913
rect 23848 21972 23900 22024
rect 24768 22015 24820 22024
rect 20444 21879 20496 21888
rect 20444 21845 20453 21879
rect 20453 21845 20487 21879
rect 20487 21845 20496 21879
rect 20444 21836 20496 21845
rect 21180 21836 21232 21888
rect 21640 21836 21692 21888
rect 22560 21879 22612 21888
rect 22560 21845 22569 21879
rect 22569 21845 22603 21879
rect 22603 21845 22612 21879
rect 22560 21836 22612 21845
rect 23296 21836 23348 21888
rect 23664 21836 23716 21888
rect 24032 21904 24084 21956
rect 24768 21981 24774 22015
rect 24774 21981 24808 22015
rect 24808 21981 24820 22015
rect 24768 21972 24820 21981
rect 24676 21947 24728 21956
rect 24676 21913 24685 21947
rect 24685 21913 24719 21947
rect 24719 21913 24728 21947
rect 24676 21904 24728 21913
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25596 22108 25648 22160
rect 26700 22219 26752 22228
rect 26700 22185 26709 22219
rect 26709 22185 26743 22219
rect 26743 22185 26752 22219
rect 26700 22176 26752 22185
rect 27896 22176 27948 22228
rect 28080 22176 28132 22228
rect 26056 22108 26108 22160
rect 25596 22015 25648 22024
rect 25596 21981 25610 22015
rect 25610 21981 25644 22015
rect 25644 21981 25648 22015
rect 25596 21972 25648 21981
rect 25780 21972 25832 22024
rect 26148 22040 26200 22092
rect 26332 22015 26384 22024
rect 26332 21981 26346 22015
rect 26346 21981 26380 22015
rect 26380 21981 26384 22015
rect 26332 21972 26384 21981
rect 26608 22015 26660 22024
rect 26608 21981 26617 22015
rect 26617 21981 26651 22015
rect 26651 21981 26660 22015
rect 26608 21972 26660 21981
rect 26792 21972 26844 22024
rect 27436 22040 27488 22092
rect 28080 22040 28132 22092
rect 26976 21972 27028 22024
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 28356 21972 28408 22024
rect 26148 21947 26200 21956
rect 26148 21913 26157 21947
rect 26157 21913 26191 21947
rect 26191 21913 26200 21947
rect 26148 21904 26200 21913
rect 27344 21904 27396 21956
rect 28816 22015 28868 22024
rect 28816 21981 28825 22015
rect 28825 21981 28859 22015
rect 28859 21981 28868 22015
rect 28816 21972 28868 21981
rect 28540 21904 28592 21956
rect 24492 21836 24544 21888
rect 24768 21836 24820 21888
rect 25872 21836 25924 21888
rect 26884 21836 26936 21888
rect 27068 21879 27120 21888
rect 27068 21845 27077 21879
rect 27077 21845 27111 21879
rect 27111 21845 27120 21879
rect 27068 21836 27120 21845
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 27988 21836 28040 21888
rect 28264 21836 28316 21888
rect 28448 21836 28500 21888
rect 29092 21879 29144 21888
rect 29092 21845 29101 21879
rect 29101 21845 29135 21879
rect 29135 21845 29144 21879
rect 29092 21836 29144 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1952 21607 2004 21616
rect 1952 21573 1961 21607
rect 1961 21573 1995 21607
rect 1995 21573 2004 21607
rect 1952 21564 2004 21573
rect 2412 21564 2464 21616
rect 2872 21632 2924 21684
rect 3700 21632 3752 21684
rect 4436 21632 4488 21684
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 1860 21292 1912 21344
rect 3516 21428 3568 21480
rect 3884 21428 3936 21480
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 4252 21539 4304 21548
rect 4252 21505 4287 21539
rect 4287 21505 4304 21539
rect 4252 21496 4304 21505
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 5448 21632 5500 21684
rect 5632 21675 5684 21684
rect 5632 21641 5641 21675
rect 5641 21641 5675 21675
rect 5675 21641 5684 21675
rect 5632 21632 5684 21641
rect 5724 21632 5776 21684
rect 6000 21632 6052 21684
rect 5264 21607 5316 21616
rect 5264 21573 5273 21607
rect 5273 21573 5307 21607
rect 5307 21573 5316 21607
rect 5264 21564 5316 21573
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 6276 21564 6328 21616
rect 7288 21564 7340 21616
rect 8024 21632 8076 21684
rect 5816 21496 5868 21548
rect 4344 21360 4396 21412
rect 4528 21360 4580 21412
rect 6092 21471 6144 21480
rect 6092 21437 6101 21471
rect 6101 21437 6135 21471
rect 6135 21437 6144 21471
rect 6092 21428 6144 21437
rect 6828 21496 6880 21548
rect 7380 21496 7432 21548
rect 8300 21607 8352 21616
rect 7012 21428 7064 21480
rect 6368 21360 6420 21412
rect 7196 21360 7248 21412
rect 7656 21360 7708 21412
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 8300 21573 8309 21607
rect 8309 21573 8343 21607
rect 8343 21573 8352 21607
rect 8300 21564 8352 21573
rect 8852 21632 8904 21684
rect 9220 21632 9272 21684
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 10600 21632 10652 21684
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11428 21632 11480 21684
rect 11520 21632 11572 21684
rect 10048 21564 10100 21616
rect 10784 21564 10836 21616
rect 11888 21632 11940 21684
rect 13084 21632 13136 21684
rect 13268 21675 13320 21684
rect 13268 21641 13277 21675
rect 13277 21641 13311 21675
rect 13311 21641 13320 21675
rect 13268 21632 13320 21641
rect 13360 21632 13412 21684
rect 12808 21564 12860 21616
rect 8208 21496 8260 21548
rect 8668 21496 8720 21548
rect 8852 21428 8904 21480
rect 8392 21360 8444 21412
rect 8944 21360 8996 21412
rect 9312 21496 9364 21548
rect 10876 21496 10928 21548
rect 11060 21539 11112 21548
rect 11060 21505 11069 21539
rect 11069 21505 11103 21539
rect 11103 21505 11112 21539
rect 11060 21496 11112 21505
rect 9496 21428 9548 21480
rect 11888 21496 11940 21548
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 12624 21539 12676 21548
rect 12624 21505 12633 21539
rect 12633 21505 12667 21539
rect 12667 21505 12676 21539
rect 13636 21607 13688 21616
rect 13636 21573 13645 21607
rect 13645 21573 13679 21607
rect 13679 21573 13688 21607
rect 13636 21564 13688 21573
rect 14832 21632 14884 21684
rect 15476 21632 15528 21684
rect 15568 21632 15620 21684
rect 15936 21632 15988 21684
rect 16304 21675 16356 21684
rect 16304 21641 16313 21675
rect 16313 21641 16347 21675
rect 16347 21641 16356 21675
rect 16304 21632 16356 21641
rect 16396 21632 16448 21684
rect 17500 21632 17552 21684
rect 12624 21496 12676 21505
rect 13544 21539 13596 21548
rect 13544 21505 13551 21539
rect 13551 21505 13596 21539
rect 12900 21428 12952 21480
rect 10600 21360 10652 21412
rect 11980 21360 12032 21412
rect 12072 21360 12124 21412
rect 2504 21292 2556 21344
rect 3424 21292 3476 21344
rect 4436 21292 4488 21344
rect 7288 21292 7340 21344
rect 8852 21292 8904 21344
rect 9036 21292 9088 21344
rect 9772 21292 9824 21344
rect 10416 21292 10468 21344
rect 12440 21292 12492 21344
rect 12716 21360 12768 21412
rect 12808 21292 12860 21344
rect 13544 21496 13596 21505
rect 14004 21496 14056 21548
rect 14280 21496 14332 21548
rect 14924 21564 14976 21616
rect 15016 21496 15068 21548
rect 15108 21539 15160 21548
rect 15108 21505 15117 21539
rect 15117 21505 15151 21539
rect 15151 21505 15160 21539
rect 15108 21496 15160 21505
rect 19340 21632 19392 21684
rect 21088 21632 21140 21684
rect 21364 21632 21416 21684
rect 18052 21564 18104 21616
rect 14740 21428 14792 21480
rect 16396 21496 16448 21548
rect 16580 21496 16632 21548
rect 16764 21496 16816 21548
rect 17132 21496 17184 21548
rect 15292 21360 15344 21412
rect 16304 21428 16356 21480
rect 15752 21360 15804 21412
rect 17040 21360 17092 21412
rect 17132 21360 17184 21412
rect 13636 21292 13688 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 14004 21292 14056 21301
rect 14372 21292 14424 21344
rect 14740 21292 14792 21344
rect 14924 21335 14976 21344
rect 14924 21301 14933 21335
rect 14933 21301 14967 21335
rect 14967 21301 14976 21335
rect 14924 21292 14976 21301
rect 15200 21292 15252 21344
rect 16672 21335 16724 21344
rect 16672 21301 16681 21335
rect 16681 21301 16715 21335
rect 16715 21301 16724 21335
rect 16672 21292 16724 21301
rect 17316 21292 17368 21344
rect 17684 21496 17736 21548
rect 18052 21428 18104 21480
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 18788 21496 18840 21548
rect 18972 21539 19024 21548
rect 18972 21505 18981 21539
rect 18981 21505 19015 21539
rect 19015 21505 19024 21539
rect 18972 21496 19024 21505
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 17500 21335 17552 21344
rect 17500 21301 17509 21335
rect 17509 21301 17543 21335
rect 17543 21301 17552 21335
rect 17500 21292 17552 21301
rect 17960 21335 18012 21344
rect 17960 21301 17969 21335
rect 17969 21301 18003 21335
rect 18003 21301 18012 21335
rect 17960 21292 18012 21301
rect 18052 21292 18104 21344
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 19156 21360 19208 21412
rect 19616 21496 19668 21548
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 20444 21564 20496 21616
rect 20812 21564 20864 21616
rect 21824 21564 21876 21616
rect 22468 21607 22520 21616
rect 22468 21573 22477 21607
rect 22477 21573 22511 21607
rect 22511 21573 22520 21607
rect 22468 21564 22520 21573
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 20536 21496 20588 21548
rect 21088 21496 21140 21548
rect 21364 21539 21416 21548
rect 21364 21505 21373 21539
rect 21373 21505 21407 21539
rect 21407 21505 21416 21539
rect 21364 21496 21416 21505
rect 21548 21496 21600 21548
rect 21916 21539 21968 21548
rect 21916 21505 21925 21539
rect 21925 21505 21959 21539
rect 21959 21505 21968 21539
rect 21916 21496 21968 21505
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 22652 21564 22704 21616
rect 22836 21539 22888 21548
rect 22836 21505 22865 21539
rect 22865 21505 22888 21539
rect 22836 21496 22888 21505
rect 19340 21292 19392 21344
rect 19800 21292 19852 21344
rect 19892 21292 19944 21344
rect 22468 21428 22520 21480
rect 22744 21428 22796 21480
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 23572 21564 23624 21616
rect 23848 21564 23900 21616
rect 24768 21632 24820 21684
rect 25596 21632 25648 21684
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 22928 21292 22980 21344
rect 23020 21292 23072 21344
rect 23572 21428 23624 21480
rect 23756 21471 23808 21480
rect 23756 21437 23765 21471
rect 23765 21437 23799 21471
rect 23799 21437 23808 21471
rect 23756 21428 23808 21437
rect 23848 21428 23900 21480
rect 23848 21292 23900 21344
rect 24584 21607 24636 21616
rect 24584 21573 24593 21607
rect 24593 21573 24627 21607
rect 24627 21573 24636 21607
rect 24584 21564 24636 21573
rect 26056 21564 26108 21616
rect 26976 21632 27028 21684
rect 27068 21632 27120 21684
rect 27344 21632 27396 21684
rect 26332 21564 26384 21616
rect 24124 21496 24176 21548
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 25872 21496 25924 21548
rect 26608 21496 26660 21548
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27436 21496 27488 21548
rect 24492 21428 24544 21480
rect 24860 21428 24912 21480
rect 24952 21428 25004 21480
rect 26792 21428 26844 21480
rect 28264 21539 28316 21548
rect 28264 21505 28278 21539
rect 28278 21505 28312 21539
rect 28312 21505 28316 21539
rect 28264 21496 28316 21505
rect 28632 21496 28684 21548
rect 28724 21496 28776 21548
rect 26700 21360 26752 21412
rect 28540 21428 28592 21480
rect 25872 21292 25924 21344
rect 26424 21335 26476 21344
rect 26424 21301 26433 21335
rect 26433 21301 26467 21335
rect 26467 21301 26476 21335
rect 26424 21292 26476 21301
rect 27160 21335 27212 21344
rect 27160 21301 27169 21335
rect 27169 21301 27203 21335
rect 27203 21301 27212 21335
rect 27160 21292 27212 21301
rect 27712 21292 27764 21344
rect 28356 21360 28408 21412
rect 28172 21335 28224 21344
rect 28172 21301 28181 21335
rect 28181 21301 28215 21335
rect 28215 21301 28224 21335
rect 28172 21292 28224 21301
rect 29184 21292 29236 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2136 21088 2188 21140
rect 2780 21088 2832 21140
rect 2964 21088 3016 21140
rect 1216 20952 1268 21004
rect 1952 20884 2004 20936
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 3332 20927 3384 20936
rect 3332 20893 3341 20927
rect 3341 20893 3375 20927
rect 3375 20893 3384 20927
rect 3332 20884 3384 20893
rect 3608 20952 3660 21004
rect 1676 20816 1728 20868
rect 4712 20952 4764 21004
rect 5540 21020 5592 21072
rect 5632 21020 5684 21072
rect 6000 21088 6052 21140
rect 6736 21088 6788 21140
rect 6276 21020 6328 21072
rect 6920 21088 6972 21140
rect 7288 21088 7340 21140
rect 7472 21088 7524 21140
rect 7840 21088 7892 21140
rect 7932 21088 7984 21140
rect 5356 20952 5408 21004
rect 3792 20884 3844 20936
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 4528 20927 4580 20936
rect 4528 20893 4537 20927
rect 4537 20893 4571 20927
rect 4571 20893 4580 20927
rect 4528 20884 4580 20893
rect 3424 20748 3476 20800
rect 4712 20816 4764 20868
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 7380 21063 7432 21072
rect 7380 21029 7389 21063
rect 7389 21029 7423 21063
rect 7423 21029 7432 21063
rect 7380 21020 7432 21029
rect 10232 21088 10284 21140
rect 10324 21088 10376 21140
rect 10416 21088 10468 21140
rect 10784 21088 10836 21140
rect 7748 20952 7800 21004
rect 8024 20952 8076 21004
rect 6920 20884 6972 20936
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 7196 20927 7248 20936
rect 7196 20893 7210 20927
rect 7210 20893 7244 20927
rect 7244 20893 7248 20927
rect 7196 20884 7248 20893
rect 5540 20859 5592 20868
rect 5540 20825 5549 20859
rect 5549 20825 5583 20859
rect 5583 20825 5592 20859
rect 5540 20816 5592 20825
rect 8024 20816 8076 20868
rect 8300 20884 8352 20936
rect 8392 20859 8444 20868
rect 8392 20825 8401 20859
rect 8401 20825 8435 20859
rect 8435 20825 8444 20859
rect 8392 20816 8444 20825
rect 8852 20884 8904 20936
rect 9036 20927 9088 20936
rect 9036 20893 9046 20927
rect 9046 20893 9080 20927
rect 9080 20893 9088 20927
rect 9036 20884 9088 20893
rect 9588 20952 9640 21004
rect 9404 20927 9456 20936
rect 9404 20893 9418 20927
rect 9418 20893 9452 20927
rect 9452 20893 9456 20927
rect 10324 20952 10376 21004
rect 11152 21020 11204 21072
rect 9404 20884 9456 20893
rect 9864 20884 9916 20936
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 9496 20816 9548 20868
rect 10232 20816 10284 20868
rect 5080 20748 5132 20800
rect 5908 20748 5960 20800
rect 6828 20748 6880 20800
rect 6920 20748 6972 20800
rect 7288 20748 7340 20800
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 9772 20748 9824 20800
rect 11060 20884 11112 20936
rect 12256 21088 12308 21140
rect 12624 21088 12676 21140
rect 17500 21088 17552 21140
rect 18696 21088 18748 21140
rect 14924 21020 14976 21072
rect 17224 21020 17276 21072
rect 10784 20859 10836 20868
rect 10784 20825 10793 20859
rect 10793 20825 10827 20859
rect 10827 20825 10836 20859
rect 10784 20816 10836 20825
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 13084 20995 13136 21004
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 13176 20927 13228 20936
rect 13176 20893 13185 20927
rect 13185 20893 13219 20927
rect 13219 20893 13228 20927
rect 13176 20884 13228 20893
rect 13820 20927 13872 20936
rect 13820 20893 13829 20927
rect 13829 20893 13863 20927
rect 13863 20893 13872 20927
rect 13820 20884 13872 20893
rect 10968 20748 11020 20800
rect 11060 20791 11112 20800
rect 11060 20757 11069 20791
rect 11069 20757 11103 20791
rect 11103 20757 11112 20791
rect 11060 20748 11112 20757
rect 11520 20748 11572 20800
rect 11612 20748 11664 20800
rect 12072 20748 12124 20800
rect 12164 20748 12216 20800
rect 14004 20816 14056 20868
rect 14188 20816 14240 20868
rect 14464 20816 14516 20868
rect 14832 20927 14884 20936
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 17592 20952 17644 21004
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 16120 20816 16172 20868
rect 16304 20816 16356 20868
rect 16488 20816 16540 20868
rect 12716 20791 12768 20800
rect 12716 20757 12725 20791
rect 12725 20757 12759 20791
rect 12759 20757 12768 20791
rect 12716 20748 12768 20757
rect 12900 20748 12952 20800
rect 13820 20748 13872 20800
rect 14832 20748 14884 20800
rect 14924 20748 14976 20800
rect 15016 20791 15068 20800
rect 15016 20757 15025 20791
rect 15025 20757 15059 20791
rect 15059 20757 15068 20791
rect 15016 20748 15068 20757
rect 15936 20748 15988 20800
rect 16580 20748 16632 20800
rect 17224 20884 17276 20936
rect 18052 20952 18104 21004
rect 18512 21020 18564 21072
rect 19616 21131 19668 21140
rect 19616 21097 19625 21131
rect 19625 21097 19659 21131
rect 19659 21097 19668 21131
rect 19616 21088 19668 21097
rect 17592 20748 17644 20800
rect 18052 20816 18104 20868
rect 18144 20816 18196 20868
rect 18788 20927 18840 20936
rect 18788 20893 18797 20927
rect 18797 20893 18831 20927
rect 18831 20893 18840 20927
rect 18788 20884 18840 20893
rect 18972 20884 19024 20936
rect 19432 20952 19484 21004
rect 21732 21088 21784 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 22008 21088 22060 21140
rect 22192 21088 22244 21140
rect 20996 21020 21048 21072
rect 19340 20884 19392 20936
rect 18604 20816 18656 20868
rect 19892 20884 19944 20936
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 20628 20884 20680 20893
rect 21180 20952 21232 21004
rect 18420 20748 18472 20800
rect 18972 20748 19024 20800
rect 19524 20748 19576 20800
rect 20260 20816 20312 20868
rect 21548 20884 21600 20936
rect 22836 21020 22888 21072
rect 22744 20952 22796 21004
rect 22192 20884 22244 20936
rect 22284 20927 22336 20936
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 19800 20748 19852 20800
rect 20076 20748 20128 20800
rect 20628 20748 20680 20800
rect 21180 20816 21232 20868
rect 22468 20884 22520 20936
rect 23296 21088 23348 21140
rect 23480 21088 23532 21140
rect 24400 21088 24452 21140
rect 23112 20884 23164 20936
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23940 20884 23992 20936
rect 23848 20859 23900 20868
rect 20812 20748 20864 20800
rect 22284 20748 22336 20800
rect 23848 20825 23857 20859
rect 23857 20825 23891 20859
rect 23891 20825 23900 20859
rect 23848 20816 23900 20825
rect 24032 20859 24084 20868
rect 24032 20825 24057 20859
rect 24057 20825 24084 20859
rect 24032 20816 24084 20825
rect 23664 20748 23716 20800
rect 23940 20748 23992 20800
rect 24216 20791 24268 20800
rect 24216 20757 24225 20791
rect 24225 20757 24259 20791
rect 24259 20757 24268 20791
rect 24216 20748 24268 20757
rect 24492 20748 24544 20800
rect 24860 20884 24912 20936
rect 25320 21131 25372 21140
rect 25320 21097 25329 21131
rect 25329 21097 25363 21131
rect 25363 21097 25372 21131
rect 25320 21088 25372 21097
rect 25872 21020 25924 21072
rect 27252 21131 27304 21140
rect 27252 21097 27261 21131
rect 27261 21097 27295 21131
rect 27295 21097 27304 21131
rect 27252 21088 27304 21097
rect 27344 21088 27396 21140
rect 26884 21020 26936 21072
rect 25228 20884 25280 20936
rect 25504 20884 25556 20936
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 26056 20927 26108 20936
rect 26056 20893 26065 20927
rect 26065 20893 26099 20927
rect 26099 20893 26108 20927
rect 26056 20884 26108 20893
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 26148 20884 26200 20893
rect 26608 20995 26660 21004
rect 26608 20961 26617 20995
rect 26617 20961 26651 20995
rect 26651 20961 26660 20995
rect 26608 20952 26660 20961
rect 27252 20952 27304 21004
rect 28080 21131 28132 21140
rect 28080 21097 28089 21131
rect 28089 21097 28123 21131
rect 28123 21097 28132 21131
rect 28080 21088 28132 21097
rect 28172 21088 28224 21140
rect 30196 21088 30248 21140
rect 27712 21020 27764 21072
rect 26424 20927 26476 20936
rect 26424 20893 26433 20927
rect 26433 20893 26467 20927
rect 26467 20893 26476 20927
rect 26424 20884 26476 20893
rect 26884 20884 26936 20936
rect 24676 20816 24728 20825
rect 28632 20884 28684 20936
rect 28816 20884 28868 20936
rect 28908 20884 28960 20936
rect 29460 20884 29512 20936
rect 25504 20748 25556 20800
rect 25596 20791 25648 20800
rect 25596 20757 25605 20791
rect 25605 20757 25639 20791
rect 25639 20757 25648 20791
rect 25596 20748 25648 20757
rect 26240 20748 26292 20800
rect 27344 20748 27396 20800
rect 27436 20748 27488 20800
rect 28632 20748 28684 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5264 20544 5316 20596
rect 5356 20544 5408 20596
rect 3424 20476 3476 20528
rect 3700 20519 3752 20528
rect 3700 20485 3709 20519
rect 3709 20485 3743 20519
rect 3743 20485 3752 20519
rect 3700 20476 3752 20485
rect 3884 20476 3936 20528
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 1860 20408 1912 20460
rect 2964 20408 3016 20460
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 4160 20408 4212 20417
rect 4896 20408 4948 20460
rect 5632 20476 5684 20528
rect 5816 20544 5868 20596
rect 6460 20544 6512 20596
rect 5540 20408 5592 20460
rect 2780 20340 2832 20392
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 6276 20408 6328 20460
rect 6184 20340 6236 20392
rect 5816 20272 5868 20324
rect 6092 20272 6144 20324
rect 6736 20451 6788 20460
rect 6736 20417 6746 20451
rect 6746 20417 6780 20451
rect 6780 20417 6788 20451
rect 7288 20544 7340 20596
rect 7932 20544 7984 20596
rect 9036 20544 9088 20596
rect 6736 20408 6788 20417
rect 7104 20408 7156 20460
rect 8392 20519 8444 20528
rect 8392 20485 8401 20519
rect 8401 20485 8435 20519
rect 8435 20485 8444 20519
rect 8392 20476 8444 20485
rect 9496 20476 9548 20528
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 7564 20383 7616 20392
rect 7564 20349 7573 20383
rect 7573 20349 7607 20383
rect 7607 20349 7616 20383
rect 7564 20340 7616 20349
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 8484 20451 8536 20460
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 8392 20340 8444 20392
rect 8852 20408 8904 20460
rect 9312 20408 9364 20460
rect 9404 20408 9456 20460
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 10416 20544 10468 20596
rect 11888 20544 11940 20596
rect 13084 20544 13136 20596
rect 14280 20544 14332 20596
rect 15108 20544 15160 20596
rect 15844 20544 15896 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 16396 20544 16448 20596
rect 17684 20544 17736 20596
rect 10508 20519 10560 20528
rect 10508 20485 10517 20519
rect 10517 20485 10551 20519
rect 10551 20485 10560 20519
rect 10508 20476 10560 20485
rect 9220 20340 9272 20392
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 10876 20451 10928 20460
rect 10876 20417 10891 20451
rect 10891 20417 10925 20451
rect 10925 20417 10928 20451
rect 10876 20408 10928 20417
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 3608 20204 3660 20256
rect 5172 20204 5224 20256
rect 6184 20247 6236 20256
rect 6184 20213 6193 20247
rect 6193 20213 6227 20247
rect 6227 20213 6236 20247
rect 6184 20204 6236 20213
rect 7288 20204 7340 20256
rect 7380 20204 7432 20256
rect 8760 20272 8812 20324
rect 8024 20247 8076 20256
rect 8024 20213 8033 20247
rect 8033 20213 8067 20247
rect 8067 20213 8076 20247
rect 8024 20204 8076 20213
rect 8300 20204 8352 20256
rect 10600 20340 10652 20392
rect 10968 20340 11020 20392
rect 11520 20408 11572 20460
rect 12072 20408 12124 20460
rect 15016 20476 15068 20528
rect 11152 20340 11204 20392
rect 12164 20340 12216 20392
rect 9772 20272 9824 20324
rect 12900 20408 12952 20460
rect 14280 20408 14332 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 14188 20340 14240 20392
rect 16028 20408 16080 20460
rect 16212 20408 16264 20460
rect 17592 20476 17644 20528
rect 17960 20544 18012 20596
rect 18144 20544 18196 20596
rect 18420 20587 18472 20596
rect 18420 20553 18429 20587
rect 18429 20553 18463 20587
rect 18463 20553 18472 20587
rect 18420 20544 18472 20553
rect 18880 20544 18932 20596
rect 21272 20544 21324 20596
rect 21640 20544 21692 20596
rect 17132 20408 17184 20460
rect 17224 20408 17276 20460
rect 17316 20408 17368 20460
rect 16856 20340 16908 20392
rect 17776 20408 17828 20460
rect 18144 20408 18196 20460
rect 18328 20408 18380 20460
rect 18420 20408 18472 20460
rect 19248 20408 19300 20460
rect 19984 20476 20036 20528
rect 21088 20476 21140 20528
rect 22008 20476 22060 20528
rect 22468 20476 22520 20528
rect 19432 20340 19484 20392
rect 19616 20408 19668 20460
rect 19708 20408 19760 20460
rect 20536 20408 20588 20460
rect 24492 20587 24544 20596
rect 24492 20553 24501 20587
rect 24501 20553 24535 20587
rect 24535 20553 24544 20587
rect 24492 20544 24544 20553
rect 22928 20451 22980 20460
rect 22928 20417 22937 20451
rect 22937 20417 22971 20451
rect 22971 20417 22980 20451
rect 22928 20408 22980 20417
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23480 20408 23532 20460
rect 24124 20408 24176 20460
rect 24216 20408 24268 20460
rect 19800 20340 19852 20392
rect 19892 20340 19944 20392
rect 20812 20340 20864 20392
rect 21088 20340 21140 20392
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 24400 20340 24452 20392
rect 17040 20272 17092 20324
rect 20352 20272 20404 20324
rect 24584 20476 24636 20528
rect 24768 20451 24820 20460
rect 24768 20417 24777 20451
rect 24777 20417 24811 20451
rect 24811 20417 24820 20451
rect 24768 20408 24820 20417
rect 25412 20544 25464 20596
rect 25596 20544 25648 20596
rect 25964 20476 26016 20528
rect 26976 20544 27028 20596
rect 28264 20544 28316 20596
rect 10232 20204 10284 20256
rect 10876 20204 10928 20256
rect 11152 20204 11204 20256
rect 12072 20204 12124 20256
rect 12532 20204 12584 20256
rect 13268 20204 13320 20256
rect 13820 20204 13872 20256
rect 16396 20204 16448 20256
rect 17500 20204 17552 20256
rect 17592 20204 17644 20256
rect 24768 20272 24820 20324
rect 21088 20204 21140 20256
rect 22192 20204 22244 20256
rect 23296 20204 23348 20256
rect 23664 20204 23716 20256
rect 23756 20247 23808 20256
rect 23756 20213 23765 20247
rect 23765 20213 23799 20247
rect 23799 20213 23808 20247
rect 23756 20204 23808 20213
rect 24308 20204 24360 20256
rect 24952 20204 25004 20256
rect 25780 20451 25832 20460
rect 25780 20417 25789 20451
rect 25789 20417 25823 20451
rect 25823 20417 25832 20451
rect 25780 20408 25832 20417
rect 26240 20408 26292 20460
rect 25504 20340 25556 20392
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 26240 20315 26292 20324
rect 26240 20281 26249 20315
rect 26249 20281 26283 20315
rect 26283 20281 26292 20315
rect 26240 20272 26292 20281
rect 27896 20476 27948 20528
rect 27068 20408 27120 20460
rect 27344 20408 27396 20460
rect 28264 20451 28316 20460
rect 28264 20417 28273 20451
rect 28273 20417 28307 20451
rect 28307 20417 28316 20451
rect 28264 20408 28316 20417
rect 28448 20451 28500 20460
rect 28448 20417 28457 20451
rect 28457 20417 28491 20451
rect 28491 20417 28500 20451
rect 28448 20408 28500 20417
rect 28540 20408 28592 20460
rect 29092 20408 29144 20460
rect 27804 20383 27856 20392
rect 27804 20349 27813 20383
rect 27813 20349 27847 20383
rect 27847 20349 27856 20383
rect 27804 20340 27856 20349
rect 28172 20340 28224 20392
rect 25320 20204 25372 20256
rect 25412 20247 25464 20256
rect 25412 20213 25421 20247
rect 25421 20213 25455 20247
rect 25455 20213 25464 20247
rect 25412 20204 25464 20213
rect 25688 20204 25740 20256
rect 26792 20204 26844 20256
rect 27344 20272 27396 20324
rect 27436 20272 27488 20324
rect 27804 20204 27856 20256
rect 28080 20204 28132 20256
rect 28172 20247 28224 20256
rect 28172 20213 28181 20247
rect 28181 20213 28215 20247
rect 28215 20213 28224 20247
rect 28172 20204 28224 20213
rect 28448 20204 28500 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2964 20000 3016 20052
rect 3792 20000 3844 20052
rect 4896 20000 4948 20052
rect 4988 20000 5040 20052
rect 5632 20000 5684 20052
rect 6000 20000 6052 20052
rect 6460 20000 6512 20052
rect 8024 20000 8076 20052
rect 9036 20000 9088 20052
rect 12900 20000 12952 20052
rect 15200 20000 15252 20052
rect 17684 20000 17736 20052
rect 18604 20000 18656 20052
rect 19156 20000 19208 20052
rect 21088 20000 21140 20052
rect 21640 20000 21692 20052
rect 22744 20000 22796 20052
rect 24124 20000 24176 20052
rect 24768 20000 24820 20052
rect 25412 20043 25464 20052
rect 25412 20009 25421 20043
rect 25421 20009 25455 20043
rect 25455 20009 25464 20043
rect 25412 20000 25464 20009
rect 25780 20043 25832 20052
rect 25780 20009 25789 20043
rect 25789 20009 25823 20043
rect 25823 20009 25832 20043
rect 25780 20000 25832 20009
rect 26424 20000 26476 20052
rect 27528 20043 27580 20052
rect 7288 19932 7340 19984
rect 1216 19864 1268 19916
rect 3056 19907 3108 19916
rect 3056 19873 3065 19907
rect 3065 19873 3099 19907
rect 3099 19873 3108 19907
rect 3056 19864 3108 19873
rect 3240 19864 3292 19916
rect 10968 19932 11020 19984
rect 11980 19932 12032 19984
rect 3700 19796 3752 19848
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 4988 19796 5040 19805
rect 5080 19839 5132 19848
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 3976 19728 4028 19780
rect 5264 19796 5316 19848
rect 9128 19864 9180 19916
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 11704 19864 11756 19916
rect 11888 19864 11940 19916
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 12992 19932 13044 19984
rect 16212 19975 16264 19984
rect 16212 19941 16221 19975
rect 16221 19941 16255 19975
rect 16255 19941 16264 19975
rect 16212 19932 16264 19941
rect 6368 19796 6420 19848
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6828 19728 6880 19780
rect 5264 19660 5316 19712
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 7472 19796 7524 19848
rect 8208 19796 8260 19848
rect 9680 19796 9732 19848
rect 10416 19796 10468 19848
rect 10784 19796 10836 19848
rect 11520 19796 11572 19848
rect 8484 19728 8536 19780
rect 8852 19728 8904 19780
rect 10692 19728 10744 19780
rect 8392 19660 8444 19712
rect 10140 19660 10192 19712
rect 10324 19660 10376 19712
rect 12348 19728 12400 19780
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 13544 19864 13596 19916
rect 13084 19796 13136 19848
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 12992 19728 13044 19780
rect 14464 19728 14516 19780
rect 12808 19660 12860 19712
rect 13084 19660 13136 19712
rect 14188 19660 14240 19712
rect 14648 19796 14700 19848
rect 14832 19796 14884 19848
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15292 19796 15344 19848
rect 15384 19796 15436 19848
rect 16764 19932 16816 19984
rect 16856 19932 16908 19984
rect 18972 19932 19024 19984
rect 15660 19728 15712 19780
rect 18604 19864 18656 19916
rect 15016 19660 15068 19712
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 17592 19796 17644 19848
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 17316 19728 17368 19780
rect 18328 19796 18380 19848
rect 18788 19796 18840 19848
rect 19340 19864 19392 19916
rect 20168 19975 20220 19984
rect 20168 19941 20177 19975
rect 20177 19941 20211 19975
rect 20211 19941 20220 19975
rect 20168 19932 20220 19941
rect 21732 19932 21784 19984
rect 22192 19932 22244 19984
rect 22468 19932 22520 19984
rect 24032 19932 24084 19984
rect 24216 19932 24268 19984
rect 24860 19932 24912 19984
rect 25136 19932 25188 19984
rect 20628 19864 20680 19916
rect 20812 19864 20864 19916
rect 22100 19864 22152 19916
rect 23296 19864 23348 19916
rect 23848 19864 23900 19916
rect 19156 19796 19208 19848
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 20076 19796 20128 19848
rect 20352 19728 20404 19780
rect 20536 19796 20588 19848
rect 18236 19660 18288 19712
rect 18420 19660 18472 19712
rect 18880 19660 18932 19712
rect 19524 19660 19576 19712
rect 19984 19660 20036 19712
rect 20904 19796 20956 19848
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 21916 19796 21968 19848
rect 24400 19796 24452 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 24676 19796 24728 19848
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 21272 19660 21324 19712
rect 22100 19660 22152 19712
rect 22744 19728 22796 19780
rect 24308 19728 24360 19780
rect 24768 19771 24820 19780
rect 24768 19737 24777 19771
rect 24777 19737 24811 19771
rect 24811 19737 24820 19771
rect 24768 19728 24820 19737
rect 25136 19796 25188 19848
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 26148 19864 26200 19916
rect 23480 19703 23532 19712
rect 23480 19669 23489 19703
rect 23489 19669 23523 19703
rect 23523 19669 23532 19703
rect 23480 19660 23532 19669
rect 23756 19660 23808 19712
rect 25044 19660 25096 19712
rect 25780 19796 25832 19848
rect 26332 19864 26384 19916
rect 26516 19839 26568 19848
rect 26516 19805 26525 19839
rect 26525 19805 26559 19839
rect 26559 19805 26568 19839
rect 26516 19796 26568 19805
rect 26608 19839 26660 19848
rect 26608 19805 26617 19839
rect 26617 19805 26651 19839
rect 26651 19805 26660 19839
rect 26608 19796 26660 19805
rect 26332 19728 26384 19780
rect 26884 19771 26936 19780
rect 26884 19737 26893 19771
rect 26893 19737 26927 19771
rect 26927 19737 26936 19771
rect 26884 19728 26936 19737
rect 26976 19728 27028 19780
rect 27528 20009 27537 20043
rect 27537 20009 27571 20043
rect 27571 20009 27580 20043
rect 27528 20000 27580 20009
rect 27896 20043 27948 20052
rect 27896 20009 27905 20043
rect 27905 20009 27939 20043
rect 27939 20009 27948 20043
rect 27896 20000 27948 20009
rect 28356 20000 28408 20052
rect 27252 19932 27304 19984
rect 27436 19864 27488 19916
rect 29184 19864 29236 19916
rect 27436 19771 27488 19780
rect 27436 19737 27445 19771
rect 27445 19737 27479 19771
rect 27479 19737 27488 19771
rect 27436 19728 27488 19737
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 28264 19796 28316 19848
rect 29092 19796 29144 19848
rect 28724 19728 28776 19780
rect 27712 19660 27764 19712
rect 28356 19703 28408 19712
rect 28356 19669 28365 19703
rect 28365 19669 28399 19703
rect 28399 19669 28408 19703
rect 28356 19660 28408 19669
rect 28816 19703 28868 19712
rect 28816 19669 28825 19703
rect 28825 19669 28859 19703
rect 28859 19669 28868 19703
rect 28816 19660 28868 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3056 19456 3108 19508
rect 3332 19456 3384 19508
rect 3792 19456 3844 19508
rect 5724 19456 5776 19508
rect 6276 19456 6328 19508
rect 6736 19456 6788 19508
rect 3516 19320 3568 19372
rect 4068 19320 4120 19372
rect 5356 19388 5408 19440
rect 4528 19320 4580 19372
rect 4804 19320 4856 19372
rect 4988 19363 5040 19372
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 1492 19252 1544 19304
rect 1768 19252 1820 19304
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 2872 19116 2924 19168
rect 4252 19184 4304 19236
rect 5172 19252 5224 19304
rect 5264 19252 5316 19304
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 5816 19320 5868 19372
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6000 19320 6052 19372
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6644 19388 6696 19440
rect 7380 19456 7432 19508
rect 8300 19456 8352 19508
rect 8484 19499 8536 19508
rect 8484 19465 8493 19499
rect 8493 19465 8527 19499
rect 8527 19465 8536 19499
rect 8484 19456 8536 19465
rect 8760 19456 8812 19508
rect 6920 19320 6972 19372
rect 7196 19320 7248 19372
rect 9404 19499 9456 19508
rect 9404 19465 9413 19499
rect 9413 19465 9447 19499
rect 9447 19465 9456 19499
rect 9404 19456 9456 19465
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 10508 19456 10560 19508
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 10140 19388 10192 19440
rect 12348 19456 12400 19508
rect 12532 19456 12584 19508
rect 12624 19499 12676 19508
rect 12624 19465 12633 19499
rect 12633 19465 12667 19499
rect 12667 19465 12676 19499
rect 12624 19456 12676 19465
rect 12716 19456 12768 19508
rect 6552 19184 6604 19236
rect 7288 19184 7340 19236
rect 7656 19184 7708 19236
rect 8760 19184 8812 19236
rect 9128 19320 9180 19372
rect 9312 19363 9364 19372
rect 9312 19329 9321 19363
rect 9321 19329 9355 19363
rect 9355 19329 9364 19363
rect 9312 19320 9364 19329
rect 10324 19320 10376 19372
rect 12072 19388 12124 19440
rect 12164 19388 12216 19440
rect 11704 19320 11756 19372
rect 11980 19363 12032 19372
rect 11980 19329 11989 19363
rect 11989 19329 12023 19363
rect 12023 19329 12032 19363
rect 11980 19320 12032 19329
rect 12256 19320 12308 19372
rect 12992 19431 13044 19440
rect 12992 19397 13001 19431
rect 13001 19397 13035 19431
rect 13035 19397 13044 19431
rect 12992 19388 13044 19397
rect 10048 19295 10100 19304
rect 10048 19261 10057 19295
rect 10057 19261 10091 19295
rect 10091 19261 10100 19295
rect 10048 19252 10100 19261
rect 10140 19252 10192 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 9036 19184 9088 19236
rect 9128 19184 9180 19236
rect 10508 19184 10560 19236
rect 3332 19159 3384 19168
rect 3332 19125 3341 19159
rect 3341 19125 3375 19159
rect 3375 19125 3384 19159
rect 3332 19116 3384 19125
rect 5540 19116 5592 19168
rect 5816 19116 5868 19168
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 8852 19116 8904 19168
rect 12624 19252 12676 19304
rect 13268 19363 13320 19372
rect 13268 19329 13277 19363
rect 13277 19329 13311 19363
rect 13311 19329 13320 19363
rect 13268 19320 13320 19329
rect 12716 19184 12768 19236
rect 15108 19456 15160 19508
rect 14096 19431 14148 19440
rect 14096 19397 14105 19431
rect 14105 19397 14139 19431
rect 14139 19397 14148 19431
rect 14096 19388 14148 19397
rect 13452 19184 13504 19236
rect 13728 19184 13780 19236
rect 14464 19320 14516 19372
rect 15384 19388 15436 19440
rect 15752 19456 15804 19508
rect 16672 19456 16724 19508
rect 16764 19499 16816 19508
rect 16764 19465 16773 19499
rect 16773 19465 16807 19499
rect 16807 19465 16816 19499
rect 16764 19456 16816 19465
rect 15936 19320 15988 19372
rect 17132 19320 17184 19372
rect 17224 19320 17276 19372
rect 18788 19456 18840 19508
rect 17776 19388 17828 19440
rect 19248 19456 19300 19508
rect 19340 19456 19392 19508
rect 18328 19363 18380 19372
rect 14924 19252 14976 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 17040 19252 17092 19304
rect 18328 19329 18337 19363
rect 18337 19329 18371 19363
rect 18371 19329 18380 19363
rect 18328 19320 18380 19329
rect 18788 19320 18840 19372
rect 19156 19388 19208 19440
rect 19340 19320 19392 19372
rect 19892 19388 19944 19440
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 17500 19184 17552 19236
rect 18236 19252 18288 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18880 19252 18932 19304
rect 20628 19388 20680 19440
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20812 19431 20864 19440
rect 20812 19397 20821 19431
rect 20821 19397 20855 19431
rect 20855 19397 20864 19431
rect 20812 19388 20864 19397
rect 21548 19388 21600 19440
rect 21916 19456 21968 19508
rect 22652 19456 22704 19508
rect 23112 19499 23164 19508
rect 23112 19465 23121 19499
rect 23121 19465 23155 19499
rect 23155 19465 23164 19499
rect 23112 19456 23164 19465
rect 23572 19388 23624 19440
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 21732 19320 21784 19372
rect 18144 19227 18196 19236
rect 18144 19193 18153 19227
rect 18153 19193 18187 19227
rect 18187 19193 18196 19227
rect 18144 19184 18196 19193
rect 12808 19116 12860 19168
rect 13820 19116 13872 19168
rect 14648 19116 14700 19168
rect 15384 19116 15436 19168
rect 19156 19184 19208 19236
rect 19708 19184 19760 19236
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 18972 19116 19024 19168
rect 20076 19116 20128 19168
rect 20812 19184 20864 19236
rect 21456 19227 21508 19236
rect 21456 19193 21465 19227
rect 21465 19193 21499 19227
rect 21499 19193 21508 19227
rect 21456 19184 21508 19193
rect 22100 19252 22152 19304
rect 22284 19252 22336 19304
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 24124 19431 24176 19440
rect 24124 19397 24133 19431
rect 24133 19397 24167 19431
rect 24167 19397 24176 19431
rect 24124 19388 24176 19397
rect 24400 19456 24452 19508
rect 25320 19456 25372 19508
rect 25596 19456 25648 19508
rect 25688 19456 25740 19508
rect 23940 19363 23992 19372
rect 23940 19329 23950 19363
rect 23950 19329 23984 19363
rect 23984 19329 23992 19363
rect 23940 19320 23992 19329
rect 21916 19116 21968 19168
rect 22652 19184 22704 19236
rect 23480 19184 23532 19236
rect 27344 19431 27396 19440
rect 27344 19397 27353 19431
rect 27353 19397 27387 19431
rect 27387 19397 27396 19431
rect 27344 19388 27396 19397
rect 27620 19388 27672 19440
rect 24676 19320 24728 19372
rect 24952 19320 25004 19372
rect 24952 19184 25004 19236
rect 25320 19320 25372 19372
rect 26608 19320 26660 19372
rect 25964 19295 26016 19304
rect 25964 19261 25973 19295
rect 25973 19261 26007 19295
rect 26007 19261 26016 19295
rect 25964 19252 26016 19261
rect 26148 19184 26200 19236
rect 24584 19116 24636 19168
rect 27252 19252 27304 19304
rect 28448 19456 28500 19508
rect 28632 19499 28684 19508
rect 28632 19465 28641 19499
rect 28641 19465 28675 19499
rect 28675 19465 28684 19499
rect 28632 19456 28684 19465
rect 27804 19295 27856 19304
rect 27804 19261 27813 19295
rect 27813 19261 27847 19295
rect 27847 19261 27856 19295
rect 27804 19252 27856 19261
rect 27252 19116 27304 19168
rect 27712 19159 27764 19168
rect 27712 19125 27721 19159
rect 27721 19125 27755 19159
rect 27755 19125 27764 19159
rect 27712 19116 27764 19125
rect 28172 19159 28224 19168
rect 28172 19125 28181 19159
rect 28181 19125 28215 19159
rect 28215 19125 28224 19159
rect 28172 19116 28224 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 4068 18912 4120 18964
rect 5172 18912 5224 18964
rect 5908 18912 5960 18964
rect 7840 18912 7892 18964
rect 8392 18955 8444 18964
rect 8392 18921 8401 18955
rect 8401 18921 8435 18955
rect 8435 18921 8444 18955
rect 8392 18912 8444 18921
rect 8760 18912 8812 18964
rect 1860 18776 1912 18828
rect 5264 18776 5316 18828
rect 6092 18844 6144 18896
rect 6184 18844 6236 18896
rect 2688 18708 2740 18760
rect 3332 18708 3384 18760
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 6368 18776 6420 18828
rect 8300 18844 8352 18896
rect 6184 18751 6236 18760
rect 6184 18717 6194 18751
rect 6194 18717 6228 18751
rect 6228 18717 6236 18751
rect 6184 18708 6236 18717
rect 1216 18640 1268 18692
rect 6552 18751 6604 18760
rect 6552 18717 6566 18751
rect 6566 18717 6600 18751
rect 6600 18717 6604 18751
rect 6552 18708 6604 18717
rect 4896 18640 4948 18692
rect 6000 18640 6052 18692
rect 6276 18640 6328 18692
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 8208 18708 8260 18760
rect 9404 18708 9456 18760
rect 7932 18683 7984 18692
rect 5080 18572 5132 18624
rect 6552 18572 6604 18624
rect 7932 18649 7941 18683
rect 7941 18649 7975 18683
rect 7975 18649 7984 18683
rect 7932 18640 7984 18649
rect 6736 18572 6788 18624
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 7380 18572 7432 18624
rect 7564 18572 7616 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 8208 18572 8260 18624
rect 8392 18572 8444 18624
rect 8852 18640 8904 18692
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 11704 18912 11756 18964
rect 12164 18912 12216 18964
rect 15016 18912 15068 18964
rect 15844 18912 15896 18964
rect 15936 18955 15988 18964
rect 15936 18921 15945 18955
rect 15945 18921 15979 18955
rect 15979 18921 15988 18955
rect 15936 18912 15988 18921
rect 16120 18912 16172 18964
rect 11520 18844 11572 18896
rect 13084 18844 13136 18896
rect 13176 18887 13228 18896
rect 13176 18853 13185 18887
rect 13185 18853 13219 18887
rect 13219 18853 13228 18887
rect 13176 18844 13228 18853
rect 10968 18776 11020 18828
rect 14280 18844 14332 18896
rect 14556 18844 14608 18896
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10876 18708 10928 18760
rect 11704 18708 11756 18760
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 12256 18708 12308 18760
rect 12716 18708 12768 18760
rect 13820 18708 13872 18760
rect 15844 18776 15896 18828
rect 17316 18844 17368 18896
rect 17868 18912 17920 18964
rect 19984 18912 20036 18964
rect 20260 18912 20312 18964
rect 22928 18912 22980 18964
rect 23388 18912 23440 18964
rect 10416 18683 10468 18692
rect 10416 18649 10425 18683
rect 10425 18649 10459 18683
rect 10459 18649 10468 18683
rect 10416 18640 10468 18649
rect 10508 18683 10560 18692
rect 10508 18649 10543 18683
rect 10543 18649 10560 18683
rect 10508 18640 10560 18649
rect 11152 18640 11204 18692
rect 13268 18640 13320 18692
rect 14280 18708 14332 18760
rect 9036 18572 9088 18624
rect 10968 18572 11020 18624
rect 11796 18572 11848 18624
rect 12164 18572 12216 18624
rect 12532 18572 12584 18624
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 14556 18640 14608 18692
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16120 18708 16172 18760
rect 16304 18708 16356 18760
rect 16488 18708 16540 18760
rect 13728 18572 13780 18624
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 14004 18572 14056 18624
rect 15844 18572 15896 18624
rect 16764 18708 16816 18760
rect 18604 18776 18656 18828
rect 18880 18776 18932 18828
rect 21364 18844 21416 18896
rect 21732 18844 21784 18896
rect 22008 18844 22060 18896
rect 22468 18844 22520 18896
rect 19248 18776 19300 18828
rect 17132 18572 17184 18624
rect 17960 18708 18012 18760
rect 18236 18708 18288 18760
rect 18328 18708 18380 18760
rect 18420 18683 18472 18692
rect 18420 18649 18429 18683
rect 18429 18649 18463 18683
rect 18463 18649 18472 18683
rect 18420 18640 18472 18649
rect 18788 18708 18840 18760
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 19524 18640 19576 18692
rect 20076 18683 20128 18692
rect 20076 18649 20085 18683
rect 20085 18649 20119 18683
rect 20119 18649 20128 18683
rect 20076 18640 20128 18649
rect 20168 18572 20220 18624
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 22192 18776 22244 18828
rect 20444 18572 20496 18624
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 21916 18708 21968 18760
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22744 18776 22796 18828
rect 23480 18844 23532 18896
rect 24216 18955 24268 18964
rect 24216 18921 24225 18955
rect 24225 18921 24259 18955
rect 24259 18921 24268 18955
rect 24216 18912 24268 18921
rect 24492 18912 24544 18964
rect 24584 18955 24636 18964
rect 24584 18921 24593 18955
rect 24593 18921 24627 18955
rect 24627 18921 24636 18955
rect 24584 18912 24636 18921
rect 25044 18912 25096 18964
rect 25688 18912 25740 18964
rect 24124 18776 24176 18828
rect 24676 18844 24728 18896
rect 26148 18844 26200 18896
rect 26884 18912 26936 18964
rect 29092 18955 29144 18964
rect 29092 18921 29101 18955
rect 29101 18921 29135 18955
rect 29135 18921 29144 18955
rect 29092 18912 29144 18921
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 23664 18708 23716 18760
rect 23756 18751 23808 18760
rect 23756 18717 23765 18751
rect 23765 18717 23799 18751
rect 23799 18717 23808 18751
rect 23756 18708 23808 18717
rect 24032 18708 24084 18760
rect 23848 18683 23900 18692
rect 23848 18649 23857 18683
rect 23857 18649 23891 18683
rect 23891 18649 23900 18683
rect 23848 18640 23900 18649
rect 22192 18572 22244 18624
rect 22468 18615 22520 18624
rect 22468 18581 22477 18615
rect 22477 18581 22511 18615
rect 22511 18581 22520 18615
rect 22468 18572 22520 18581
rect 23112 18572 23164 18624
rect 23940 18572 23992 18624
rect 24308 18708 24360 18760
rect 24400 18751 24452 18760
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 24952 18640 25004 18692
rect 25044 18572 25096 18624
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 26976 18844 27028 18896
rect 26148 18683 26200 18692
rect 26148 18649 26157 18683
rect 26157 18649 26191 18683
rect 26191 18649 26200 18683
rect 26148 18640 26200 18649
rect 25964 18572 26016 18624
rect 26056 18572 26108 18624
rect 27252 18708 27304 18760
rect 27620 18708 27672 18760
rect 27988 18751 28040 18760
rect 27988 18717 28022 18751
rect 28022 18717 28040 18751
rect 27988 18708 28040 18717
rect 26700 18572 26752 18624
rect 28908 18640 28960 18692
rect 27252 18615 27304 18624
rect 27252 18581 27261 18615
rect 27261 18581 27295 18615
rect 27295 18581 27304 18615
rect 27252 18572 27304 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 4896 18411 4948 18420
rect 4896 18377 4905 18411
rect 4905 18377 4939 18411
rect 4939 18377 4948 18411
rect 4896 18368 4948 18377
rect 5080 18368 5132 18420
rect 5632 18368 5684 18420
rect 6000 18368 6052 18420
rect 2596 18300 2648 18352
rect 4804 18300 4856 18352
rect 1768 18232 1820 18284
rect 3240 18232 3292 18284
rect 5908 18300 5960 18352
rect 6368 18300 6420 18352
rect 6920 18300 6972 18352
rect 7380 18368 7432 18420
rect 7932 18411 7984 18420
rect 7932 18377 7941 18411
rect 7941 18377 7975 18411
rect 7975 18377 7984 18411
rect 7932 18368 7984 18377
rect 8484 18368 8536 18420
rect 5816 18275 5868 18284
rect 3700 18164 3752 18216
rect 3884 18164 3936 18216
rect 4620 18164 4672 18216
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 5816 18232 5868 18241
rect 5448 18164 5500 18216
rect 6092 18232 6144 18284
rect 6460 18164 6512 18216
rect 5908 18096 5960 18148
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 6920 18164 6972 18216
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 8208 18300 8260 18352
rect 6736 18096 6788 18148
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 8392 18275 8444 18284
rect 8392 18241 8405 18275
rect 8405 18241 8439 18275
rect 8439 18241 8444 18275
rect 8392 18232 8444 18241
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 3884 18028 3936 18080
rect 4712 18028 4764 18080
rect 7196 18028 7248 18080
rect 7288 18028 7340 18080
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 9036 18368 9088 18420
rect 9956 18368 10008 18420
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 7748 18028 7800 18080
rect 8852 18139 8904 18148
rect 8852 18105 8861 18139
rect 8861 18105 8895 18139
rect 8895 18105 8904 18139
rect 8852 18096 8904 18105
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9588 18232 9640 18284
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 10600 18300 10652 18352
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 12808 18368 12860 18420
rect 12992 18368 13044 18420
rect 13544 18368 13596 18420
rect 13820 18368 13872 18420
rect 14556 18368 14608 18420
rect 14740 18368 14792 18420
rect 15936 18368 15988 18420
rect 16488 18411 16540 18420
rect 16488 18377 16497 18411
rect 16497 18377 16531 18411
rect 16531 18377 16540 18411
rect 16488 18368 16540 18377
rect 16672 18368 16724 18420
rect 11152 18300 11204 18352
rect 11980 18343 12032 18352
rect 10416 18232 10468 18284
rect 11980 18309 11989 18343
rect 11989 18309 12023 18343
rect 12023 18309 12032 18343
rect 11980 18300 12032 18309
rect 12624 18300 12676 18352
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 11704 18164 11756 18216
rect 9220 18096 9272 18148
rect 10416 18096 10468 18148
rect 10876 18096 10928 18148
rect 11520 18096 11572 18148
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 13176 18164 13228 18216
rect 13452 18232 13504 18284
rect 14004 18232 14056 18284
rect 9036 18028 9088 18080
rect 9128 18028 9180 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 11612 18071 11664 18080
rect 11612 18037 11621 18071
rect 11621 18037 11655 18071
rect 11655 18037 11664 18071
rect 11612 18028 11664 18037
rect 11980 18028 12032 18080
rect 12900 18028 12952 18080
rect 13452 18096 13504 18148
rect 13728 18096 13780 18148
rect 14280 18164 14332 18216
rect 14648 18232 14700 18284
rect 14648 18096 14700 18148
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 15016 18232 15068 18284
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 16580 18300 16632 18352
rect 17960 18368 18012 18420
rect 18328 18368 18380 18420
rect 18788 18368 18840 18420
rect 15844 18232 15896 18284
rect 15476 18164 15528 18216
rect 16028 18164 16080 18216
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17500 18232 17552 18284
rect 17684 18232 17736 18284
rect 18052 18232 18104 18284
rect 19432 18300 19484 18352
rect 19708 18300 19760 18352
rect 19892 18368 19944 18420
rect 20444 18368 20496 18420
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 21180 18368 21232 18420
rect 21364 18368 21416 18420
rect 17408 18164 17460 18216
rect 19156 18275 19208 18284
rect 19156 18241 19165 18275
rect 19165 18241 19199 18275
rect 19199 18241 19208 18275
rect 19156 18232 19208 18241
rect 19984 18232 20036 18284
rect 20628 18232 20680 18284
rect 20904 18232 20956 18284
rect 14924 18096 14976 18148
rect 15292 18096 15344 18148
rect 13084 18028 13136 18080
rect 13544 18028 13596 18080
rect 14004 18028 14056 18080
rect 14372 18028 14424 18080
rect 14556 18028 14608 18080
rect 17040 18096 17092 18148
rect 17592 18139 17644 18148
rect 17592 18105 17601 18139
rect 17601 18105 17635 18139
rect 17635 18105 17644 18139
rect 17592 18096 17644 18105
rect 18052 18096 18104 18148
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 18604 18096 18656 18148
rect 20168 18096 20220 18148
rect 20720 18096 20772 18148
rect 21548 18275 21600 18284
rect 21548 18241 21557 18275
rect 21557 18241 21591 18275
rect 21591 18241 21600 18275
rect 21548 18232 21600 18241
rect 24124 18368 24176 18420
rect 22652 18343 22704 18352
rect 22652 18309 22661 18343
rect 22661 18309 22695 18343
rect 22695 18309 22704 18343
rect 22652 18300 22704 18309
rect 23296 18300 23348 18352
rect 25228 18368 25280 18420
rect 25412 18368 25464 18420
rect 26056 18368 26108 18420
rect 26424 18368 26476 18420
rect 28080 18368 28132 18420
rect 21824 18232 21876 18284
rect 21916 18232 21968 18284
rect 21732 18096 21784 18148
rect 23940 18232 23992 18284
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 22468 18164 22520 18216
rect 22928 18164 22980 18216
rect 23020 18164 23072 18216
rect 24400 18275 24452 18284
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 24676 18232 24728 18284
rect 24584 18164 24636 18216
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 25412 18232 25464 18284
rect 28172 18300 28224 18352
rect 25596 18232 25648 18284
rect 25688 18164 25740 18216
rect 26884 18164 26936 18216
rect 27620 18232 27672 18284
rect 18512 18028 18564 18080
rect 18696 18028 18748 18080
rect 19800 18028 19852 18080
rect 22008 18028 22060 18080
rect 24032 18028 24084 18080
rect 24492 18096 24544 18148
rect 25044 18028 25096 18080
rect 26056 18071 26108 18080
rect 26056 18037 26065 18071
rect 26065 18037 26099 18071
rect 26099 18037 26108 18071
rect 26056 18028 26108 18037
rect 26700 18139 26752 18148
rect 26700 18105 26709 18139
rect 26709 18105 26743 18139
rect 26743 18105 26752 18139
rect 26700 18096 26752 18105
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3516 17824 3568 17876
rect 4620 17824 4672 17876
rect 5540 17824 5592 17876
rect 6828 17824 6880 17876
rect 1216 17688 1268 17740
rect 1676 17620 1728 17672
rect 2964 17731 3016 17740
rect 2964 17697 2973 17731
rect 2973 17697 3007 17731
rect 3007 17697 3016 17731
rect 2964 17688 3016 17697
rect 3608 17688 3660 17740
rect 4620 17688 4672 17740
rect 3424 17620 3476 17672
rect 3884 17620 3936 17672
rect 4436 17620 4488 17672
rect 5816 17756 5868 17808
rect 6460 17756 6512 17808
rect 6644 17756 6696 17808
rect 4804 17688 4856 17740
rect 5632 17688 5684 17740
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 7380 17731 7432 17740
rect 7380 17697 7389 17731
rect 7389 17697 7423 17731
rect 7423 17697 7432 17731
rect 7380 17688 7432 17697
rect 7932 17824 7984 17876
rect 8760 17824 8812 17876
rect 8116 17756 8168 17808
rect 9036 17756 9088 17808
rect 8300 17688 8352 17740
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 5908 17663 5960 17672
rect 5908 17629 5917 17663
rect 5917 17629 5951 17663
rect 5951 17629 5960 17663
rect 5908 17620 5960 17629
rect 5724 17595 5776 17604
rect 5724 17561 5733 17595
rect 5733 17561 5767 17595
rect 5767 17561 5776 17595
rect 5724 17552 5776 17561
rect 5632 17484 5684 17536
rect 6092 17620 6144 17672
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 7840 17663 7892 17672
rect 7840 17629 7849 17663
rect 7849 17629 7883 17663
rect 7883 17629 7892 17663
rect 7840 17620 7892 17629
rect 8852 17688 8904 17740
rect 6644 17552 6696 17604
rect 6092 17527 6144 17536
rect 6092 17493 6101 17527
rect 6101 17493 6135 17527
rect 6135 17493 6144 17527
rect 6092 17484 6144 17493
rect 6552 17484 6604 17536
rect 7748 17552 7800 17604
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 13452 17824 13504 17876
rect 14280 17824 14332 17876
rect 10232 17756 10284 17808
rect 10876 17688 10928 17740
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 10324 17620 10376 17672
rect 10416 17620 10468 17672
rect 13544 17756 13596 17808
rect 17040 17824 17092 17876
rect 17960 17824 18012 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 19064 17824 19116 17876
rect 21180 17867 21232 17876
rect 21180 17833 21189 17867
rect 21189 17833 21223 17867
rect 21223 17833 21232 17867
rect 21180 17824 21232 17833
rect 21548 17824 21600 17876
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 23204 17824 23256 17876
rect 11520 17688 11572 17740
rect 11612 17688 11664 17740
rect 12808 17688 12860 17740
rect 13360 17688 13412 17740
rect 7932 17484 7984 17536
rect 8392 17484 8444 17536
rect 8576 17484 8628 17536
rect 9404 17484 9456 17536
rect 9772 17484 9824 17536
rect 10508 17552 10560 17604
rect 11888 17620 11940 17672
rect 12900 17620 12952 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 15292 17756 15344 17808
rect 14648 17688 14700 17740
rect 15752 17688 15804 17740
rect 16948 17756 17000 17808
rect 17592 17799 17644 17808
rect 17592 17765 17601 17799
rect 17601 17765 17635 17799
rect 17635 17765 17644 17799
rect 17592 17756 17644 17765
rect 18696 17799 18748 17808
rect 18696 17765 18705 17799
rect 18705 17765 18739 17799
rect 18739 17765 18748 17799
rect 18696 17756 18748 17765
rect 18052 17731 18104 17740
rect 18052 17697 18061 17731
rect 18061 17697 18095 17731
rect 18095 17697 18104 17731
rect 18052 17688 18104 17697
rect 18420 17688 18472 17740
rect 10876 17552 10928 17604
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 13636 17595 13688 17604
rect 13636 17561 13645 17595
rect 13645 17561 13679 17595
rect 13679 17561 13688 17595
rect 13636 17552 13688 17561
rect 14280 17552 14332 17604
rect 14372 17595 14424 17604
rect 14372 17561 14381 17595
rect 14381 17561 14415 17595
rect 14415 17561 14424 17595
rect 14372 17552 14424 17561
rect 14832 17620 14884 17672
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 15476 17620 15528 17672
rect 15844 17620 15896 17672
rect 14924 17484 14976 17536
rect 15108 17484 15160 17536
rect 15292 17484 15344 17536
rect 16580 17620 16632 17672
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 16488 17595 16540 17604
rect 16488 17561 16497 17595
rect 16497 17561 16531 17595
rect 16531 17561 16540 17595
rect 16488 17552 16540 17561
rect 16212 17484 16264 17536
rect 16304 17484 16356 17536
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 17684 17620 17736 17672
rect 17592 17552 17644 17604
rect 17500 17484 17552 17536
rect 21916 17799 21968 17808
rect 21916 17765 21925 17799
rect 21925 17765 21959 17799
rect 21959 17765 21968 17799
rect 21916 17756 21968 17765
rect 22008 17756 22060 17808
rect 23296 17756 23348 17808
rect 24676 17824 24728 17876
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 19432 17552 19484 17604
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 19800 17620 19852 17672
rect 19984 17620 20036 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 20996 17620 21048 17672
rect 20720 17552 20772 17604
rect 21180 17663 21232 17672
rect 21180 17629 21189 17663
rect 21189 17629 21223 17663
rect 21223 17629 21232 17663
rect 21180 17620 21232 17629
rect 21364 17731 21416 17740
rect 21364 17697 21373 17731
rect 21373 17697 21407 17731
rect 21407 17697 21416 17731
rect 21364 17688 21416 17697
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 24768 17688 24820 17740
rect 21916 17620 21968 17672
rect 22376 17663 22428 17672
rect 22376 17629 22385 17663
rect 22385 17629 22419 17663
rect 22419 17629 22428 17663
rect 22376 17620 22428 17629
rect 23112 17620 23164 17672
rect 23480 17620 23532 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 25136 17824 25188 17876
rect 25412 17867 25464 17876
rect 25412 17833 25421 17867
rect 25421 17833 25455 17867
rect 25455 17833 25464 17867
rect 25412 17824 25464 17833
rect 25596 17824 25648 17876
rect 26148 17824 26200 17876
rect 26792 17867 26844 17876
rect 26792 17833 26801 17867
rect 26801 17833 26835 17867
rect 26835 17833 26844 17867
rect 26792 17824 26844 17833
rect 21364 17552 21416 17604
rect 22928 17552 22980 17604
rect 23388 17484 23440 17536
rect 23480 17484 23532 17536
rect 23664 17595 23716 17604
rect 23664 17561 23673 17595
rect 23673 17561 23707 17595
rect 23707 17561 23716 17595
rect 23664 17552 23716 17561
rect 24492 17552 24544 17604
rect 24676 17595 24728 17604
rect 24676 17561 24685 17595
rect 24685 17561 24719 17595
rect 24719 17561 24728 17595
rect 24676 17552 24728 17561
rect 24768 17595 24820 17604
rect 24768 17561 24777 17595
rect 24777 17561 24811 17595
rect 24811 17561 24820 17595
rect 24768 17552 24820 17561
rect 25320 17620 25372 17672
rect 26332 17688 26384 17740
rect 26976 17688 27028 17740
rect 25780 17620 25832 17672
rect 27252 17620 27304 17672
rect 27436 17620 27488 17672
rect 25504 17595 25556 17604
rect 25504 17561 25513 17595
rect 25513 17561 25547 17595
rect 25547 17561 25556 17595
rect 25504 17552 25556 17561
rect 25596 17552 25648 17604
rect 25872 17552 25924 17604
rect 25964 17595 26016 17604
rect 25964 17561 25973 17595
rect 25973 17561 26007 17595
rect 26007 17561 26016 17595
rect 25964 17552 26016 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 3240 17280 3292 17332
rect 4804 17280 4856 17332
rect 3332 17144 3384 17196
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 3792 17144 3844 17196
rect 4896 17144 4948 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 2872 17076 2924 17128
rect 6092 17280 6144 17332
rect 6368 17323 6420 17332
rect 6368 17289 6377 17323
rect 6377 17289 6411 17323
rect 6411 17289 6420 17323
rect 6368 17280 6420 17289
rect 5448 17255 5500 17264
rect 5448 17221 5457 17255
rect 5457 17221 5491 17255
rect 5491 17221 5500 17255
rect 5448 17212 5500 17221
rect 5540 17255 5592 17264
rect 5540 17221 5549 17255
rect 5549 17221 5583 17255
rect 5583 17221 5592 17255
rect 5540 17212 5592 17221
rect 5632 17255 5684 17264
rect 5632 17221 5667 17255
rect 5667 17221 5684 17255
rect 5632 17212 5684 17221
rect 6000 17212 6052 17264
rect 5632 17076 5684 17128
rect 5908 17076 5960 17128
rect 6092 17187 6144 17196
rect 6092 17153 6101 17187
rect 6101 17153 6135 17187
rect 6135 17153 6144 17187
rect 6092 17144 6144 17153
rect 6460 17144 6512 17196
rect 6828 17280 6880 17332
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 7840 17323 7892 17332
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 7104 17212 7156 17264
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 3240 16940 3292 16992
rect 4068 16940 4120 16992
rect 4436 16940 4488 16992
rect 5448 17008 5500 17060
rect 5724 17008 5776 17060
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 7564 17076 7616 17128
rect 7932 17212 7984 17264
rect 8484 17280 8536 17332
rect 8116 17255 8168 17264
rect 8116 17221 8125 17255
rect 8125 17221 8159 17255
rect 8159 17221 8168 17255
rect 8116 17212 8168 17221
rect 10508 17280 10560 17332
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 11336 17280 11388 17332
rect 10232 17212 10284 17264
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 9680 17144 9732 17196
rect 9772 17144 9824 17196
rect 10784 17187 10836 17196
rect 8484 17119 8536 17128
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 8300 17008 8352 17060
rect 11704 17280 11756 17332
rect 12072 17280 12124 17332
rect 12348 17280 12400 17332
rect 12716 17280 12768 17332
rect 12900 17323 12952 17332
rect 12900 17289 12909 17323
rect 12909 17289 12943 17323
rect 12943 17289 12952 17323
rect 12900 17280 12952 17289
rect 13084 17323 13136 17332
rect 13084 17289 13093 17323
rect 13093 17289 13127 17323
rect 13127 17289 13136 17323
rect 13084 17280 13136 17289
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 14556 17280 14608 17332
rect 14924 17280 14976 17332
rect 17500 17280 17552 17332
rect 18880 17280 18932 17332
rect 13268 17212 13320 17264
rect 12532 17144 12584 17196
rect 13176 17144 13228 17196
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11520 17076 11572 17085
rect 14004 17144 14056 17196
rect 14372 17144 14424 17196
rect 15292 17144 15344 17196
rect 15936 17212 15988 17264
rect 16304 17212 16356 17264
rect 7012 16940 7064 16992
rect 14004 17008 14056 17060
rect 15016 17008 15068 17060
rect 16304 17008 16356 17060
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 17684 17144 17736 17196
rect 18328 17144 18380 17196
rect 18512 17144 18564 17196
rect 18604 17076 18656 17128
rect 19156 17144 19208 17196
rect 20628 17323 20680 17332
rect 20628 17289 20637 17323
rect 20637 17289 20671 17323
rect 20671 17289 20680 17323
rect 20628 17280 20680 17289
rect 20904 17280 20956 17332
rect 21088 17212 21140 17264
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 19892 17144 19944 17196
rect 20076 17187 20128 17196
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 19248 17008 19300 17060
rect 21364 17255 21416 17264
rect 21364 17221 21373 17255
rect 21373 17221 21407 17255
rect 21407 17221 21416 17255
rect 21364 17212 21416 17221
rect 22468 17323 22520 17332
rect 22468 17289 22477 17323
rect 22477 17289 22511 17323
rect 22511 17289 22520 17323
rect 22468 17280 22520 17289
rect 22836 17323 22888 17332
rect 22836 17289 22845 17323
rect 22845 17289 22879 17323
rect 22879 17289 22888 17323
rect 22836 17280 22888 17289
rect 22928 17280 22980 17332
rect 23296 17280 23348 17332
rect 24768 17280 24820 17332
rect 43260 17323 43312 17332
rect 43260 17289 43269 17323
rect 43269 17289 43303 17323
rect 43303 17289 43312 17323
rect 43260 17280 43312 17289
rect 22652 17212 22704 17264
rect 21732 17144 21784 17196
rect 21456 17119 21508 17128
rect 21456 17085 21490 17119
rect 21490 17085 21508 17119
rect 21456 17076 21508 17085
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23480 17212 23532 17264
rect 24308 17212 24360 17264
rect 23572 17187 23624 17196
rect 23572 17153 23581 17187
rect 23581 17153 23615 17187
rect 23615 17153 23624 17187
rect 23572 17144 23624 17153
rect 43168 17187 43220 17196
rect 43168 17153 43177 17187
rect 43177 17153 43211 17187
rect 43211 17153 43220 17187
rect 43168 17144 43220 17153
rect 22008 17051 22060 17060
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 11796 16940 11848 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 14648 16940 14700 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 17684 16940 17736 16992
rect 19156 16940 19208 16992
rect 19984 16940 20036 16992
rect 20260 16940 20312 16992
rect 21088 16940 21140 16992
rect 22008 17017 22017 17051
rect 22017 17017 22051 17051
rect 22051 17017 22060 17051
rect 22008 17008 22060 17017
rect 21916 16940 21968 16992
rect 23112 17008 23164 17060
rect 24676 17076 24728 17128
rect 24492 17008 24544 17060
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3332 16736 3384 16788
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 5172 16736 5224 16788
rect 5632 16736 5684 16788
rect 3608 16600 3660 16652
rect 3792 16643 3844 16652
rect 3792 16609 3801 16643
rect 3801 16609 3835 16643
rect 3835 16609 3844 16643
rect 3792 16600 3844 16609
rect 1216 16464 1268 16516
rect 3056 16532 3108 16584
rect 7196 16668 7248 16720
rect 7012 16600 7064 16652
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 6552 16532 6604 16584
rect 8668 16736 8720 16788
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 11520 16736 11572 16788
rect 12256 16736 12308 16788
rect 13820 16736 13872 16788
rect 14280 16736 14332 16788
rect 15016 16736 15068 16788
rect 15660 16736 15712 16788
rect 16764 16736 16816 16788
rect 17040 16736 17092 16788
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 17592 16736 17644 16788
rect 18604 16736 18656 16788
rect 18880 16779 18932 16788
rect 18880 16745 18889 16779
rect 18889 16745 18923 16779
rect 18923 16745 18932 16779
rect 18880 16736 18932 16745
rect 10324 16668 10376 16720
rect 10784 16668 10836 16720
rect 7472 16532 7524 16584
rect 8392 16532 8444 16584
rect 8484 16532 8536 16584
rect 8300 16464 8352 16516
rect 9404 16532 9456 16584
rect 10692 16532 10744 16584
rect 11428 16532 11480 16584
rect 11980 16600 12032 16652
rect 11612 16575 11664 16584
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 12072 16532 12124 16584
rect 12808 16600 12860 16652
rect 13360 16668 13412 16720
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 13912 16600 13964 16652
rect 14004 16600 14056 16652
rect 15384 16668 15436 16720
rect 15936 16668 15988 16720
rect 17316 16668 17368 16720
rect 16304 16600 16356 16652
rect 11060 16396 11112 16448
rect 11980 16396 12032 16448
rect 12900 16439 12952 16448
rect 12900 16405 12909 16439
rect 12909 16405 12943 16439
rect 12943 16405 12952 16439
rect 12900 16396 12952 16405
rect 13268 16507 13320 16516
rect 13268 16473 13277 16507
rect 13277 16473 13311 16507
rect 13311 16473 13320 16507
rect 13268 16464 13320 16473
rect 13360 16464 13412 16516
rect 14004 16464 14056 16516
rect 13636 16396 13688 16448
rect 14464 16532 14516 16584
rect 14648 16575 14700 16584
rect 14648 16541 14682 16575
rect 14682 16541 14700 16575
rect 14648 16532 14700 16541
rect 15384 16532 15436 16584
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 19892 16736 19944 16788
rect 25504 16736 25556 16788
rect 19800 16668 19852 16720
rect 18328 16600 18380 16652
rect 19064 16600 19116 16652
rect 20444 16668 20496 16720
rect 24400 16668 24452 16720
rect 19156 16532 19208 16584
rect 20260 16532 20312 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 20812 16600 20864 16652
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 21088 16532 21140 16584
rect 21456 16532 21508 16584
rect 22376 16600 22428 16652
rect 22100 16575 22152 16584
rect 22100 16541 22109 16575
rect 22109 16541 22143 16575
rect 22143 16541 22152 16575
rect 22100 16532 22152 16541
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 22560 16532 22612 16584
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 16488 16396 16540 16448
rect 19248 16396 19300 16448
rect 19340 16396 19392 16448
rect 21364 16464 21416 16516
rect 22652 16464 22704 16516
rect 20720 16396 20772 16448
rect 21916 16396 21968 16448
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2872 16192 2924 16244
rect 4068 16192 4120 16244
rect 4988 16192 5040 16244
rect 6000 16192 6052 16244
rect 7564 16192 7616 16244
rect 8484 16192 8536 16244
rect 9680 16192 9732 16244
rect 9864 16192 9916 16244
rect 10048 16192 10100 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11612 16192 11664 16244
rect 12900 16192 12952 16244
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 16120 16235 16172 16244
rect 16120 16201 16129 16235
rect 16129 16201 16163 16235
rect 16163 16201 16172 16235
rect 16120 16192 16172 16201
rect 16764 16192 16816 16244
rect 19432 16192 19484 16244
rect 20352 16192 20404 16244
rect 22468 16192 22520 16244
rect 23020 16192 23072 16244
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 1860 16056 1912 16108
rect 2780 15852 2832 15904
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3700 15988 3752 16040
rect 3884 15988 3936 16040
rect 4896 16056 4948 16108
rect 4712 15988 4764 16040
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 6092 16056 6144 16108
rect 6460 16099 6512 16108
rect 6460 16065 6469 16099
rect 6469 16065 6503 16099
rect 6503 16065 6512 16099
rect 6460 16056 6512 16065
rect 7380 16056 7432 16108
rect 6000 15988 6052 16040
rect 7472 15988 7524 16040
rect 8208 16056 8260 16108
rect 8760 16031 8812 16040
rect 8760 15997 8769 16031
rect 8769 15997 8803 16031
rect 8803 15997 8812 16031
rect 8760 15988 8812 15997
rect 11704 16124 11756 16176
rect 13820 16167 13872 16176
rect 13820 16133 13829 16167
rect 13829 16133 13863 16167
rect 13863 16133 13872 16167
rect 13820 16124 13872 16133
rect 14280 16124 14332 16176
rect 15476 16124 15528 16176
rect 21364 16124 21416 16176
rect 10968 16056 11020 16108
rect 12256 16056 12308 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 19064 16056 19116 16108
rect 19156 16056 19208 16108
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 17132 15988 17184 16040
rect 4068 15852 4120 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 7748 15852 7800 15904
rect 8484 15852 8536 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 11336 15852 11388 15904
rect 20260 16031 20312 16040
rect 20260 15997 20269 16031
rect 20269 15997 20303 16031
rect 20303 15997 20312 16031
rect 20260 15988 20312 15997
rect 21640 15963 21692 15972
rect 21640 15929 21649 15963
rect 21649 15929 21683 15963
rect 21683 15929 21692 15963
rect 21640 15920 21692 15929
rect 13176 15852 13228 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 17408 15852 17460 15904
rect 17960 15895 18012 15904
rect 17960 15861 17969 15895
rect 17969 15861 18003 15895
rect 18003 15861 18012 15895
rect 17960 15852 18012 15861
rect 19248 15895 19300 15904
rect 19248 15861 19257 15895
rect 19257 15861 19291 15895
rect 19291 15861 19300 15895
rect 19248 15852 19300 15861
rect 26884 16124 26936 16176
rect 28356 16124 28408 16176
rect 28816 15852 28868 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3424 15648 3476 15700
rect 3884 15648 3936 15700
rect 1216 15512 1268 15564
rect 3148 15512 3200 15564
rect 5632 15648 5684 15700
rect 7288 15648 7340 15700
rect 8024 15648 8076 15700
rect 8760 15648 8812 15700
rect 5264 15580 5316 15632
rect 6184 15512 6236 15564
rect 8116 15512 8168 15564
rect 9220 15512 9272 15564
rect 9772 15512 9824 15564
rect 9956 15512 10008 15564
rect 3792 15376 3844 15428
rect 4068 15444 4120 15496
rect 5264 15444 5316 15496
rect 5356 15444 5408 15496
rect 4804 15376 4856 15428
rect 5540 15308 5592 15360
rect 5908 15444 5960 15496
rect 8944 15444 8996 15496
rect 11336 15648 11388 15700
rect 12808 15648 12860 15700
rect 13728 15648 13780 15700
rect 17132 15648 17184 15700
rect 20260 15648 20312 15700
rect 22468 15648 22520 15700
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 13912 15512 13964 15564
rect 6828 15308 6880 15360
rect 7380 15308 7432 15360
rect 9404 15351 9456 15360
rect 9404 15317 9413 15351
rect 9413 15317 9447 15351
rect 9447 15317 9456 15351
rect 9404 15308 9456 15317
rect 12256 15444 12308 15496
rect 15016 15580 15068 15632
rect 15568 15580 15620 15632
rect 16028 15623 16080 15632
rect 16028 15589 16037 15623
rect 16037 15589 16071 15623
rect 16071 15589 16080 15623
rect 16028 15580 16080 15589
rect 16304 15623 16356 15632
rect 16304 15589 16313 15623
rect 16313 15589 16347 15623
rect 16347 15589 16356 15623
rect 16304 15580 16356 15589
rect 14740 15512 14792 15564
rect 18512 15623 18564 15632
rect 18512 15589 18521 15623
rect 18521 15589 18555 15623
rect 18555 15589 18564 15623
rect 18512 15580 18564 15589
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 11520 15376 11572 15428
rect 10876 15308 10928 15360
rect 11060 15308 11112 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13452 15308 13504 15360
rect 17408 15487 17460 15496
rect 17408 15453 17442 15487
rect 17442 15453 17460 15487
rect 17408 15444 17460 15453
rect 26056 15444 26108 15496
rect 17960 15376 18012 15428
rect 22744 15376 22796 15428
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 2780 15104 2832 15156
rect 3056 15104 3108 15156
rect 3976 15147 4028 15156
rect 3976 15113 3985 15147
rect 3985 15113 4019 15147
rect 4019 15113 4028 15147
rect 3976 15104 4028 15113
rect 6184 15104 6236 15156
rect 2044 15036 2096 15088
rect 3240 14968 3292 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4620 14968 4672 15020
rect 5816 15036 5868 15088
rect 7472 15104 7524 15156
rect 7564 15104 7616 15156
rect 8024 15104 8076 15156
rect 6736 15079 6788 15088
rect 6736 15045 6745 15079
rect 6745 15045 6779 15079
rect 6779 15045 6788 15079
rect 6736 15036 6788 15045
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10784 15104 10836 15156
rect 3516 14900 3568 14952
rect 5816 14900 5868 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7380 14968 7432 15020
rect 8208 14968 8260 15020
rect 8484 14968 8536 15020
rect 12532 15104 12584 15156
rect 12992 15104 13044 15156
rect 14740 15104 14792 15156
rect 15016 15147 15068 15156
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11796 15011 11848 15020
rect 11520 14968 11572 14977
rect 11796 14977 11830 15011
rect 11830 14977 11848 15011
rect 11796 14968 11848 14977
rect 13452 15011 13504 15020
rect 13452 14977 13486 15011
rect 13486 14977 13504 15011
rect 13452 14968 13504 14977
rect 14464 14968 14516 15020
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 3240 14764 3292 14816
rect 3700 14764 3752 14816
rect 4712 14764 4764 14816
rect 7012 14764 7064 14816
rect 7380 14764 7432 14816
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 11796 14764 11848 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 4620 14560 4672 14612
rect 5172 14492 5224 14544
rect 6920 14560 6972 14612
rect 8116 14603 8168 14612
rect 8116 14569 8125 14603
rect 8125 14569 8159 14603
rect 8159 14569 8168 14603
rect 8116 14560 8168 14569
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 10048 14560 10100 14612
rect 10876 14560 10928 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 9772 14492 9824 14544
rect 13176 14492 13228 14544
rect 1216 14424 1268 14476
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 6644 14424 6696 14476
rect 4804 14356 4856 14408
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 7012 14399 7064 14408
rect 5264 14356 5316 14365
rect 5356 14288 5408 14340
rect 6184 14288 6236 14340
rect 7012 14365 7046 14399
rect 7046 14365 7064 14399
rect 7012 14356 7064 14365
rect 7564 14356 7616 14408
rect 6092 14220 6144 14272
rect 7656 14220 7708 14272
rect 8116 14220 8168 14272
rect 13360 14220 13412 14272
rect 14556 14220 14608 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14016 1728 14068
rect 2504 14016 2556 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 3240 13948 3292 14000
rect 4620 13948 4672 14000
rect 6092 13948 6144 14000
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 7104 14016 7156 14068
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 8208 14016 8260 14068
rect 10876 14016 10928 14068
rect 6920 13948 6972 14000
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 4620 13744 4672 13796
rect 6736 13744 6788 13796
rect 7840 13744 7892 13796
rect 6920 13676 6972 13728
rect 7380 13676 7432 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3792 13472 3844 13524
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 6276 13472 6328 13524
rect 8484 13472 8536 13524
rect 7380 13404 7432 13456
rect 1216 13336 1268 13388
rect 7840 13379 7892 13388
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 4712 13268 4764 13320
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 5172 12928 5224 12980
rect 6920 12928 6972 12980
rect 5816 12860 5868 12912
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1216 12248 1268 12300
rect 6828 12180 6880 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4620 11704 4672 11756
rect 11980 11704 12032 11756
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 7748 11092 7800 11144
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1216 10072 1268 10124
rect 9404 10004 9456 10056
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 11612 9596 11664 9648
rect 13360 9596 13412 9648
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1216 8984 1268 9036
rect 11152 8916 11204 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1216 7896 1268 7948
rect 4620 7828 4672 7880
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1216 6808 1268 6860
rect 11612 6740 11664 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 18512 5516 18564 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 1216 4632 1268 4684
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 1216 3544 1268 3596
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 24676 2635 24728 2644
rect 24676 2601 24685 2635
rect 24685 2601 24719 2635
rect 24719 2601 24728 2635
rect 24676 2592 24728 2601
rect 22468 2456 22520 2508
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 1490 44200 1546 45000
rect 2686 44200 2742 45000
rect 3882 44200 3938 45000
rect 5078 44200 5134 45000
rect 6274 44200 6330 45000
rect 7470 44200 7526 45000
rect 8666 44200 8722 45000
rect 9862 44200 9918 45000
rect 11058 44200 11114 45000
rect 12254 44200 12310 45000
rect 13450 44200 13506 45000
rect 14646 44200 14702 45000
rect 15842 44200 15898 45000
rect 17038 44200 17094 45000
rect 18234 44200 18290 45000
rect 19430 44200 19486 45000
rect 20626 44200 20682 45000
rect 21822 44200 21878 45000
rect 23018 44200 23074 45000
rect 24214 44200 24270 45000
rect 25410 44200 25466 45000
rect 26606 44200 26662 45000
rect 27802 44200 27858 45000
rect 28998 44200 29054 45000
rect 30194 44200 30250 45000
rect 31390 44200 31446 45000
rect 32586 44200 32642 45000
rect 33782 44200 33838 45000
rect 34978 44200 35034 45000
rect 36174 44200 36230 45000
rect 37370 44200 37426 45000
rect 38566 44200 38622 45000
rect 39762 44200 39818 45000
rect 40958 44200 41014 45000
rect 42154 44200 42210 45000
rect 43350 44200 43406 45000
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 24228 42362 24256 44200
rect 25424 42362 25452 44200
rect 26620 42362 26648 44200
rect 27816 42362 27844 44200
rect 29012 42362 29040 44200
rect 30208 42362 30236 44200
rect 31404 42362 31432 44200
rect 32600 42362 32628 44200
rect 24216 42356 24268 42362
rect 24216 42298 24268 42304
rect 25412 42356 25464 42362
rect 25412 42298 25464 42304
rect 26608 42356 26660 42362
rect 26608 42298 26660 42304
rect 27804 42356 27856 42362
rect 27804 42298 27856 42304
rect 29000 42356 29052 42362
rect 29000 42298 29052 42304
rect 30196 42356 30248 42362
rect 30196 42298 30248 42304
rect 31392 42356 31444 42362
rect 31392 42298 31444 42304
rect 32588 42356 32640 42362
rect 32588 42298 32640 42304
rect 34992 42294 35020 44200
rect 36188 42362 36216 44200
rect 37384 42362 37412 44200
rect 36176 42356 36228 42362
rect 36176 42298 36228 42304
rect 37372 42356 37424 42362
rect 37372 42298 37424 42304
rect 34980 42288 35032 42294
rect 34980 42230 35032 42236
rect 23940 42084 23992 42090
rect 23940 42026 23992 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 940 41608 992 41614
rect 940 41550 992 41556
rect 952 41449 980 41550
rect 938 41440 994 41449
rect 17696 41414 17724 41754
rect 938 41375 994 41384
rect 17328 41386 17724 41414
rect 8116 41064 8168 41070
rect 8116 41006 8168 41012
rect 9128 41064 9180 41070
rect 9128 41006 9180 41012
rect 10048 41064 10100 41070
rect 10048 41006 10100 41012
rect 11152 41064 11204 41070
rect 11152 41006 11204 41012
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 13544 41064 13596 41070
rect 13544 41006 13596 41012
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 940 40520 992 40526
rect 940 40462 992 40468
rect 952 40361 980 40462
rect 8024 40452 8076 40458
rect 8024 40394 8076 40400
rect 938 40352 994 40361
rect 938 40287 994 40296
rect 6276 40044 6328 40050
rect 6276 39986 6328 39992
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 1216 39500 1268 39506
rect 1216 39442 1268 39448
rect 1228 39273 1256 39442
rect 6000 39432 6052 39438
rect 6000 39374 6052 39380
rect 1214 39264 1270 39273
rect 1214 39199 1270 39208
rect 6012 39098 6040 39374
rect 6000 39092 6052 39098
rect 6000 39034 6052 39040
rect 5632 38888 5684 38894
rect 5632 38830 5684 38836
rect 5908 38888 5960 38894
rect 5908 38830 5960 38836
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 1216 38412 1268 38418
rect 1216 38354 1268 38360
rect 1228 38185 1256 38354
rect 4160 38344 4212 38350
rect 4160 38286 4212 38292
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 1214 38176 1270 38185
rect 1214 38111 1270 38120
rect 4172 38010 4200 38286
rect 4712 38208 4764 38214
rect 4712 38150 4764 38156
rect 4160 38004 4212 38010
rect 4160 37946 4212 37952
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4160 37256 4212 37262
rect 4160 37198 4212 37204
rect 1216 37120 1268 37126
rect 1214 37088 1216 37097
rect 1268 37088 1270 37097
rect 1214 37023 1270 37032
rect 4172 36786 4200 37198
rect 4724 37194 4752 38150
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4160 36780 4212 36786
rect 4160 36722 4212 36728
rect 4068 36576 4120 36582
rect 4068 36518 4120 36524
rect 4080 36378 4108 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4908 36378 4936 38286
rect 5448 38208 5500 38214
rect 5448 38150 5500 38156
rect 5264 37800 5316 37806
rect 5264 37742 5316 37748
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 4896 36372 4948 36378
rect 4896 36314 4948 36320
rect 940 36168 992 36174
rect 940 36110 992 36116
rect 4436 36168 4488 36174
rect 4436 36110 4488 36116
rect 952 36009 980 36110
rect 938 36000 994 36009
rect 938 35935 994 35944
rect 4448 35834 4476 36110
rect 4988 36032 5040 36038
rect 4988 35974 5040 35980
rect 4436 35828 4488 35834
rect 4436 35770 4488 35776
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34921 980 35022
rect 5000 35018 5028 35974
rect 5276 35630 5304 37742
rect 5460 36854 5488 38150
rect 5644 38010 5672 38830
rect 5632 38004 5684 38010
rect 5632 37946 5684 37952
rect 5920 37806 5948 38830
rect 6184 38752 6236 38758
rect 6184 38694 6236 38700
rect 6196 38010 6224 38694
rect 6184 38004 6236 38010
rect 6184 37946 6236 37952
rect 5908 37800 5960 37806
rect 5908 37742 5960 37748
rect 5632 37732 5684 37738
rect 5632 37674 5684 37680
rect 5644 37466 5672 37674
rect 5632 37460 5684 37466
rect 5632 37402 5684 37408
rect 5448 36848 5500 36854
rect 5448 36790 5500 36796
rect 5644 36786 5672 37402
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5632 36372 5684 36378
rect 5632 36314 5684 36320
rect 5644 36242 5672 36314
rect 5632 36236 5684 36242
rect 5552 36196 5632 36224
rect 5264 35624 5316 35630
rect 5264 35566 5316 35572
rect 4988 35012 5040 35018
rect 4988 34954 5040 34960
rect 3332 34944 3384 34950
rect 938 34912 994 34921
rect 3332 34886 3384 34892
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 938 34847 994 34856
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 2136 34536 2188 34542
rect 2136 34478 2188 34484
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2872 34536 2924 34542
rect 2872 34478 2924 34484
rect 940 33992 992 33998
rect 940 33934 992 33940
rect 952 33833 980 33934
rect 938 33824 994 33833
rect 938 33759 994 33768
rect 1780 32978 1808 34478
rect 2148 34202 2176 34478
rect 2136 34196 2188 34202
rect 2136 34138 2188 34144
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1964 33658 1992 34002
rect 2044 33992 2096 33998
rect 2044 33934 2096 33940
rect 2056 33658 2084 33934
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 2044 33652 2096 33658
rect 2044 33594 2096 33600
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1768 32972 1820 32978
rect 1768 32914 1820 32920
rect 1872 32910 1900 33390
rect 1860 32904 1912 32910
rect 2240 32858 2268 34478
rect 2596 33856 2648 33862
rect 2596 33798 2648 33804
rect 2608 33658 2636 33798
rect 2596 33652 2648 33658
rect 2596 33594 2648 33600
rect 2884 33114 2912 34478
rect 3344 34066 3372 34886
rect 3516 34536 3568 34542
rect 3516 34478 3568 34484
rect 3424 34400 3476 34406
rect 3424 34342 3476 34348
rect 3332 34060 3384 34066
rect 3332 34002 3384 34008
rect 3436 33930 3464 34342
rect 3424 33924 3476 33930
rect 3424 33866 3476 33872
rect 3528 33658 3556 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 34202 4660 34886
rect 4712 34740 4764 34746
rect 4712 34682 4764 34688
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 3608 33856 3660 33862
rect 3608 33798 3660 33804
rect 3884 33856 3936 33862
rect 3884 33798 3936 33804
rect 3516 33652 3568 33658
rect 3516 33594 3568 33600
rect 3424 33312 3476 33318
rect 3424 33254 3476 33260
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2686 33008 2742 33017
rect 2686 32943 2742 32952
rect 2700 32910 2728 32943
rect 1860 32846 1912 32852
rect 940 32768 992 32774
rect 938 32736 940 32745
rect 992 32736 994 32745
rect 938 32671 994 32680
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1504 31657 1532 32302
rect 1490 31648 1546 31657
rect 1490 31583 1546 31592
rect 1216 30796 1268 30802
rect 1216 30738 1268 30744
rect 1228 30569 1256 30738
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 1214 30560 1270 30569
rect 1214 30495 1270 30504
rect 1596 29782 1624 30670
rect 1584 29776 1636 29782
rect 1584 29718 1636 29724
rect 1216 29708 1268 29714
rect 1216 29650 1268 29656
rect 1228 29481 1256 29650
rect 1214 29472 1270 29481
rect 1214 29407 1270 29416
rect 1490 29200 1546 29209
rect 1490 29135 1546 29144
rect 1504 29034 1532 29135
rect 1492 29028 1544 29034
rect 1492 28970 1544 28976
rect 1216 28620 1268 28626
rect 1216 28562 1268 28568
rect 1228 28393 1256 28562
rect 1214 28384 1270 28393
rect 1214 28319 1270 28328
rect 1216 27532 1268 27538
rect 1216 27474 1268 27480
rect 1228 27305 1256 27474
rect 1214 27296 1270 27305
rect 1214 27231 1270 27240
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 1412 25294 1440 25774
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1504 25158 1532 28970
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1596 28121 1624 28494
rect 1582 28112 1638 28121
rect 1582 28047 1638 28056
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 26518 1624 27270
rect 1688 27169 1716 32370
rect 1872 32026 1900 32846
rect 2148 32842 2268 32858
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2136 32836 2268 32842
rect 2188 32830 2268 32836
rect 2136 32778 2188 32784
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 1860 32020 1912 32026
rect 1860 31962 1912 31968
rect 1872 31754 1900 31962
rect 1872 31726 1992 31754
rect 1964 31346 1992 31726
rect 2976 31482 3004 32302
rect 3436 31754 3464 33254
rect 3516 32224 3568 32230
rect 3516 32166 3568 32172
rect 3528 32026 3556 32166
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3424 31748 3476 31754
rect 3424 31690 3476 31696
rect 2964 31476 3016 31482
rect 2964 31418 3016 31424
rect 3148 31408 3200 31414
rect 3148 31350 3200 31356
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 2504 31340 2556 31346
rect 2504 31282 2556 31288
rect 2516 30938 2544 31282
rect 2504 30932 2556 30938
rect 2504 30874 2556 30880
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 2056 30394 2084 30738
rect 3056 30592 3108 30598
rect 2870 30560 2926 30569
rect 3056 30534 3108 30540
rect 2870 30495 2926 30504
rect 2044 30388 2096 30394
rect 2044 30330 2096 30336
rect 2884 30258 2912 30495
rect 2962 30424 3018 30433
rect 2962 30359 3018 30368
rect 2136 30252 2188 30258
rect 2136 30194 2188 30200
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2504 30252 2556 30258
rect 2504 30194 2556 30200
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1860 29504 1912 29510
rect 1860 29446 1912 29452
rect 1872 29238 1900 29446
rect 1860 29232 1912 29238
rect 1860 29174 1912 29180
rect 1768 28960 1820 28966
rect 1768 28902 1820 28908
rect 1780 28218 1808 28902
rect 1860 28416 1912 28422
rect 1860 28358 1912 28364
rect 1872 28218 1900 28358
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 1872 28082 1900 28154
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 2056 27606 2084 29582
rect 2148 28014 2176 30194
rect 2424 29646 2452 30194
rect 2516 29850 2544 30194
rect 2688 30116 2740 30122
rect 2688 30058 2740 30064
rect 2504 29844 2556 29850
rect 2504 29786 2556 29792
rect 2700 29714 2728 30058
rect 2976 30054 3004 30359
rect 2964 30048 3016 30054
rect 2964 29990 3016 29996
rect 3068 29866 3096 30534
rect 3160 30258 3188 31350
rect 3424 30728 3476 30734
rect 3330 30696 3386 30705
rect 3424 30670 3476 30676
rect 3330 30631 3332 30640
rect 3384 30631 3386 30640
rect 3332 30602 3384 30608
rect 3344 30394 3372 30602
rect 3332 30388 3384 30394
rect 3332 30330 3384 30336
rect 3240 30320 3292 30326
rect 3240 30262 3292 30268
rect 3148 30252 3200 30258
rect 3148 30194 3200 30200
rect 2884 29838 3096 29866
rect 2688 29708 2740 29714
rect 2688 29650 2740 29656
rect 2412 29640 2464 29646
rect 2412 29582 2464 29588
rect 2780 29504 2832 29510
rect 2780 29446 2832 29452
rect 2318 29336 2374 29345
rect 2318 29271 2374 29280
rect 2688 29300 2740 29306
rect 2332 29034 2360 29271
rect 2688 29242 2740 29248
rect 2504 29096 2556 29102
rect 2504 29038 2556 29044
rect 2596 29096 2648 29102
rect 2596 29038 2648 29044
rect 2320 29028 2372 29034
rect 2320 28970 2372 28976
rect 2228 28960 2280 28966
rect 2228 28902 2280 28908
rect 2412 28960 2464 28966
rect 2412 28902 2464 28908
rect 2240 28801 2268 28902
rect 2226 28792 2282 28801
rect 2226 28727 2282 28736
rect 2424 28218 2452 28902
rect 2516 28762 2544 29038
rect 2504 28756 2556 28762
rect 2504 28698 2556 28704
rect 2608 28558 2636 29038
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 2136 28008 2188 28014
rect 2136 27950 2188 27956
rect 2504 28008 2556 28014
rect 2504 27950 2556 27956
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 2516 27334 2544 27950
rect 2700 27878 2728 29242
rect 2792 28966 2820 29446
rect 2780 28960 2832 28966
rect 2780 28902 2832 28908
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 1674 27160 1730 27169
rect 2884 27130 2912 29838
rect 2964 29776 3016 29782
rect 2964 29718 3016 29724
rect 2976 27985 3004 29718
rect 3160 29696 3188 30194
rect 3252 29850 3280 30262
rect 3332 30116 3384 30122
rect 3332 30058 3384 30064
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3160 29668 3280 29696
rect 3252 29492 3280 29668
rect 3344 29646 3372 30058
rect 3436 29850 3464 30670
rect 3516 30252 3568 30258
rect 3516 30194 3568 30200
rect 3424 29844 3476 29850
rect 3424 29786 3476 29792
rect 3528 29714 3556 30194
rect 3516 29708 3568 29714
rect 3516 29650 3568 29656
rect 3332 29640 3384 29646
rect 3332 29582 3384 29588
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3436 29492 3464 29582
rect 3054 29472 3110 29481
rect 3252 29464 3464 29492
rect 3054 29407 3110 29416
rect 3068 29170 3096 29407
rect 3330 29336 3386 29345
rect 3386 29294 3464 29322
rect 3330 29271 3386 29280
rect 3332 29232 3384 29238
rect 3332 29174 3384 29180
rect 3056 29164 3108 29170
rect 3056 29106 3108 29112
rect 3068 28558 3096 29106
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3056 28552 3108 28558
rect 3056 28494 3108 28500
rect 3056 28144 3108 28150
rect 3160 28132 3188 28970
rect 3252 28422 3280 29038
rect 3344 28966 3372 29174
rect 3436 29102 3464 29294
rect 3528 29288 3556 29650
rect 3620 29458 3648 33798
rect 3896 33386 3924 33798
rect 4080 33454 4108 34002
rect 4724 33522 4752 34682
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 5000 34134 5028 34546
rect 5356 34400 5408 34406
rect 5356 34342 5408 34348
rect 4988 34128 5040 34134
rect 4988 34070 5040 34076
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4896 33448 4948 33454
rect 4896 33390 4948 33396
rect 3884 33380 3936 33386
rect 3884 33322 3936 33328
rect 3988 33114 4016 33390
rect 3976 33108 4028 33114
rect 3976 33050 4028 33056
rect 4080 32774 4108 33390
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4528 32904 4580 32910
rect 4580 32864 4660 32892
rect 4528 32846 4580 32852
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 3988 31754 4016 32710
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 4080 32008 4108 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4080 31980 4200 32008
rect 4172 31929 4200 31980
rect 4158 31920 4214 31929
rect 4158 31855 4214 31864
rect 4344 31884 4396 31890
rect 4172 31754 4200 31855
rect 4344 31826 4396 31832
rect 3896 31726 4016 31754
rect 4160 31748 4212 31754
rect 3896 31686 3924 31726
rect 4160 31690 4212 31696
rect 3884 31680 3936 31686
rect 3884 31622 3936 31628
rect 3896 31346 3924 31622
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 3700 31136 3752 31142
rect 3700 31078 3752 31084
rect 3712 30734 3740 31078
rect 3700 30728 3752 30734
rect 3752 30688 3832 30716
rect 3700 30670 3752 30676
rect 3620 29430 3740 29458
rect 3608 29300 3660 29306
rect 3528 29260 3608 29288
rect 3608 29242 3660 29248
rect 3424 29096 3476 29102
rect 3424 29038 3476 29044
rect 3332 28960 3384 28966
rect 3332 28902 3384 28908
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3344 28472 3372 28902
rect 3436 28762 3464 28902
rect 3712 28762 3740 29430
rect 3424 28756 3476 28762
rect 3424 28698 3476 28704
rect 3700 28756 3752 28762
rect 3700 28698 3752 28704
rect 3606 28656 3662 28665
rect 3606 28591 3662 28600
rect 3424 28484 3476 28490
rect 3344 28444 3424 28472
rect 3424 28426 3476 28432
rect 3240 28416 3292 28422
rect 3238 28384 3240 28393
rect 3292 28384 3294 28393
rect 3238 28319 3294 28328
rect 3252 28150 3280 28319
rect 3108 28104 3188 28132
rect 3240 28144 3292 28150
rect 3056 28086 3108 28092
rect 3240 28086 3292 28092
rect 2962 27976 3018 27985
rect 2962 27911 3018 27920
rect 3148 27872 3200 27878
rect 3148 27814 3200 27820
rect 3160 27470 3188 27814
rect 3332 27600 3384 27606
rect 3332 27542 3384 27548
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 1674 27095 1730 27104
rect 2872 27124 2924 27130
rect 2924 27084 3004 27112
rect 2872 27066 2924 27072
rect 1860 26920 1912 26926
rect 1860 26862 1912 26868
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1584 26376 1636 26382
rect 1582 26344 1584 26353
rect 1636 26344 1638 26353
rect 1582 26279 1638 26288
rect 1872 26217 1900 26862
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 1858 26208 1914 26217
rect 1858 26143 1914 26152
rect 2688 25356 2740 25362
rect 2688 25298 2740 25304
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1768 25220 1820 25226
rect 1768 25162 1820 25168
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 24750 1532 25094
rect 1780 24954 1808 25162
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 2056 24886 2084 25230
rect 2044 24880 2096 24886
rect 2044 24822 2096 24828
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1216 24268 1268 24274
rect 1216 24210 1268 24216
rect 1228 24041 1256 24210
rect 1214 24032 1270 24041
rect 1214 23967 1270 23976
rect 1216 23180 1268 23186
rect 1216 23122 1268 23128
rect 1228 22953 1256 23122
rect 1214 22944 1270 22953
rect 1214 22879 1270 22888
rect 1216 22092 1268 22098
rect 1216 22034 1268 22040
rect 1228 21865 1256 22034
rect 1214 21856 1270 21865
rect 1214 21791 1270 21800
rect 1216 21004 1268 21010
rect 1216 20946 1268 20952
rect 1228 20777 1256 20946
rect 1214 20768 1270 20777
rect 1214 20703 1270 20712
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 1228 19689 1256 19858
rect 1214 19680 1270 19689
rect 1214 19615 1270 19624
rect 1504 19310 1532 24686
rect 1582 24304 1638 24313
rect 1582 24239 1638 24248
rect 1596 24206 1624 24239
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 2056 23662 2084 24822
rect 2596 24676 2648 24682
rect 2596 24618 2648 24624
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1768 23656 1820 23662
rect 1768 23598 1820 23604
rect 2044 23656 2096 23662
rect 2044 23598 2096 23604
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1596 22030 1624 22918
rect 1780 22438 1808 23598
rect 2148 23050 2176 23666
rect 2136 23044 2188 23050
rect 2136 22986 2188 22992
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1780 21332 1808 22374
rect 2042 22128 2098 22137
rect 2042 22063 2098 22072
rect 1952 21616 2004 21622
rect 1950 21584 1952 21593
rect 2004 21584 2006 21593
rect 1950 21519 2006 21528
rect 1860 21344 1912 21350
rect 1780 21304 1860 21332
rect 1860 21286 1912 21292
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20466 1716 20810
rect 1872 20466 1900 21286
rect 1964 20942 1992 21519
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1216 18692 1268 18698
rect 1216 18634 1268 18640
rect 1228 18601 1256 18634
rect 1214 18592 1270 18601
rect 1214 18527 1270 18536
rect 1780 18290 1808 19246
rect 1872 18834 1900 20402
rect 1860 18828 1912 18834
rect 1860 18770 1912 18776
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17513 1256 17682
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1214 17504 1270 17513
rect 1214 17439 1270 17448
rect 1688 17338 1716 17614
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1780 17134 1808 18226
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1216 16516 1268 16522
rect 1216 16458 1268 16464
rect 1228 16425 1256 16458
rect 1214 16416 1270 16425
rect 1214 16351 1270 16360
rect 1676 16108 1728 16114
rect 1780 16096 1808 17070
rect 1860 16108 1912 16114
rect 1780 16068 1860 16096
rect 1676 16050 1728 16056
rect 1860 16050 1912 16056
rect 1216 15564 1268 15570
rect 1216 15506 1268 15512
rect 1228 15337 1256 15506
rect 1214 15328 1270 15337
rect 1214 15263 1270 15272
rect 1688 15162 1716 16050
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1216 14476 1268 14482
rect 1216 14418 1268 14424
rect 1228 14249 1256 14418
rect 1214 14240 1270 14249
rect 1214 14175 1270 14184
rect 1688 14074 1716 15098
rect 2056 15094 2084 22063
rect 2424 21622 2452 22374
rect 2412 21616 2464 21622
rect 2412 21558 2464 21564
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2148 21146 2176 21422
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 2516 21049 2544 21286
rect 2502 21040 2558 21049
rect 2502 20975 2558 20984
rect 2502 20768 2558 20777
rect 2502 20703 2558 20712
rect 2044 15088 2096 15094
rect 2044 15030 2096 15036
rect 2516 14074 2544 20703
rect 2608 18358 2636 24618
rect 2700 18766 2728 25298
rect 2792 25129 2820 26250
rect 2778 25120 2834 25129
rect 2778 25055 2834 25064
rect 2872 24608 2924 24614
rect 2872 24550 2924 24556
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2792 21146 2820 24210
rect 2884 23322 2912 24550
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2976 22953 3004 27084
rect 3344 26217 3372 27542
rect 3436 27130 3464 28426
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 3330 26208 3386 26217
rect 3330 26143 3386 26152
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 3252 25498 3280 25842
rect 3240 25492 3292 25498
rect 3240 25434 3292 25440
rect 3332 25424 3384 25430
rect 3332 25366 3384 25372
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3068 24410 3096 25230
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 3068 23089 3096 24074
rect 3344 23730 3372 25366
rect 3436 25265 3464 26930
rect 3528 26926 3556 28018
rect 3516 26920 3568 26926
rect 3516 26862 3568 26868
rect 3422 25256 3478 25265
rect 3422 25191 3478 25200
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3054 23080 3110 23089
rect 3054 23015 3110 23024
rect 3068 22982 3096 23015
rect 3056 22976 3108 22982
rect 2962 22944 3018 22953
rect 3056 22918 3108 22924
rect 2962 22879 3018 22888
rect 3160 22778 3188 23666
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3252 23118 3280 23530
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 3344 23322 3372 23462
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 3330 23216 3386 23225
rect 3330 23151 3386 23160
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3054 22672 3110 22681
rect 3054 22607 3110 22616
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 2884 21690 2912 22170
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2976 21146 3004 22510
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2792 20398 2820 21082
rect 3068 20482 3096 22607
rect 3148 22500 3200 22506
rect 3148 22442 3200 22448
rect 3160 20584 3188 22442
rect 3252 20942 3280 22918
rect 3344 20942 3372 23151
rect 3436 22098 3464 25094
rect 3620 24936 3648 28591
rect 3712 27470 3740 28698
rect 3804 28626 3832 30688
rect 3792 28620 3844 28626
rect 3792 28562 3844 28568
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3804 28218 3832 28426
rect 3896 28234 3924 31282
rect 4356 31278 4384 31826
rect 4632 31754 4660 32864
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 4724 32026 4752 32778
rect 4908 32026 4936 33390
rect 5368 33318 5396 34342
rect 5552 34134 5580 36196
rect 5632 36178 5684 36184
rect 5632 35760 5684 35766
rect 5632 35702 5684 35708
rect 5644 35290 5672 35702
rect 5632 35284 5684 35290
rect 5632 35226 5684 35232
rect 5540 34128 5592 34134
rect 5540 34070 5592 34076
rect 5448 33856 5500 33862
rect 5448 33798 5500 33804
rect 5460 33658 5488 33798
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5356 33312 5408 33318
rect 5356 33254 5408 33260
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5368 32026 5396 32710
rect 5644 32434 5672 33254
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 4896 32020 4948 32026
rect 4896 31962 4948 31968
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 5368 31890 5396 31962
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 4632 31726 4752 31754
rect 4344 31272 4396 31278
rect 4344 31214 4396 31220
rect 4068 31204 4120 31210
rect 4068 31146 4120 31152
rect 4080 30938 4108 31146
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 3988 30734 4016 30874
rect 4632 30734 4660 31078
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4540 30598 4568 30670
rect 3976 30592 4028 30598
rect 3976 30534 4028 30540
rect 4528 30592 4580 30598
rect 4528 30534 4580 30540
rect 3988 30326 4016 30534
rect 4724 30326 4752 31726
rect 4908 31346 4936 31826
rect 4988 31680 5040 31686
rect 4988 31622 5040 31628
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 5000 31346 5028 31622
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4816 30938 4844 31214
rect 5000 30938 5028 31282
rect 4804 30932 4856 30938
rect 4804 30874 4856 30880
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 4896 30728 4948 30734
rect 4894 30696 4896 30705
rect 4988 30728 5040 30734
rect 4948 30696 4950 30705
rect 4988 30670 5040 30676
rect 4894 30631 4950 30640
rect 4802 30424 4858 30433
rect 4802 30359 4804 30368
rect 4856 30359 4858 30368
rect 4804 30330 4856 30336
rect 3976 30320 4028 30326
rect 3976 30262 4028 30268
rect 4160 30320 4212 30326
rect 4344 30320 4396 30326
rect 4160 30262 4212 30268
rect 4264 30280 4344 30308
rect 4172 30190 4200 30262
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4172 30054 4200 30126
rect 4264 30122 4292 30280
rect 4712 30320 4764 30326
rect 4344 30262 4396 30268
rect 4526 30288 4582 30297
rect 5000 30297 5028 30670
rect 5184 30433 5212 31622
rect 5460 31414 5488 31826
rect 5448 31408 5500 31414
rect 5448 31350 5500 31356
rect 5538 31376 5594 31385
rect 5460 30870 5488 31350
rect 5538 31311 5594 31320
rect 5552 31278 5580 31311
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5448 30864 5500 30870
rect 5448 30806 5500 30812
rect 5540 30864 5592 30870
rect 5540 30806 5592 30812
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 5170 30424 5226 30433
rect 5170 30359 5226 30368
rect 5276 30326 5304 30602
rect 5264 30320 5316 30326
rect 4712 30262 4764 30268
rect 4986 30288 5042 30297
rect 4526 30223 4582 30232
rect 4540 30190 4568 30223
rect 4528 30184 4580 30190
rect 4528 30126 4580 30132
rect 4252 30116 4304 30122
rect 4252 30058 4304 30064
rect 4620 30116 4672 30122
rect 4620 30058 4672 30064
rect 4160 30048 4212 30054
rect 3988 30008 4160 30036
rect 3988 29714 4016 30008
rect 4160 29990 4212 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4066 29744 4122 29753
rect 3976 29708 4028 29714
rect 4066 29679 4122 29688
rect 3976 29650 4028 29656
rect 3976 29504 4028 29510
rect 3976 29446 4028 29452
rect 3988 29186 4016 29446
rect 4080 29306 4108 29679
rect 4632 29306 4660 30058
rect 4724 29850 4752 30262
rect 4896 30252 4948 30258
rect 5264 30262 5316 30268
rect 4986 30223 5042 30232
rect 4896 30194 4948 30200
rect 4908 30036 4936 30194
rect 5368 30190 5396 30670
rect 5446 30560 5502 30569
rect 5446 30495 5502 30504
rect 5460 30394 5488 30495
rect 5448 30388 5500 30394
rect 5448 30330 5500 30336
rect 5172 30184 5224 30190
rect 5172 30126 5224 30132
rect 5356 30184 5408 30190
rect 5356 30126 5408 30132
rect 4908 30008 5120 30036
rect 4712 29844 4764 29850
rect 4712 29786 4764 29792
rect 4724 29646 4752 29786
rect 4712 29640 4764 29646
rect 4712 29582 4764 29588
rect 5092 29578 5120 30008
rect 5184 29850 5212 30126
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 5276 29730 5304 29990
rect 5368 29753 5396 30126
rect 5552 30122 5580 30806
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5644 30394 5672 30670
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 5540 30116 5592 30122
rect 5540 30058 5592 30064
rect 5184 29702 5304 29730
rect 5354 29744 5410 29753
rect 5080 29572 5132 29578
rect 5080 29514 5132 29520
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4620 29300 4672 29306
rect 4620 29242 4672 29248
rect 4526 29200 4582 29209
rect 3988 29158 4108 29186
rect 3974 28792 4030 28801
rect 3974 28727 3976 28736
rect 4028 28727 4030 28736
rect 3976 28698 4028 28704
rect 4080 28404 4108 29158
rect 4526 29135 4528 29144
rect 4580 29135 4582 29144
rect 4528 29106 4580 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4344 28620 4396 28626
rect 4344 28562 4396 28568
rect 4160 28416 4212 28422
rect 4080 28376 4160 28404
rect 4160 28358 4212 28364
rect 3974 28248 4030 28257
rect 3792 28212 3844 28218
rect 3896 28206 3974 28234
rect 4356 28218 4384 28562
rect 4434 28520 4490 28529
rect 4434 28455 4436 28464
rect 4488 28455 4490 28464
rect 4436 28426 4488 28432
rect 3974 28183 4030 28192
rect 4068 28212 4120 28218
rect 3792 28154 3844 28160
rect 4068 28154 4120 28160
rect 4344 28212 4396 28218
rect 4344 28154 4396 28160
rect 3804 27674 3832 28154
rect 3884 27940 3936 27946
rect 3884 27882 3936 27888
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 3896 27470 3924 27882
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3792 26988 3844 26994
rect 3896 26976 3924 27406
rect 4080 26994 4108 28154
rect 4632 28064 4660 29242
rect 4712 29164 4764 29170
rect 4712 29106 4764 29112
rect 4724 28218 4752 29106
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4816 28801 4844 28902
rect 4802 28792 4858 28801
rect 4802 28727 4858 28736
rect 4908 28744 4936 29446
rect 5092 29306 5120 29514
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4986 29200 5042 29209
rect 4986 29135 4988 29144
rect 5040 29135 5042 29144
rect 4988 29106 5040 29112
rect 5080 28756 5132 28762
rect 4908 28716 5080 28744
rect 4908 28490 4936 28716
rect 5080 28698 5132 28704
rect 5184 28506 5212 29702
rect 5354 29679 5410 29688
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 5276 29306 5304 29582
rect 5264 29300 5316 29306
rect 5264 29242 5316 29248
rect 5448 29164 5500 29170
rect 5448 29106 5500 29112
rect 5460 28762 5488 29106
rect 5630 28792 5686 28801
rect 5448 28756 5500 28762
rect 5630 28727 5632 28736
rect 5448 28698 5500 28704
rect 5684 28727 5686 28736
rect 5632 28698 5684 28704
rect 5460 28558 5488 28698
rect 4896 28484 4948 28490
rect 4896 28426 4948 28432
rect 5000 28478 5212 28506
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5264 28484 5316 28490
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4540 28036 4660 28064
rect 4540 27946 4568 28036
rect 4804 28008 4856 28014
rect 4724 27968 4804 27996
rect 4528 27940 4580 27946
rect 4528 27882 4580 27888
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 4172 27130 4200 27610
rect 4344 27532 4396 27538
rect 4344 27474 4396 27480
rect 4356 27402 4384 27474
rect 4344 27396 4396 27402
rect 4344 27338 4396 27344
rect 4436 27396 4488 27402
rect 4436 27338 4488 27344
rect 4252 27328 4304 27334
rect 4252 27270 4304 27276
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3844 26948 3924 26976
rect 4068 26988 4120 26994
rect 3792 26930 3844 26936
rect 4068 26930 4120 26936
rect 4264 26908 4292 27270
rect 4356 27033 4384 27338
rect 4448 27062 4476 27338
rect 4436 27056 4488 27062
rect 4342 27024 4398 27033
rect 4436 26998 4488 27004
rect 4342 26959 4398 26968
rect 4344 26920 4396 26926
rect 4264 26888 4344 26908
rect 4396 26888 4398 26897
rect 4264 26880 4342 26888
rect 4632 26874 4660 27882
rect 4724 27470 4752 27968
rect 4804 27950 4856 27956
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4724 27062 4752 27406
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 4816 27130 4844 27338
rect 4804 27124 4856 27130
rect 4804 27066 4856 27072
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4802 27024 4858 27033
rect 4802 26959 4804 26968
rect 4856 26959 4858 26968
rect 4804 26930 4856 26936
rect 4632 26858 4844 26874
rect 4632 26852 4856 26858
rect 4632 26846 4804 26852
rect 4342 26823 4398 26832
rect 4804 26794 4856 26800
rect 4816 26761 4844 26794
rect 4802 26752 4858 26761
rect 4214 26684 4522 26693
rect 4802 26687 4858 26696
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4436 26512 4488 26518
rect 4436 26454 4488 26460
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3700 26240 3752 26246
rect 3700 26182 3752 26188
rect 3712 25974 3740 26182
rect 3700 25968 3752 25974
rect 3700 25910 3752 25916
rect 3712 25498 3740 25910
rect 3700 25492 3752 25498
rect 3700 25434 3752 25440
rect 3528 24908 3648 24936
rect 3528 24274 3556 24908
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3620 24410 3648 24754
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3516 24268 3568 24274
rect 3568 24228 3648 24256
rect 3516 24210 3568 24216
rect 3620 23186 3648 24228
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3528 21486 3556 22918
rect 3712 22574 3740 24754
rect 3804 23730 3832 26250
rect 3896 26042 3924 26318
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3896 25430 3924 25842
rect 3988 25702 4016 26250
rect 4356 25906 4384 26386
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 4448 25809 4476 26454
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 4620 25832 4672 25838
rect 4434 25800 4490 25809
rect 4620 25774 4672 25780
rect 4434 25735 4490 25744
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3884 25424 3936 25430
rect 3884 25366 3936 25372
rect 3988 25294 4016 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3896 24206 3924 24346
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3792 23724 3844 23730
rect 3844 23684 3924 23712
rect 3792 23666 3844 23672
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3606 21992 3662 22001
rect 3606 21927 3662 21936
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3436 20806 3464 21286
rect 3620 21010 3648 21927
rect 3712 21690 3740 22102
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3608 21004 3660 21010
rect 3528 20964 3608 20992
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3160 20556 3372 20584
rect 2964 20460 3016 20466
rect 3068 20454 3188 20482
rect 2964 20402 3016 20408
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2976 20058 3004 20402
rect 3054 20360 3110 20369
rect 3054 20295 3110 20304
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3068 19922 3096 20295
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3068 19514 3096 19858
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3054 19272 3110 19281
rect 3054 19207 3110 19216
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2884 17134 2912 19110
rect 3068 18426 3096 19207
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3068 18306 3096 18362
rect 2976 18278 3096 18306
rect 2976 17746 3004 18278
rect 3160 18170 3188 20454
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3252 19922 3280 20198
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3344 19514 3372 20556
rect 3424 20528 3476 20534
rect 3422 20496 3424 20505
rect 3476 20496 3478 20505
rect 3422 20431 3478 20440
rect 3332 19508 3384 19514
rect 3528 19496 3556 20964
rect 3608 20946 3660 20952
rect 3804 20942 3832 22986
rect 3896 22778 3924 23684
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3988 22710 4016 25230
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 4080 24206 4108 25094
rect 4632 24818 4660 25774
rect 4724 25362 4752 25842
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4724 24993 4752 25298
rect 4710 24984 4766 24993
rect 4710 24919 4766 24928
rect 4816 24818 4844 26522
rect 4908 26042 4936 28426
rect 5000 28422 5028 28478
rect 5264 28426 5316 28432
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 5080 28416 5132 28422
rect 5080 28358 5132 28364
rect 5172 28416 5224 28422
rect 5172 28358 5224 28364
rect 5092 27674 5120 28358
rect 5184 28218 5212 28358
rect 5172 28212 5224 28218
rect 5172 28154 5224 28160
rect 5276 28064 5304 28426
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5368 28082 5396 28358
rect 5460 28218 5488 28494
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5184 28036 5304 28064
rect 5356 28076 5408 28082
rect 5080 27668 5132 27674
rect 5080 27610 5132 27616
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 5000 27130 5028 27406
rect 5184 27282 5212 28036
rect 5356 28018 5408 28024
rect 5552 28014 5580 28494
rect 5632 28416 5684 28422
rect 5630 28384 5632 28393
rect 5684 28384 5686 28393
rect 5630 28319 5686 28328
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5264 27872 5316 27878
rect 5264 27814 5316 27820
rect 5448 27872 5500 27878
rect 5552 27849 5580 27950
rect 5448 27814 5500 27820
rect 5538 27840 5594 27849
rect 5276 27470 5304 27814
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5262 27296 5318 27305
rect 5184 27254 5262 27282
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 5184 26994 5212 27254
rect 5262 27231 5318 27240
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5264 26988 5316 26994
rect 5264 26930 5316 26936
rect 4988 26920 5040 26926
rect 5040 26868 5212 26874
rect 4988 26862 5212 26868
rect 5000 26858 5212 26862
rect 5000 26852 5224 26858
rect 5000 26846 5172 26852
rect 5172 26794 5224 26800
rect 5276 26761 5304 26930
rect 5368 26897 5396 27542
rect 5460 26926 5488 27814
rect 5538 27775 5594 27784
rect 5644 27674 5672 28018
rect 5632 27668 5684 27674
rect 5632 27610 5684 27616
rect 5644 27470 5672 27610
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5540 27396 5592 27402
rect 5540 27338 5592 27344
rect 5552 27305 5580 27338
rect 5632 27328 5684 27334
rect 5538 27296 5594 27305
rect 5632 27270 5684 27276
rect 5538 27231 5594 27240
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5448 26920 5500 26926
rect 5354 26888 5410 26897
rect 5448 26862 5500 26868
rect 5354 26823 5410 26832
rect 5262 26752 5318 26761
rect 5262 26687 5318 26696
rect 4988 26512 5040 26518
rect 5172 26512 5224 26518
rect 4988 26454 5040 26460
rect 5170 26480 5172 26489
rect 5224 26480 5226 26489
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 5000 25906 5028 26454
rect 5170 26415 5226 26424
rect 5184 26382 5212 26415
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5092 26042 5120 26318
rect 5172 26240 5224 26246
rect 5224 26200 5304 26228
rect 5172 26182 5224 26188
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5092 25906 5120 25978
rect 5172 25968 5224 25974
rect 5276 25945 5304 26200
rect 5172 25910 5224 25916
rect 5262 25936 5318 25945
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5000 25226 5028 25842
rect 5080 25696 5132 25702
rect 5080 25638 5132 25644
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4896 25152 4948 25158
rect 5092 25106 5120 25638
rect 5184 25537 5212 25910
rect 5262 25871 5264 25880
rect 5316 25871 5318 25880
rect 5264 25842 5316 25848
rect 5170 25528 5226 25537
rect 5276 25498 5304 25842
rect 5170 25463 5226 25472
rect 5264 25492 5316 25498
rect 5184 25294 5212 25463
rect 5264 25434 5316 25440
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 4896 25094 4948 25100
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4528 24744 4580 24750
rect 4618 24712 4674 24721
rect 4580 24692 4618 24698
rect 4528 24686 4618 24692
rect 4540 24670 4618 24686
rect 4618 24647 4674 24656
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4528 24336 4580 24342
rect 4528 24278 4580 24284
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4080 23866 4108 24006
rect 4158 23896 4214 23905
rect 4068 23860 4120 23866
rect 4158 23831 4214 23840
rect 4068 23802 4120 23808
rect 4172 23662 4200 23831
rect 4160 23656 4212 23662
rect 4540 23633 4568 24278
rect 4724 24274 4752 24550
rect 4712 24268 4764 24274
rect 4632 24228 4712 24256
rect 4160 23598 4212 23604
rect 4526 23624 4582 23633
rect 4526 23559 4582 23568
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4080 23118 4108 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 24228
rect 4712 24210 4764 24216
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4724 23361 4752 23802
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4710 23352 4766 23361
rect 4710 23287 4766 23296
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3896 21729 3924 22578
rect 4264 22545 4292 22918
rect 4250 22536 4306 22545
rect 4068 22500 4120 22506
rect 4250 22471 4306 22480
rect 4068 22442 4120 22448
rect 3882 21720 3938 21729
rect 3882 21655 3938 21664
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3792 20936 3844 20942
rect 3698 20904 3754 20913
rect 3792 20878 3844 20884
rect 3698 20839 3754 20848
rect 3712 20534 3740 20839
rect 3896 20534 3924 21422
rect 4080 20942 4108 22442
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22166 4660 22986
rect 4724 22234 4752 23054
rect 4816 22817 4844 23598
rect 4802 22808 4858 22817
rect 4802 22743 4858 22752
rect 4816 22642 4844 22743
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4908 22522 4936 25094
rect 5000 25078 5120 25106
rect 5000 24410 5028 25078
rect 5184 24954 5212 25230
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 5092 24290 5120 24822
rect 5276 24818 5304 25094
rect 5368 24954 5396 26823
rect 5460 26790 5488 26862
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5460 25498 5488 26726
rect 5552 26246 5580 26930
rect 5644 26586 5672 27270
rect 5736 26994 5764 37130
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5828 34490 5856 37062
rect 5920 36106 5948 37742
rect 6288 37670 6316 39986
rect 6736 39976 6788 39982
rect 6736 39918 6788 39924
rect 6368 39500 6420 39506
rect 6368 39442 6420 39448
rect 6380 37806 6408 39442
rect 6552 39296 6604 39302
rect 6552 39238 6604 39244
rect 6564 38282 6592 39238
rect 6748 38554 6776 39918
rect 7104 39840 7156 39846
rect 7104 39782 7156 39788
rect 7840 39840 7892 39846
rect 7840 39782 7892 39788
rect 7116 39098 7144 39782
rect 7380 39500 7432 39506
rect 7380 39442 7432 39448
rect 7104 39092 7156 39098
rect 7104 39034 7156 39040
rect 7392 38894 7420 39442
rect 7380 38888 7432 38894
rect 7380 38830 7432 38836
rect 7104 38752 7156 38758
rect 7104 38694 7156 38700
rect 6736 38548 6788 38554
rect 6736 38490 6788 38496
rect 6552 38276 6604 38282
rect 6552 38218 6604 38224
rect 6748 38010 6776 38490
rect 7116 38282 7144 38694
rect 7852 38350 7880 39782
rect 7840 38344 7892 38350
rect 7840 38286 7892 38292
rect 7104 38276 7156 38282
rect 7104 38218 7156 38224
rect 7472 38276 7524 38282
rect 7472 38218 7524 38224
rect 6828 38208 6880 38214
rect 6828 38150 6880 38156
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6840 37942 6868 38150
rect 6828 37936 6880 37942
rect 6828 37878 6880 37884
rect 7484 37806 7512 38218
rect 8036 37942 8064 40394
rect 8128 40186 8156 41006
rect 8668 40928 8720 40934
rect 8668 40870 8720 40876
rect 8576 40520 8628 40526
rect 8576 40462 8628 40468
rect 8116 40180 8168 40186
rect 8116 40122 8168 40128
rect 8588 39098 8616 40462
rect 8576 39092 8628 39098
rect 8576 39034 8628 39040
rect 8680 39030 8708 40870
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 8852 40384 8904 40390
rect 8852 40326 8904 40332
rect 8864 40050 8892 40326
rect 8852 40044 8904 40050
rect 8852 39986 8904 39992
rect 8668 39024 8720 39030
rect 8668 38966 8720 38972
rect 8208 38752 8260 38758
rect 8208 38694 8260 38700
rect 8024 37936 8076 37942
rect 8024 37878 8076 37884
rect 8116 37936 8168 37942
rect 8116 37878 8168 37884
rect 6368 37800 6420 37806
rect 6368 37742 6420 37748
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 7012 37800 7064 37806
rect 7012 37742 7064 37748
rect 7472 37800 7524 37806
rect 7472 37742 7524 37748
rect 6276 37664 6328 37670
rect 6276 37606 6328 37612
rect 6460 37664 6512 37670
rect 6460 37606 6512 37612
rect 6472 37194 6500 37606
rect 6736 37324 6788 37330
rect 6736 37266 6788 37272
rect 6460 37188 6512 37194
rect 6460 37130 6512 37136
rect 6092 37120 6144 37126
rect 6092 37062 6144 37068
rect 6644 37120 6696 37126
rect 6644 37062 6696 37068
rect 6104 36582 6132 37062
rect 6656 36922 6684 37062
rect 6644 36916 6696 36922
rect 6644 36858 6696 36864
rect 6644 36712 6696 36718
rect 6748 36666 6776 37266
rect 6696 36660 6776 36666
rect 6644 36654 6776 36660
rect 6656 36638 6776 36654
rect 6932 36666 6960 37742
rect 7024 36786 7052 37742
rect 7484 37262 7512 37742
rect 7472 37256 7524 37262
rect 7472 37198 7524 37204
rect 7012 36780 7064 36786
rect 7012 36722 7064 36728
rect 8128 36718 8156 37878
rect 8220 36786 8248 38694
rect 8760 38208 8812 38214
rect 8760 38150 8812 38156
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8116 36712 8168 36718
rect 8036 36672 8116 36700
rect 6932 36638 7052 36666
rect 6092 36576 6144 36582
rect 6092 36518 6144 36524
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 5908 36100 5960 36106
rect 5908 36042 5960 36048
rect 6012 35834 6040 36110
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 5908 35624 5960 35630
rect 5960 35584 6040 35612
rect 5908 35566 5960 35572
rect 5906 34504 5962 34513
rect 5828 34462 5906 34490
rect 5906 34439 5962 34448
rect 6012 34406 6040 35584
rect 6104 35290 6132 36518
rect 6552 36032 6604 36038
rect 6552 35974 6604 35980
rect 6276 35556 6328 35562
rect 6276 35498 6328 35504
rect 6092 35284 6144 35290
rect 6092 35226 6144 35232
rect 6184 34468 6236 34474
rect 6184 34410 6236 34416
rect 6000 34400 6052 34406
rect 6000 34342 6052 34348
rect 6012 33522 6040 34342
rect 6196 34241 6224 34410
rect 6182 34232 6238 34241
rect 6182 34167 6238 34176
rect 6288 34066 6316 35498
rect 6460 35488 6512 35494
rect 6460 35430 6512 35436
rect 6472 34066 6500 35430
rect 6564 35018 6592 35974
rect 6552 35012 6604 35018
rect 6552 34954 6604 34960
rect 6552 34400 6604 34406
rect 6552 34342 6604 34348
rect 6276 34060 6328 34066
rect 6276 34002 6328 34008
rect 6460 34060 6512 34066
rect 6460 34002 6512 34008
rect 6000 33516 6052 33522
rect 6000 33458 6052 33464
rect 6276 33108 6328 33114
rect 6276 33050 6328 33056
rect 5908 32768 5960 32774
rect 5908 32710 5960 32716
rect 5920 32298 5948 32710
rect 6288 32298 6316 33050
rect 5908 32292 5960 32298
rect 5908 32234 5960 32240
rect 6276 32292 6328 32298
rect 6276 32234 6328 32240
rect 5920 31754 5948 32234
rect 5908 31748 5960 31754
rect 5908 31690 5960 31696
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5828 28694 5856 28902
rect 5816 28688 5868 28694
rect 5816 28630 5868 28636
rect 5816 28552 5868 28558
rect 5816 28494 5868 28500
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5644 25906 5672 26250
rect 5736 25906 5764 26930
rect 5828 26489 5856 28494
rect 5920 26994 5948 31690
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 6196 29850 6224 30194
rect 6184 29844 6236 29850
rect 6184 29786 6236 29792
rect 6092 28484 6144 28490
rect 6092 28426 6144 28432
rect 6104 28150 6132 28426
rect 6092 28144 6144 28150
rect 6092 28086 6144 28092
rect 6196 27946 6224 29786
rect 6184 27940 6236 27946
rect 6184 27882 6236 27888
rect 6184 27600 6236 27606
rect 6184 27542 6236 27548
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 6092 27328 6144 27334
rect 6092 27270 6144 27276
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 5920 26897 5948 26930
rect 5906 26888 5962 26897
rect 5906 26823 5962 26832
rect 5908 26512 5960 26518
rect 5814 26480 5870 26489
rect 5908 26454 5960 26460
rect 5814 26415 5870 26424
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5828 26042 5856 26182
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5644 25294 5672 25638
rect 5814 25392 5870 25401
rect 5814 25327 5870 25336
rect 5828 25294 5856 25327
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5092 24262 5212 24290
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 4816 22494 4936 22522
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4250 21992 4306 22001
rect 4250 21927 4306 21936
rect 4158 21856 4214 21865
rect 4158 21791 4214 21800
rect 4172 21554 4200 21791
rect 4264 21554 4292 21927
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4264 21457 4292 21490
rect 4250 21448 4306 21457
rect 4356 21418 4384 22034
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21690 4476 21898
rect 4526 21720 4582 21729
rect 4436 21684 4488 21690
rect 4526 21655 4582 21664
rect 4436 21626 4488 21632
rect 4448 21554 4476 21626
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4250 21383 4306 21392
rect 4344 21412 4396 21418
rect 4344 21354 4396 21360
rect 4448 21350 4476 21490
rect 4540 21418 4568 21655
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4158 20632 4214 20641
rect 4158 20567 4214 20576
rect 3700 20528 3752 20534
rect 3700 20470 3752 20476
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 20262 3648 20402
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3712 19854 3740 20470
rect 4172 20466 4200 20567
rect 4540 20505 4568 20878
rect 4526 20496 4582 20505
rect 4160 20460 4212 20466
rect 4526 20431 4582 20440
rect 4160 20402 4212 20408
rect 3792 20392 3844 20398
rect 3844 20352 3924 20380
rect 3792 20334 3844 20340
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3804 19514 3832 19994
rect 3332 19450 3384 19456
rect 3436 19468 3556 19496
rect 3792 19508 3844 19514
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18766 3372 19110
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3068 18142 3188 18170
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 16250 2912 17070
rect 3068 16590 3096 18142
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15162 2820 15846
rect 3068 15162 3096 16526
rect 3160 15570 3188 18022
rect 3252 17338 3280 18226
rect 3436 17678 3464 19468
rect 3792 19450 3844 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 18970 3556 19314
rect 3896 19310 3924 20352
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19825 4660 21490
rect 4724 21010 4752 22170
rect 4816 22030 4844 22494
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4908 21842 4936 22374
rect 5000 22137 5028 24142
rect 5092 23905 5120 24142
rect 5078 23896 5134 23905
rect 5078 23831 5134 23840
rect 5184 23730 5212 24262
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5276 23905 5304 24142
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5262 23896 5318 23905
rect 5262 23831 5318 23840
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5092 23610 5120 23666
rect 5092 23594 5304 23610
rect 5092 23588 5316 23594
rect 5092 23582 5264 23588
rect 5092 22642 5120 23582
rect 5264 23530 5316 23536
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5262 23488 5318 23497
rect 5184 22982 5212 23462
rect 5368 23474 5396 24074
rect 5318 23446 5396 23474
rect 5262 23423 5318 23432
rect 5460 23066 5488 24890
rect 5552 24818 5580 25094
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 5552 24177 5580 24618
rect 5538 24168 5594 24177
rect 5538 24103 5594 24112
rect 5552 23866 5580 24103
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5538 23624 5594 23633
rect 5538 23559 5594 23568
rect 5276 23038 5488 23066
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 5170 22536 5226 22545
rect 5170 22471 5226 22480
rect 5078 22400 5134 22409
rect 5078 22335 5134 22344
rect 4986 22128 5042 22137
rect 4986 22063 5042 22072
rect 5092 22030 5120 22335
rect 5080 22024 5132 22030
rect 4986 21992 5042 22001
rect 5080 21966 5132 21972
rect 4986 21927 4988 21936
rect 5040 21927 5042 21936
rect 4988 21898 5040 21904
rect 4816 21814 4936 21842
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4724 20777 4752 20810
rect 4710 20768 4766 20777
rect 4710 20703 4766 20712
rect 4816 19854 4844 21814
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4894 21312 4950 21321
rect 4894 21247 4950 21256
rect 4908 21049 4936 21247
rect 4894 21040 4950 21049
rect 4894 20975 4950 20984
rect 4908 20466 4936 20975
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4894 20224 4950 20233
rect 4894 20159 4950 20168
rect 4908 20058 4936 20159
rect 5000 20058 5028 21490
rect 5092 20806 5120 21966
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5184 20505 5212 22471
rect 5276 22098 5304 23038
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5368 22817 5396 22918
rect 5354 22808 5410 22817
rect 5410 22766 5488 22794
rect 5354 22743 5410 22752
rect 5354 22536 5410 22545
rect 5460 22506 5488 22766
rect 5552 22642 5580 23559
rect 5644 23526 5672 24006
rect 5736 23866 5764 25230
rect 5814 25120 5870 25129
rect 5814 25055 5870 25064
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5828 23730 5856 25055
rect 5920 24886 5948 26454
rect 6012 26246 6040 27270
rect 6104 27130 6132 27270
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6196 27010 6224 27542
rect 6288 27130 6316 32234
rect 6368 31816 6420 31822
rect 6368 31758 6420 31764
rect 6380 30054 6408 31758
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 6472 30870 6500 31282
rect 6460 30864 6512 30870
rect 6460 30806 6512 30812
rect 6460 30592 6512 30598
rect 6460 30534 6512 30540
rect 6472 30297 6500 30534
rect 6458 30288 6514 30297
rect 6458 30223 6514 30232
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6460 29776 6512 29782
rect 6460 29718 6512 29724
rect 6472 29510 6500 29718
rect 6460 29504 6512 29510
rect 6460 29446 6512 29452
rect 6564 28994 6592 34342
rect 6656 34066 6684 36638
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6644 34060 6696 34066
rect 6644 34002 6696 34008
rect 6644 33516 6696 33522
rect 6644 33458 6696 33464
rect 6656 33114 6684 33458
rect 6644 33108 6696 33114
rect 6644 33050 6696 33056
rect 6644 29232 6696 29238
rect 6644 29174 6696 29180
rect 6472 28966 6592 28994
rect 6366 28792 6422 28801
rect 6366 28727 6422 28736
rect 6380 28626 6408 28727
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 6366 28520 6422 28529
rect 6366 28455 6422 28464
rect 6380 27606 6408 28455
rect 6368 27600 6420 27606
rect 6368 27542 6420 27548
rect 6380 27441 6408 27542
rect 6366 27432 6422 27441
rect 6366 27367 6422 27376
rect 6276 27124 6328 27130
rect 6276 27066 6328 27072
rect 6104 26982 6224 27010
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 5998 25664 6054 25673
rect 5998 25599 6054 25608
rect 6012 25294 6040 25599
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 5908 24880 5960 24886
rect 5960 24840 6040 24868
rect 5908 24822 5960 24828
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 5920 24449 5948 24686
rect 5906 24440 5962 24449
rect 5906 24375 5962 24384
rect 5920 24206 5948 24375
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 6012 23730 6040 24840
rect 6104 24206 6132 26982
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6196 25498 6224 26726
rect 6288 26382 6316 27066
rect 6472 26994 6500 28966
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6460 26988 6512 26994
rect 6460 26930 6512 26936
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 6104 23610 6132 24142
rect 6196 23644 6224 25434
rect 6288 24818 6316 26318
rect 6380 25838 6408 26930
rect 6472 26790 6500 26930
rect 6460 26784 6512 26790
rect 6460 26726 6512 26732
rect 6460 26512 6512 26518
rect 6564 26500 6592 28562
rect 6656 28234 6684 29174
rect 6748 28626 6776 36518
rect 6920 36100 6972 36106
rect 6920 36042 6972 36048
rect 6828 35012 6880 35018
rect 6828 34954 6880 34960
rect 6840 34202 6868 34954
rect 6932 34610 6960 36042
rect 7024 35630 7052 36638
rect 7104 36644 7156 36650
rect 7104 36586 7156 36592
rect 7012 35624 7064 35630
rect 7012 35566 7064 35572
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 7024 34610 7052 35022
rect 6920 34604 6972 34610
rect 6920 34546 6972 34552
rect 7012 34604 7064 34610
rect 7012 34546 7064 34552
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 7024 33930 7052 34546
rect 7116 34406 7144 36586
rect 7656 36236 7708 36242
rect 7656 36178 7708 36184
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7288 36032 7340 36038
rect 7288 35974 7340 35980
rect 7300 35834 7328 35974
rect 7392 35834 7420 36110
rect 7484 35834 7512 36110
rect 7288 35828 7340 35834
rect 7288 35770 7340 35776
rect 7380 35828 7432 35834
rect 7380 35770 7432 35776
rect 7472 35828 7524 35834
rect 7472 35770 7524 35776
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 7104 34400 7156 34406
rect 7104 34342 7156 34348
rect 7208 33998 7236 35430
rect 7392 35290 7420 35770
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7668 35222 7696 36178
rect 7748 35760 7800 35766
rect 7748 35702 7800 35708
rect 7656 35216 7708 35222
rect 7656 35158 7708 35164
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7576 34202 7604 35022
rect 7760 34746 7788 35702
rect 8036 35630 8064 36672
rect 8116 36654 8168 36660
rect 8116 36168 8168 36174
rect 8312 36145 8340 37810
rect 8392 37460 8444 37466
rect 8392 37402 8444 37408
rect 8116 36110 8168 36116
rect 8298 36136 8354 36145
rect 8128 35834 8156 36110
rect 8298 36071 8354 36080
rect 8116 35828 8168 35834
rect 8116 35770 8168 35776
rect 8300 35760 8352 35766
rect 8404 35748 8432 37402
rect 8484 37324 8536 37330
rect 8484 37266 8536 37272
rect 8496 36378 8524 37266
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8484 36372 8536 36378
rect 8484 36314 8536 36320
rect 8352 35720 8432 35748
rect 8300 35702 8352 35708
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 8588 35154 8616 37198
rect 8668 37188 8720 37194
rect 8668 37130 8720 37136
rect 8680 35290 8708 37130
rect 8772 36582 8800 38150
rect 8956 37806 8984 40462
rect 9140 39642 9168 41006
rect 9680 40928 9732 40934
rect 9680 40870 9732 40876
rect 9588 40112 9640 40118
rect 9588 40054 9640 40060
rect 9496 40044 9548 40050
rect 9496 39986 9548 39992
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 9312 39976 9364 39982
rect 9312 39918 9364 39924
rect 9404 39976 9456 39982
rect 9404 39918 9456 39924
rect 9128 39636 9180 39642
rect 9128 39578 9180 39584
rect 9232 38894 9260 39918
rect 9220 38888 9272 38894
rect 9220 38830 9272 38836
rect 9232 38486 9260 38830
rect 9220 38480 9272 38486
rect 9220 38422 9272 38428
rect 9036 38344 9088 38350
rect 9036 38286 9088 38292
rect 8944 37800 8996 37806
rect 8944 37742 8996 37748
rect 9048 37466 9076 38286
rect 9036 37460 9088 37466
rect 9036 37402 9088 37408
rect 8944 37120 8996 37126
rect 8944 37062 8996 37068
rect 8760 36576 8812 36582
rect 8760 36518 8812 36524
rect 8760 36032 8812 36038
rect 8760 35974 8812 35980
rect 8772 35834 8800 35974
rect 8760 35828 8812 35834
rect 8760 35770 8812 35776
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8576 35148 8628 35154
rect 8576 35090 8628 35096
rect 8208 34944 8260 34950
rect 8208 34886 8260 34892
rect 7748 34740 7800 34746
rect 7748 34682 7800 34688
rect 7564 34196 7616 34202
rect 7564 34138 7616 34144
rect 7196 33992 7248 33998
rect 7196 33934 7248 33940
rect 7472 33992 7524 33998
rect 7472 33934 7524 33940
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 7024 32910 7052 33866
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 7024 32230 7052 32846
rect 7012 32224 7064 32230
rect 7012 32166 7064 32172
rect 7024 31890 7052 32166
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6840 31482 6868 31758
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 6932 30938 6960 31350
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7116 30938 7144 31282
rect 6920 30932 6972 30938
rect 6920 30874 6972 30880
rect 7104 30932 7156 30938
rect 7104 30874 7156 30880
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 6932 30394 6960 30534
rect 6920 30388 6972 30394
rect 6920 30330 6972 30336
rect 7116 30326 7144 30534
rect 7300 30374 7328 33798
rect 7380 33448 7432 33454
rect 7380 33390 7432 33396
rect 7392 32570 7420 33390
rect 7484 32774 7512 33934
rect 7932 33312 7984 33318
rect 7932 33254 7984 33260
rect 7944 32910 7972 33254
rect 7932 32904 7984 32910
rect 7932 32846 7984 32852
rect 7472 32768 7524 32774
rect 7472 32710 7524 32716
rect 7380 32564 7432 32570
rect 7380 32506 7432 32512
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7392 32026 7420 32370
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7472 31680 7524 31686
rect 7472 31622 7524 31628
rect 7484 31278 7512 31622
rect 7576 31414 7604 31758
rect 7564 31408 7616 31414
rect 7564 31350 7616 31356
rect 7748 31408 7800 31414
rect 7748 31350 7800 31356
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 7300 30346 7420 30374
rect 7104 30320 7156 30326
rect 7104 30262 7156 30268
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 6840 29850 6868 30194
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6828 29640 6880 29646
rect 7196 29640 7248 29646
rect 6880 29588 6960 29594
rect 6828 29582 6960 29588
rect 7196 29582 7248 29588
rect 6840 29566 6960 29582
rect 6736 28620 6788 28626
rect 6736 28562 6788 28568
rect 6736 28484 6788 28490
rect 6932 28472 6960 29566
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 7024 29306 7052 29514
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 7024 28966 7052 29106
rect 7012 28960 7064 28966
rect 7012 28902 7064 28908
rect 7208 28762 7236 29582
rect 7286 29472 7342 29481
rect 7286 29407 7342 29416
rect 7300 29170 7328 29407
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7196 28484 7248 28490
rect 6932 28444 7196 28472
rect 6736 28426 6788 28432
rect 7248 28444 7328 28472
rect 7196 28426 7248 28432
rect 6647 28206 6684 28234
rect 6748 28218 6776 28426
rect 6736 28212 6788 28218
rect 6647 28082 6675 28206
rect 6736 28154 6788 28160
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6642 27976 6698 27985
rect 6642 27911 6698 27920
rect 6512 26472 6592 26500
rect 6460 26454 6512 26460
rect 6458 26072 6514 26081
rect 6458 26007 6514 26016
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6366 25664 6422 25673
rect 6366 25599 6422 25608
rect 6380 24970 6408 25599
rect 6472 25294 6500 26007
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6564 25673 6592 25842
rect 6656 25702 6684 27911
rect 6748 27520 6776 28018
rect 6840 27878 6868 28018
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 7010 27840 7066 27849
rect 7010 27775 7066 27784
rect 6748 27492 6868 27520
rect 6734 27432 6790 27441
rect 6734 27367 6790 27376
rect 6748 26994 6776 27367
rect 6840 27334 6868 27492
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6840 26382 6868 26930
rect 7024 26790 7052 27775
rect 7116 27674 7144 28086
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 7208 27334 7236 28018
rect 7300 27470 7328 28444
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7194 27160 7250 27169
rect 7194 27095 7250 27104
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 6828 26376 6880 26382
rect 6734 26344 6790 26353
rect 6828 26318 6880 26324
rect 6734 26279 6790 26288
rect 6748 26042 6776 26279
rect 7104 26240 7156 26246
rect 7104 26182 7156 26188
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 7116 25906 7144 26182
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 6644 25696 6696 25702
rect 6550 25664 6606 25673
rect 6644 25638 6696 25644
rect 6550 25599 6606 25608
rect 6564 25294 6592 25599
rect 6656 25401 6684 25638
rect 6748 25486 6960 25514
rect 6642 25392 6698 25401
rect 6642 25327 6698 25336
rect 6748 25294 6776 25486
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6460 25152 6512 25158
rect 6458 25120 6460 25129
rect 6736 25152 6788 25158
rect 6512 25120 6514 25129
rect 6736 25094 6788 25100
rect 6458 25055 6514 25064
rect 6550 24984 6606 24993
rect 6380 24942 6500 24970
rect 6276 24812 6328 24818
rect 6472 24800 6500 24942
rect 6606 24942 6684 24970
rect 6748 24954 6776 25094
rect 6550 24919 6606 24928
rect 6656 24818 6684 24942
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6552 24812 6604 24818
rect 6328 24772 6408 24800
rect 6472 24772 6552 24800
rect 6276 24754 6328 24760
rect 6274 24712 6330 24721
rect 6274 24647 6330 24656
rect 6380 24664 6408 24772
rect 6552 24754 6604 24760
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6288 24614 6316 24647
rect 6380 24636 6500 24664
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6366 24576 6422 24585
rect 6366 24511 6422 24520
rect 6380 24206 6408 24511
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6472 23712 6500 24636
rect 6564 24188 6592 24754
rect 6644 24200 6696 24206
rect 6564 24160 6644 24188
rect 6644 24142 6696 24148
rect 6748 23730 6776 24754
rect 6840 24342 6868 25298
rect 6932 25208 6960 25486
rect 6932 25180 6965 25208
rect 6937 24970 6965 25180
rect 7024 24993 7052 25842
rect 7208 25430 7236 27095
rect 7300 26926 7328 27406
rect 7288 26920 7340 26926
rect 7288 26862 7340 26868
rect 7392 26382 7420 30346
rect 7484 27962 7512 31214
rect 7656 31136 7708 31142
rect 7656 31078 7708 31084
rect 7668 30870 7696 31078
rect 7656 30864 7708 30870
rect 7656 30806 7708 30812
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 7576 30190 7604 30670
rect 7564 30184 7616 30190
rect 7564 30126 7616 30132
rect 7668 30054 7696 30806
rect 7760 30734 7788 31350
rect 7748 30728 7800 30734
rect 7748 30670 7800 30676
rect 7760 30258 7788 30670
rect 7852 30598 7880 32302
rect 8220 32298 8248 34886
rect 8668 34536 8720 34542
rect 8668 34478 8720 34484
rect 8574 34232 8630 34241
rect 8574 34167 8576 34176
rect 8628 34167 8630 34176
rect 8576 34138 8628 34144
rect 8680 34066 8708 34478
rect 8668 34060 8720 34066
rect 8668 34002 8720 34008
rect 8680 33658 8708 34002
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 8772 33658 8800 33934
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 8864 33402 8892 35634
rect 8956 35154 8984 37062
rect 9036 36576 9088 36582
rect 9036 36518 9088 36524
rect 9048 36310 9076 36518
rect 9036 36304 9088 36310
rect 9036 36246 9088 36252
rect 9048 36174 9076 36246
rect 9036 36168 9088 36174
rect 9036 36110 9088 36116
rect 9048 35698 9076 36110
rect 9036 35692 9088 35698
rect 9036 35634 9088 35640
rect 9048 35222 9076 35634
rect 9232 35612 9260 38422
rect 9324 38010 9352 39918
rect 9416 39302 9444 39918
rect 9404 39296 9456 39302
rect 9404 39238 9456 39244
rect 9312 38004 9364 38010
rect 9312 37946 9364 37952
rect 9416 37806 9444 39238
rect 9508 39030 9536 39986
rect 9496 39024 9548 39030
rect 9496 38966 9548 38972
rect 9496 38888 9548 38894
rect 9496 38830 9548 38836
rect 9404 37800 9456 37806
rect 9404 37742 9456 37748
rect 9416 37126 9444 37742
rect 9404 37120 9456 37126
rect 9404 37062 9456 37068
rect 9312 36168 9364 36174
rect 9310 36136 9312 36145
rect 9364 36136 9366 36145
rect 9310 36071 9366 36080
rect 9416 35834 9444 37062
rect 9508 36718 9536 38830
rect 9600 38010 9628 40054
rect 9692 39438 9720 40870
rect 10060 40186 10088 41006
rect 10600 40928 10652 40934
rect 10600 40870 10652 40876
rect 10416 40520 10468 40526
rect 10416 40462 10468 40468
rect 10048 40180 10100 40186
rect 10048 40122 10100 40128
rect 9772 39840 9824 39846
rect 9772 39782 9824 39788
rect 9784 39574 9812 39782
rect 9772 39568 9824 39574
rect 9772 39510 9824 39516
rect 9680 39432 9732 39438
rect 9680 39374 9732 39380
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9692 39098 9720 39374
rect 9680 39092 9732 39098
rect 9680 39034 9732 39040
rect 9784 38894 9812 39374
rect 9772 38888 9824 38894
rect 9772 38830 9824 38836
rect 9680 38208 9732 38214
rect 9680 38150 9732 38156
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 9600 36786 9628 37946
rect 9692 37194 9720 38150
rect 9784 37262 9812 38830
rect 10428 38554 10456 40462
rect 10612 39438 10640 40870
rect 10876 40452 10928 40458
rect 10876 40394 10928 40400
rect 10784 39976 10836 39982
rect 10784 39918 10836 39924
rect 10600 39432 10652 39438
rect 10600 39374 10652 39380
rect 10232 38548 10284 38554
rect 10232 38490 10284 38496
rect 10416 38548 10468 38554
rect 10416 38490 10468 38496
rect 9864 37664 9916 37670
rect 9864 37606 9916 37612
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9680 37188 9732 37194
rect 9680 37130 9732 37136
rect 9692 36922 9720 37130
rect 9680 36916 9732 36922
rect 9680 36858 9732 36864
rect 9784 36786 9812 37198
rect 9588 36780 9640 36786
rect 9588 36722 9640 36728
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9496 36712 9548 36718
rect 9876 36666 9904 37606
rect 9496 36654 9548 36660
rect 9508 36038 9536 36654
rect 9692 36638 9904 36666
rect 9496 36032 9548 36038
rect 9496 35974 9548 35980
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9692 35737 9720 36638
rect 9772 36304 9824 36310
rect 9772 36246 9824 36252
rect 9678 35728 9734 35737
rect 9784 35698 9812 36246
rect 10140 36100 10192 36106
rect 10140 36042 10192 36048
rect 10152 35766 10180 36042
rect 10140 35760 10192 35766
rect 10140 35702 10192 35708
rect 9678 35663 9680 35672
rect 9732 35663 9734 35672
rect 9772 35692 9824 35698
rect 9680 35634 9732 35640
rect 9772 35634 9824 35640
rect 9404 35624 9456 35630
rect 9232 35584 9404 35612
rect 9404 35566 9456 35572
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9036 35216 9088 35222
rect 9036 35158 9088 35164
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 9220 35080 9272 35086
rect 9220 35022 9272 35028
rect 9232 34542 9260 35022
rect 9600 34678 9628 35430
rect 9692 35193 9720 35634
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9956 35488 10008 35494
rect 9956 35430 10008 35436
rect 9876 35290 9904 35430
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9678 35184 9734 35193
rect 9678 35119 9734 35128
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9588 34672 9640 34678
rect 9588 34614 9640 34620
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 9232 34218 9260 34478
rect 9232 34202 9352 34218
rect 9128 34196 9180 34202
rect 9232 34196 9364 34202
rect 9232 34190 9312 34196
rect 9128 34138 9180 34144
rect 9312 34138 9364 34144
rect 9140 33640 9168 34138
rect 9140 33612 9352 33640
rect 9324 33522 9352 33612
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 9220 33516 9272 33522
rect 9220 33458 9272 33464
rect 9312 33516 9364 33522
rect 9312 33458 9364 33464
rect 8772 33374 8892 33402
rect 8392 33312 8444 33318
rect 8392 33254 8444 33260
rect 8404 32910 8432 33254
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 8312 32570 8340 32710
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8208 32292 8260 32298
rect 8208 32234 8260 32240
rect 8220 31906 8248 32234
rect 7944 31878 8248 31906
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7852 30394 7880 30534
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7748 30252 7800 30258
rect 7748 30194 7800 30200
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7840 29640 7892 29646
rect 7838 29608 7840 29617
rect 7892 29608 7894 29617
rect 7838 29543 7894 29552
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7576 28422 7604 29106
rect 7852 28762 7880 29242
rect 7944 28994 7972 31878
rect 8220 31822 8248 31878
rect 8024 31816 8076 31822
rect 8208 31816 8260 31822
rect 8076 31764 8156 31770
rect 8024 31758 8156 31764
rect 8208 31758 8260 31764
rect 8036 31742 8156 31758
rect 8128 31498 8156 31742
rect 8128 31470 8248 31498
rect 8116 31408 8168 31414
rect 8116 31350 8168 31356
rect 8128 30394 8156 31350
rect 8220 31346 8248 31470
rect 8404 31362 8432 32846
rect 8680 32502 8708 32914
rect 8668 32496 8720 32502
rect 8668 32438 8720 32444
rect 8576 32360 8628 32366
rect 8576 32302 8628 32308
rect 8588 32026 8616 32302
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8484 31748 8536 31754
rect 8484 31690 8536 31696
rect 8496 31482 8524 31690
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8208 31340 8260 31346
rect 8404 31334 8524 31362
rect 8208 31282 8260 31288
rect 8220 30870 8248 31282
rect 8208 30864 8260 30870
rect 8208 30806 8260 30812
rect 8116 30388 8168 30394
rect 8116 30330 8168 30336
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8128 29646 8156 30126
rect 8220 29850 8248 30126
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8128 29306 8156 29582
rect 8116 29300 8168 29306
rect 8116 29242 8168 29248
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 7944 28966 8156 28994
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7564 28416 7616 28422
rect 7564 28358 7616 28364
rect 8024 28008 8076 28014
rect 7484 27934 7880 27962
rect 8024 27950 8076 27956
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7576 27470 7604 27814
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7484 26790 7512 27406
rect 7748 27328 7800 27334
rect 7746 27296 7748 27305
rect 7800 27296 7802 27305
rect 7746 27231 7802 27240
rect 7656 27056 7708 27062
rect 7654 27024 7656 27033
rect 7708 27024 7710 27033
rect 7564 26988 7616 26994
rect 7760 26994 7788 27231
rect 7654 26959 7710 26968
rect 7748 26988 7800 26994
rect 7564 26930 7616 26936
rect 7748 26930 7800 26936
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7576 26518 7604 26930
rect 7760 26586 7788 26930
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7380 26376 7432 26382
rect 7380 26318 7432 26324
rect 7300 25702 7328 26318
rect 7288 25696 7340 25702
rect 7392 25673 7420 26318
rect 7576 26314 7604 26454
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7748 26240 7800 26246
rect 7470 26208 7526 26217
rect 7748 26182 7800 26188
rect 7470 26143 7526 26152
rect 7288 25638 7340 25644
rect 7378 25664 7434 25673
rect 7378 25599 7434 25608
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 6932 24942 6965 24970
rect 7010 24984 7066 24993
rect 6932 24886 6960 24942
rect 7010 24919 7066 24928
rect 6920 24880 6972 24886
rect 6920 24822 6972 24828
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6932 24410 6960 24550
rect 7024 24410 7052 24754
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 6828 24336 6880 24342
rect 6828 24278 6880 24284
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6840 23866 6868 24074
rect 6932 24041 6960 24074
rect 6918 24032 6974 24041
rect 6918 23967 6974 23976
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6736 23724 6788 23730
rect 6472 23684 6684 23712
rect 6196 23616 6500 23644
rect 6012 23582 6132 23610
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5828 23225 5856 23462
rect 6012 23361 6040 23582
rect 5998 23352 6054 23361
rect 5998 23287 6054 23296
rect 6368 23248 6420 23254
rect 5814 23216 5870 23225
rect 6368 23190 6420 23196
rect 5814 23151 5870 23160
rect 5908 23180 5960 23186
rect 5828 23118 5856 23151
rect 5960 23140 6096 23168
rect 5908 23122 5960 23128
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 6068 23066 6096 23140
rect 6380 23089 6408 23190
rect 6366 23080 6422 23089
rect 5632 23044 5684 23050
rect 6068 23038 6132 23066
rect 5684 23004 5764 23032
rect 5632 22986 5684 22992
rect 5736 22964 5764 23004
rect 5736 22936 5856 22964
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5354 22471 5410 22480
rect 5448 22500 5500 22506
rect 5368 22234 5396 22471
rect 5448 22442 5500 22448
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5354 22128 5410 22137
rect 5264 22092 5316 22098
rect 5354 22063 5410 22072
rect 5264 22034 5316 22040
rect 5368 22030 5396 22063
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 5264 21956 5316 21962
rect 5264 21898 5316 21904
rect 5276 21622 5304 21898
rect 5448 21888 5500 21894
rect 5354 21856 5410 21865
rect 5448 21830 5500 21836
rect 5354 21791 5410 21800
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 5368 21554 5396 21791
rect 5460 21690 5488 21830
rect 5552 21729 5580 22578
rect 5644 22234 5672 22578
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5736 22098 5764 22578
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5828 21894 5856 22936
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 5920 22409 5948 22578
rect 6104 22545 6132 23038
rect 6366 23015 6422 23024
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6090 22536 6146 22545
rect 6000 22500 6052 22506
rect 6090 22471 6146 22480
rect 6000 22442 6052 22448
rect 5906 22400 5962 22409
rect 5906 22335 5962 22344
rect 5908 22160 5960 22166
rect 5906 22128 5908 22137
rect 5960 22128 5962 22137
rect 5906 22063 5962 22072
rect 6012 22030 6040 22442
rect 6092 22432 6144 22438
rect 6288 22409 6316 22578
rect 6092 22374 6144 22380
rect 6274 22400 6330 22409
rect 6104 22030 6132 22374
rect 6274 22335 6330 22344
rect 6288 22098 6316 22335
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5538 21720 5594 21729
rect 5448 21684 5500 21690
rect 5538 21655 5594 21664
rect 5632 21684 5684 21690
rect 5448 21626 5500 21632
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5262 21176 5318 21185
rect 5262 21111 5318 21120
rect 5276 20602 5304 21111
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 5368 20602 5396 20946
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5170 20496 5226 20505
rect 5170 20431 5226 20440
rect 5276 20448 5304 20538
rect 5276 20420 5396 20448
rect 5172 20256 5224 20262
rect 5224 20216 5304 20244
rect 5172 20198 5224 20204
rect 5276 20097 5304 20216
rect 5262 20088 5318 20097
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4988 20052 5040 20058
rect 5262 20023 5318 20032
rect 4988 19994 5040 20000
rect 4986 19952 5042 19961
rect 5262 19952 5318 19961
rect 4986 19887 5042 19896
rect 5092 19910 5262 19938
rect 5000 19854 5028 19887
rect 5092 19854 5120 19910
rect 5262 19887 5318 19896
rect 4804 19848 4856 19854
rect 4250 19816 4306 19825
rect 3976 19780 4028 19786
rect 4250 19751 4306 19760
rect 4618 19816 4674 19825
rect 4804 19790 4856 19796
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5080 19848 5132 19854
rect 5264 19848 5316 19854
rect 5080 19790 5132 19796
rect 5262 19816 5264 19825
rect 5316 19816 5318 19825
rect 4618 19751 4674 19760
rect 5262 19751 5318 19760
rect 3976 19722 4028 19728
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3514 18864 3570 18873
rect 3514 18799 3570 18808
rect 3528 18426 3556 18799
rect 3606 18456 3662 18465
rect 3516 18420 3568 18426
rect 3606 18391 3608 18400
rect 3516 18362 3568 18368
rect 3660 18391 3662 18400
rect 3608 18362 3660 18368
rect 3528 17882 3556 18362
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3620 17746 3648 18362
rect 3896 18222 3924 19246
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3252 15026 3280 16934
rect 3344 16794 3372 17138
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3436 15706 3464 17138
rect 3608 16652 3660 16658
rect 3712 16640 3740 18158
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17678 3924 18022
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3804 16658 3832 17138
rect 3660 16612 3740 16640
rect 3608 16594 3660 16600
rect 3712 16046 3740 16612
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3528 14958 3556 15846
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3712 14822 3740 15982
rect 3804 15434 3832 16594
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3896 15706 3924 15982
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3252 14618 3280 14758
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 3252 14006 3280 14554
rect 3804 14482 3832 15370
rect 3988 15162 4016 19722
rect 4066 19680 4122 19689
rect 4066 19615 4122 19624
rect 4080 19378 4108 19615
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 18970 4108 19314
rect 4264 19242 4292 19751
rect 5264 19712 5316 19718
rect 4908 19672 5264 19700
rect 4526 19544 4582 19553
rect 4526 19479 4582 19488
rect 4540 19378 4568 19479
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4804 19372 4856 19378
rect 4908 19360 4936 19672
rect 5264 19654 5316 19660
rect 5170 19544 5226 19553
rect 5170 19479 5226 19488
rect 4856 19332 4936 19360
rect 4986 19408 5042 19417
rect 4986 19343 4988 19352
rect 4804 19314 4856 19320
rect 5040 19343 5042 19352
rect 4988 19314 5040 19320
rect 5184 19310 5212 19479
rect 5368 19446 5396 20420
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5460 19378 5488 21626
rect 5552 21078 5580 21655
rect 5632 21626 5684 21632
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5644 21593 5672 21626
rect 5630 21584 5686 21593
rect 5630 21519 5686 21528
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5632 21072 5684 21078
rect 5632 21014 5684 21020
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5552 20466 5580 20810
rect 5644 20534 5672 21014
rect 5632 20528 5684 20534
rect 5632 20470 5684 20476
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4908 18426 4936 18634
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 18426 5120 18566
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18158
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 4620 17740 4672 17746
rect 4080 16998 4108 17711
rect 4724 17728 4752 18022
rect 4816 17746 4844 18294
rect 4672 17700 4752 17728
rect 4804 17740 4856 17746
rect 4620 17682 4672 17688
rect 4804 17682 4856 17688
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 16998 4476 17614
rect 4816 17338 4844 17682
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4908 16794 4936 17138
rect 5184 17082 5212 18906
rect 5276 18834 5304 19246
rect 5552 19174 5580 20402
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5644 18766 5672 19994
rect 5736 19514 5764 21626
rect 5828 21554 5856 21830
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6012 21298 6040 21626
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 5828 21270 6040 21298
rect 5828 21185 5856 21270
rect 5814 21176 5870 21185
rect 5814 21111 5870 21120
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5828 20602 5856 20878
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5828 19378 5856 20266
rect 5920 19961 5948 20742
rect 6012 20058 6040 21082
rect 6104 20330 6132 21422
rect 6196 20777 6224 21830
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6288 21321 6316 21558
rect 6380 21418 6408 22918
rect 6472 22098 6500 23616
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6564 22778 6592 22918
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6564 22545 6592 22714
rect 6656 22710 6684 23684
rect 6736 23666 6788 23672
rect 6734 23624 6790 23633
rect 6734 23559 6790 23568
rect 6748 23254 6776 23559
rect 6840 23526 6868 23802
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6736 23248 6788 23254
rect 6736 23190 6788 23196
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6656 22574 6684 22646
rect 6644 22568 6696 22574
rect 6550 22536 6606 22545
rect 6644 22510 6696 22516
rect 6550 22471 6606 22480
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6550 21856 6606 21865
rect 6550 21791 6606 21800
rect 6564 21457 6592 21791
rect 6550 21448 6606 21457
rect 6368 21412 6420 21418
rect 6550 21383 6606 21392
rect 6368 21354 6420 21360
rect 6274 21312 6330 21321
rect 6274 21247 6330 21256
rect 6366 21176 6422 21185
rect 6288 21134 6366 21162
rect 6288 21078 6316 21134
rect 6366 21111 6422 21120
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6182 20768 6238 20777
rect 6564 20754 6592 21383
rect 6182 20703 6238 20712
rect 6472 20726 6592 20754
rect 6472 20602 6500 20726
rect 6550 20632 6606 20641
rect 6460 20596 6512 20602
rect 6550 20567 6606 20576
rect 6460 20538 6512 20544
rect 6276 20460 6328 20466
rect 6328 20420 6500 20448
rect 6276 20402 6328 20408
rect 6184 20392 6236 20398
rect 6236 20340 6316 20346
rect 6184 20334 6316 20340
rect 6092 20324 6144 20330
rect 6196 20318 6316 20334
rect 6092 20266 6144 20272
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6196 19961 6224 20198
rect 5906 19952 5962 19961
rect 5906 19887 5962 19896
rect 6182 19952 6238 19961
rect 6182 19887 6238 19896
rect 6288 19514 6316 20318
rect 6472 20058 6500 20420
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6564 19854 6592 20567
rect 6368 19848 6420 19854
rect 6366 19816 6368 19825
rect 6552 19848 6604 19854
rect 6420 19816 6422 19825
rect 6552 19790 6604 19796
rect 6366 19751 6422 19760
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5460 17270 5488 18158
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5552 17270 5580 17818
rect 5644 17746 5672 18362
rect 5828 18290 5856 19110
rect 5920 18970 5948 19314
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6012 18698 6040 19314
rect 6090 19136 6146 19145
rect 6090 19071 6146 19080
rect 6104 18902 6132 19071
rect 6196 18902 6224 19314
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6380 18834 6408 19751
rect 6656 19446 6684 22510
rect 6748 22438 6776 23054
rect 6840 22642 6868 23462
rect 6932 23089 6960 23967
rect 7024 23798 7052 24142
rect 7116 24070 7144 25230
rect 7194 25120 7250 25129
rect 7194 25055 7250 25064
rect 7208 24818 7236 25055
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7102 23896 7158 23905
rect 7102 23831 7158 23840
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7024 23361 7052 23462
rect 7010 23352 7066 23361
rect 7116 23322 7144 23831
rect 7208 23322 7236 24754
rect 7392 24138 7420 25366
rect 7484 25158 7512 26143
rect 7562 26072 7618 26081
rect 7562 26007 7618 26016
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7576 24936 7604 26007
rect 7760 25702 7788 26182
rect 7748 25696 7800 25702
rect 7748 25638 7800 25644
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7484 24908 7604 24936
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7010 23287 7066 23296
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7104 23112 7156 23118
rect 6918 23080 6974 23089
rect 7104 23054 7156 23060
rect 6918 23015 6974 23024
rect 6920 22976 6972 22982
rect 6918 22944 6920 22953
rect 6972 22944 6974 22953
rect 6918 22879 6974 22888
rect 7116 22642 7144 23054
rect 7196 22704 7248 22710
rect 7300 22692 7328 23598
rect 7392 23361 7420 24074
rect 7484 24052 7512 24908
rect 7668 24886 7696 25094
rect 7760 24970 7788 25638
rect 7852 25106 7880 27934
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7944 27470 7972 27814
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 8036 26926 8064 27950
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 7932 25968 7984 25974
rect 7932 25910 7984 25916
rect 7944 25226 7972 25910
rect 8036 25838 8064 26862
rect 8128 26314 8156 28966
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8312 28626 8340 28902
rect 8300 28620 8352 28626
rect 8300 28562 8352 28568
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 8208 27940 8260 27946
rect 8208 27882 8260 27888
rect 8220 27606 8248 27882
rect 8312 27713 8340 28018
rect 8298 27704 8354 27713
rect 8298 27639 8300 27648
rect 8352 27639 8354 27648
rect 8300 27610 8352 27616
rect 8404 27606 8432 29174
rect 8208 27600 8260 27606
rect 8208 27542 8260 27548
rect 8392 27600 8444 27606
rect 8392 27542 8444 27548
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8298 27432 8354 27441
rect 8220 27305 8248 27406
rect 8496 27418 8524 31334
rect 8680 31210 8708 32438
rect 8772 32212 8800 33374
rect 8852 32904 8904 32910
rect 8852 32846 8904 32852
rect 8864 32774 8892 32846
rect 8852 32768 8904 32774
rect 8852 32710 8904 32716
rect 9140 32298 9168 33458
rect 9232 33114 9260 33458
rect 9220 33108 9272 33114
rect 9220 33050 9272 33056
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9232 32502 9260 32846
rect 9324 32570 9352 33458
rect 9416 33114 9444 34614
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9600 33930 9628 34478
rect 9784 34202 9812 35090
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 9876 34610 9904 34886
rect 9968 34746 9996 35430
rect 10152 34746 10180 35702
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 10140 34740 10192 34746
rect 10140 34682 10192 34688
rect 10152 34610 10180 34682
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 9968 34202 9996 34546
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9588 33924 9640 33930
rect 9588 33866 9640 33872
rect 9600 33658 9628 33866
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9770 33144 9826 33153
rect 9404 33108 9456 33114
rect 9770 33079 9826 33088
rect 9404 33050 9456 33056
rect 9784 32910 9812 33079
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9220 32496 9272 32502
rect 9220 32438 9272 32444
rect 10244 32366 10272 38490
rect 10796 38418 10824 39918
rect 10784 38412 10836 38418
rect 10784 38354 10836 38360
rect 10416 38208 10468 38214
rect 10416 38150 10468 38156
rect 10428 38010 10456 38150
rect 10416 38004 10468 38010
rect 10416 37946 10468 37952
rect 10796 37874 10824 38354
rect 10888 38350 10916 40394
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 10980 39030 11008 40326
rect 11164 39642 11192 41006
rect 11336 40928 11388 40934
rect 11336 40870 11388 40876
rect 11244 40520 11296 40526
rect 11244 40462 11296 40468
rect 11152 39636 11204 39642
rect 11152 39578 11204 39584
rect 10968 39024 11020 39030
rect 10968 38966 11020 38972
rect 11060 38752 11112 38758
rect 11060 38694 11112 38700
rect 11072 38554 11100 38694
rect 11060 38548 11112 38554
rect 11060 38490 11112 38496
rect 10876 38344 10928 38350
rect 10876 38286 10928 38292
rect 11060 38276 11112 38282
rect 11060 38218 11112 38224
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 10968 37800 11020 37806
rect 10968 37742 11020 37748
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10428 36242 10456 37606
rect 10980 37312 11008 37742
rect 11072 37466 11100 38218
rect 11164 37806 11192 39578
rect 11256 39098 11284 40462
rect 11348 40186 11376 40870
rect 12268 40730 12296 41006
rect 12808 40928 12860 40934
rect 12808 40870 12860 40876
rect 12992 40928 13044 40934
rect 12992 40870 13044 40876
rect 12256 40724 12308 40730
rect 12256 40666 12308 40672
rect 11888 40520 11940 40526
rect 11888 40462 11940 40468
rect 11336 40180 11388 40186
rect 11336 40122 11388 40128
rect 11520 39432 11572 39438
rect 11520 39374 11572 39380
rect 11336 39296 11388 39302
rect 11336 39238 11388 39244
rect 11244 39092 11296 39098
rect 11244 39034 11296 39040
rect 11256 38010 11284 39034
rect 11244 38004 11296 38010
rect 11244 37946 11296 37952
rect 11152 37800 11204 37806
rect 11152 37742 11204 37748
rect 11348 37466 11376 39238
rect 11532 39098 11560 39374
rect 11900 39098 11928 40462
rect 12440 40384 12492 40390
rect 12440 40326 12492 40332
rect 11980 39976 12032 39982
rect 11980 39918 12032 39924
rect 11992 39438 12020 39918
rect 12452 39438 12480 40326
rect 12820 40118 12848 40870
rect 12808 40112 12860 40118
rect 12808 40054 12860 40060
rect 11980 39432 12032 39438
rect 11980 39374 12032 39380
rect 12440 39432 12492 39438
rect 12440 39374 12492 39380
rect 11520 39092 11572 39098
rect 11520 39034 11572 39040
rect 11888 39092 11940 39098
rect 11888 39034 11940 39040
rect 11992 38418 12020 39374
rect 12532 39296 12584 39302
rect 12532 39238 12584 39244
rect 12348 38888 12400 38894
rect 12348 38830 12400 38836
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 12256 38412 12308 38418
rect 12256 38354 12308 38360
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 11428 37664 11480 37670
rect 11428 37606 11480 37612
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 11336 37460 11388 37466
rect 11336 37402 11388 37408
rect 11440 37398 11468 37606
rect 11428 37392 11480 37398
rect 11428 37334 11480 37340
rect 10980 37284 11100 37312
rect 11072 37194 11100 37284
rect 10968 37188 11020 37194
rect 10968 37130 11020 37136
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 10980 36378 11008 37130
rect 11336 37120 11388 37126
rect 11336 37062 11388 37068
rect 11348 36922 11376 37062
rect 11336 36916 11388 36922
rect 11336 36858 11388 36864
rect 11532 36854 11560 37606
rect 11808 37262 11836 37810
rect 11796 37256 11848 37262
rect 11796 37198 11848 37204
rect 11520 36848 11572 36854
rect 11520 36790 11572 36796
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 11072 36378 11100 36722
rect 11520 36576 11572 36582
rect 11520 36518 11572 36524
rect 10968 36372 11020 36378
rect 10968 36314 11020 36320
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 10416 36236 10468 36242
rect 10416 36178 10468 36184
rect 10966 36136 11022 36145
rect 10966 36071 10968 36080
rect 11020 36071 11022 36080
rect 10968 36042 11020 36048
rect 10508 35488 10560 35494
rect 10508 35430 10560 35436
rect 10520 35086 10548 35430
rect 10324 35080 10376 35086
rect 10324 35022 10376 35028
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10876 35080 10928 35086
rect 10876 35022 10928 35028
rect 10336 34474 10364 35022
rect 10324 34468 10376 34474
rect 10324 34410 10376 34416
rect 10888 34406 10916 35022
rect 10980 34950 11008 36042
rect 11336 35760 11388 35766
rect 11336 35702 11388 35708
rect 11152 35692 11204 35698
rect 11152 35634 11204 35640
rect 11164 35290 11192 35634
rect 11152 35284 11204 35290
rect 11152 35226 11204 35232
rect 11348 35222 11376 35702
rect 11428 35624 11480 35630
rect 11428 35566 11480 35572
rect 11336 35216 11388 35222
rect 11336 35158 11388 35164
rect 11440 35154 11468 35566
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 10968 34944 11020 34950
rect 10968 34886 11020 34892
rect 10980 34785 11008 34886
rect 10966 34776 11022 34785
rect 10966 34711 11022 34720
rect 10876 34400 10928 34406
rect 10876 34342 10928 34348
rect 10968 34400 11020 34406
rect 10968 34342 11020 34348
rect 10888 34066 10916 34342
rect 10980 34202 11008 34342
rect 11256 34202 11284 34954
rect 11440 34746 11468 35090
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 10876 34060 10928 34066
rect 10876 34002 10928 34008
rect 11060 33992 11112 33998
rect 10506 33960 10562 33969
rect 11060 33934 11112 33940
rect 10428 33904 10506 33912
rect 10428 33884 10508 33904
rect 10322 32872 10378 32881
rect 10322 32807 10324 32816
rect 10376 32807 10378 32816
rect 10324 32778 10376 32784
rect 10336 32434 10364 32778
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 9128 32292 9180 32298
rect 9128 32234 9180 32240
rect 8772 32184 8984 32212
rect 8956 31754 8984 32184
rect 9324 32026 9352 32302
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 9324 31754 9352 31962
rect 8956 31726 9076 31754
rect 9324 31726 9444 31754
rect 8760 31680 8812 31686
rect 8760 31622 8812 31628
rect 8772 31346 8800 31622
rect 8942 31376 8998 31385
rect 8760 31340 8812 31346
rect 8942 31311 8944 31320
rect 8760 31282 8812 31288
rect 8996 31311 8998 31320
rect 8944 31282 8996 31288
rect 8668 31204 8720 31210
rect 8668 31146 8720 31152
rect 8956 30938 8984 31282
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 8576 30796 8628 30802
rect 8576 30738 8628 30744
rect 8588 29850 8616 30738
rect 8956 30598 8984 30874
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8758 30288 8814 30297
rect 8668 30252 8720 30258
rect 8814 30246 8892 30274
rect 8758 30223 8814 30232
rect 8668 30194 8720 30200
rect 8680 29850 8708 30194
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8668 29844 8720 29850
rect 8668 29786 8720 29792
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8354 27390 8524 27418
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8298 27367 8354 27376
rect 8206 27296 8262 27305
rect 8206 27231 8262 27240
rect 8298 27160 8354 27169
rect 8208 27124 8260 27130
rect 8588 27130 8616 27406
rect 8576 27124 8628 27130
rect 8354 27104 8524 27112
rect 8298 27095 8300 27104
rect 8208 27066 8260 27072
rect 8352 27084 8524 27104
rect 8300 27066 8352 27072
rect 8220 26586 8248 27066
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 8312 26450 8340 26862
rect 8404 26450 8432 26930
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7852 25078 8064 25106
rect 7760 24942 7880 24970
rect 7656 24880 7708 24886
rect 7562 24848 7618 24857
rect 7656 24822 7708 24828
rect 7562 24783 7618 24792
rect 7576 24614 7604 24783
rect 7748 24744 7800 24750
rect 7654 24712 7710 24721
rect 7748 24686 7800 24692
rect 7654 24647 7710 24656
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7564 24064 7616 24070
rect 7484 24024 7564 24052
rect 7564 24006 7616 24012
rect 7668 23866 7696 24647
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7378 23352 7434 23361
rect 7378 23287 7434 23296
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7248 22664 7328 22692
rect 7196 22646 7248 22652
rect 7392 22642 7420 23054
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 6828 22500 6880 22506
rect 6828 22442 6880 22448
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6748 21146 6776 22102
rect 6840 21962 6868 22442
rect 6932 22137 6960 22578
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6918 22128 6974 22137
rect 6918 22063 6974 22072
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 6840 21554 6868 21898
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6932 21185 6960 21830
rect 7024 21593 7052 22374
rect 7116 22166 7144 22578
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7392 22030 7420 22578
rect 7380 22024 7432 22030
rect 7286 21992 7342 22001
rect 7104 21956 7156 21962
rect 7380 21966 7432 21972
rect 7286 21927 7342 21936
rect 7104 21898 7156 21904
rect 7010 21584 7066 21593
rect 7010 21519 7066 21528
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 6918 21176 6974 21185
rect 6736 21140 6788 21146
rect 6918 21111 6920 21120
rect 6736 21082 6788 21088
rect 6972 21111 6974 21120
rect 6920 21082 6972 21088
rect 7024 20942 7052 21422
rect 7116 20942 7144 21898
rect 7300 21622 7328 21927
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7196 21412 7248 21418
rect 7196 21354 7248 21360
rect 7208 21049 7236 21354
rect 7288 21344 7340 21350
rect 7392 21321 7420 21490
rect 7288 21286 7340 21292
rect 7378 21312 7434 21321
rect 7300 21146 7328 21286
rect 7378 21247 7434 21256
rect 7484 21146 7512 23598
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7576 22545 7604 22918
rect 7668 22642 7696 22918
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7562 22536 7618 22545
rect 7562 22471 7618 22480
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7576 22273 7604 22374
rect 7562 22264 7618 22273
rect 7562 22199 7618 22208
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7380 21072 7432 21078
rect 7194 21040 7250 21049
rect 7380 21014 7432 21020
rect 7194 20975 7250 20984
rect 7208 20942 7236 20975
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7196 20936 7248 20942
rect 7392 20913 7420 21014
rect 7196 20878 7248 20884
rect 7378 20904 7434 20913
rect 6932 20806 6960 20878
rect 6828 20800 6880 20806
rect 6826 20768 6828 20777
rect 6920 20800 6972 20806
rect 6880 20768 6882 20777
rect 6920 20742 6972 20748
rect 6826 20703 6882 20712
rect 6826 20632 6882 20641
rect 6826 20567 6882 20576
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6748 19514 6776 20402
rect 6840 19786 6868 20567
rect 6918 20496 6974 20505
rect 6918 20431 6974 20440
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6274 18728 6330 18737
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 6012 18426 6040 18634
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5908 18352 5960 18358
rect 5960 18300 6040 18306
rect 5908 18294 6040 18300
rect 5816 18284 5868 18290
rect 5920 18278 6040 18294
rect 5816 18226 5868 18232
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5828 17678 5856 17750
rect 5920 17678 5948 18090
rect 5816 17672 5868 17678
rect 5722 17640 5778 17649
rect 5816 17614 5868 17620
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5722 17575 5724 17584
rect 5776 17575 5778 17584
rect 5724 17546 5776 17552
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5644 17270 5672 17478
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5184 17054 5396 17082
rect 5460 17066 5488 17206
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16794 5212 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 16250 5028 16526
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4080 16153 4108 16186
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4908 15994 4936 16050
rect 5172 16040 5224 16046
rect 4908 15988 5172 15994
rect 5224 15988 5304 15994
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15502 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4080 15026 4108 15438
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14618 4660 14962
rect 4724 14822 4752 15982
rect 4908 15966 5304 15988
rect 5276 15638 5304 15966
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5368 15502 5396 17054
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5644 16794 5672 17070
rect 5736 17066 5764 17546
rect 5920 17134 5948 17614
rect 6012 17270 6040 18278
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6104 17678 6132 18226
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 17338 6132 17478
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5998 17096 6054 17105
rect 5724 17060 5776 17066
rect 5998 17031 6054 17040
rect 5724 17002 5776 17008
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3804 13938 3832 14418
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3804 13530 3832 13874
rect 4632 13802 4660 13942
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 13738
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 1216 13388 1268 13394
rect 1216 13330 1268 13336
rect 1228 13161 1256 13330
rect 1214 13152 1270 13161
rect 1214 13087 1270 13096
rect 4264 12986 4292 13466
rect 4724 13326 4752 14758
rect 4816 14414 4844 15370
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5184 13530 5212 14486
rect 5276 14414 5304 15438
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5368 14346 5396 15438
rect 5552 15366 5580 16050
rect 5644 15706 5672 16390
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5736 15076 5764 17002
rect 5906 16960 5962 16969
rect 5906 16895 5962 16904
rect 5920 15502 5948 16895
rect 6012 16250 6040 17031
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6012 16046 6040 16186
rect 6104 16114 6132 17138
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6196 15570 6224 18702
rect 6274 18663 6276 18672
rect 6328 18663 6330 18672
rect 6276 18634 6328 18640
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 6196 15162 6224 15506
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5816 15088 5868 15094
rect 5736 15048 5816 15076
rect 5816 15030 5868 15036
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5828 13938 5856 14894
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6104 14006 6132 14214
rect 6196 14074 6224 14282
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 5184 12986 5212 13466
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5828 12918 5856 13874
rect 6288 13530 6316 18634
rect 6380 18358 6408 18770
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6472 18222 6500 19110
rect 6564 18766 6592 19178
rect 6552 18760 6604 18766
rect 6748 18714 6776 19450
rect 6932 19378 6960 20431
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6918 19136 6974 19145
rect 7024 19122 7052 20878
rect 7378 20839 7434 20848
rect 7288 20800 7340 20806
rect 7194 20768 7250 20777
rect 7116 20726 7194 20754
rect 7116 20466 7144 20726
rect 7576 20777 7604 21898
rect 7656 21412 7708 21418
rect 7656 21354 7708 21360
rect 7288 20742 7340 20748
rect 7562 20768 7618 20777
rect 7194 20703 7250 20712
rect 7300 20602 7328 20742
rect 7562 20703 7618 20712
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7300 20482 7328 20538
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7232 20454 7328 20482
rect 7378 20496 7434 20505
rect 7232 20244 7260 20454
rect 7378 20431 7434 20440
rect 7392 20398 7420 20431
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7208 20216 7260 20244
rect 7288 20256 7340 20262
rect 7208 19378 7236 20216
rect 7288 20198 7340 20204
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7300 19990 7328 20198
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7300 19553 7328 19790
rect 7286 19544 7342 19553
rect 7392 19514 7420 20198
rect 7472 19848 7524 19854
rect 7470 19816 7472 19825
rect 7524 19816 7526 19825
rect 7576 19802 7604 20334
rect 7668 20097 7696 21354
rect 7760 21010 7788 24686
rect 7852 23662 7880 24942
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7944 24614 7972 24754
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7944 24342 7972 24550
rect 7932 24336 7984 24342
rect 7932 24278 7984 24284
rect 7932 24200 7984 24206
rect 7930 24168 7932 24177
rect 7984 24168 7986 24177
rect 7930 24103 7986 24112
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7852 22506 7880 23462
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7944 22710 7972 23258
rect 8036 22710 8064 25078
rect 8128 24426 8156 26250
rect 8220 25838 8248 26318
rect 8298 26072 8354 26081
rect 8298 26007 8354 26016
rect 8312 25906 8340 26007
rect 8496 25974 8524 27084
rect 8576 27066 8628 27072
rect 8680 26994 8708 28562
rect 8760 27872 8812 27878
rect 8760 27814 8812 27820
rect 8772 27674 8800 27814
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 8864 26994 8892 30246
rect 8944 29096 8996 29102
rect 8944 29038 8996 29044
rect 8956 28490 8984 29038
rect 8944 28484 8996 28490
rect 8944 28426 8996 28432
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8956 27130 8984 27882
rect 9048 27849 9076 31726
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9220 30728 9272 30734
rect 9220 30670 9272 30676
rect 9232 30258 9260 30670
rect 9324 30666 9352 31214
rect 9312 30660 9364 30666
rect 9312 30602 9364 30608
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9232 29850 9260 30194
rect 9324 30190 9352 30602
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 9220 29844 9272 29850
rect 9220 29786 9272 29792
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9324 29306 9352 29582
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9126 29200 9182 29209
rect 9126 29135 9182 29144
rect 9220 29164 9272 29170
rect 9140 29034 9168 29135
rect 9220 29106 9272 29112
rect 9128 29028 9180 29034
rect 9128 28970 9180 28976
rect 9232 28558 9260 29106
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9324 28762 9352 29038
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9232 28218 9260 28494
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9220 28212 9272 28218
rect 9220 28154 9272 28160
rect 9034 27840 9090 27849
rect 9034 27775 9090 27784
rect 9140 27690 9168 28154
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9140 27662 9260 27690
rect 9232 27606 9260 27662
rect 9220 27600 9272 27606
rect 9220 27542 9272 27548
rect 9232 27470 9260 27542
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9140 27130 9168 27406
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 9232 27062 9260 27270
rect 9220 27056 9272 27062
rect 9220 26998 9272 27004
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8484 25968 8536 25974
rect 8482 25936 8484 25945
rect 8536 25936 8538 25945
rect 8300 25900 8352 25906
rect 8482 25871 8538 25880
rect 8300 25842 8352 25848
rect 8208 25832 8260 25838
rect 8208 25774 8260 25780
rect 8206 25528 8262 25537
rect 8206 25463 8262 25472
rect 8220 25294 8248 25463
rect 8312 25430 8340 25842
rect 8484 25764 8536 25770
rect 8484 25706 8536 25712
rect 8496 25498 8524 25706
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8300 25424 8352 25430
rect 8300 25366 8352 25372
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8220 24818 8248 25094
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8128 24398 8248 24426
rect 8220 24206 8248 24398
rect 8116 24200 8168 24206
rect 8114 24168 8116 24177
rect 8208 24200 8260 24206
rect 8168 24168 8170 24177
rect 8208 24142 8260 24148
rect 8114 24103 8170 24112
rect 8220 24041 8248 24142
rect 8206 24032 8262 24041
rect 8206 23967 8262 23976
rect 8208 23520 8260 23526
rect 8312 23508 8340 25366
rect 8588 25294 8616 25638
rect 8680 25480 8708 26930
rect 8772 26858 8800 26930
rect 9126 26888 9182 26897
rect 8760 26852 8812 26858
rect 9324 26858 9352 27950
rect 9126 26823 9182 26832
rect 9312 26852 9364 26858
rect 8760 26794 8812 26800
rect 8772 25770 8800 26794
rect 9140 26364 9168 26823
rect 9312 26794 9364 26800
rect 9416 26382 9444 31726
rect 9508 31686 9536 32302
rect 10324 32224 10376 32230
rect 10428 32212 10456 33884
rect 10560 33895 10562 33904
rect 10508 33866 10560 33872
rect 11072 33658 11100 33934
rect 11244 33856 11296 33862
rect 11532 33844 11560 36518
rect 11808 35714 11836 37198
rect 11888 37120 11940 37126
rect 11888 37062 11940 37068
rect 11900 36582 11928 37062
rect 11888 36576 11940 36582
rect 11888 36518 11940 36524
rect 11716 35686 11836 35714
rect 11900 35698 11928 36518
rect 11992 36242 12020 38354
rect 12164 37800 12216 37806
rect 12164 37742 12216 37748
rect 12176 37330 12204 37742
rect 12268 37738 12296 38354
rect 12256 37732 12308 37738
rect 12256 37674 12308 37680
rect 12164 37324 12216 37330
rect 12164 37266 12216 37272
rect 12164 37120 12216 37126
rect 12164 37062 12216 37068
rect 12072 36712 12124 36718
rect 12072 36654 12124 36660
rect 11980 36236 12032 36242
rect 11980 36178 12032 36184
rect 12084 36174 12112 36654
rect 12176 36378 12204 37062
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12072 36168 12124 36174
rect 12072 36110 12124 36116
rect 11888 35692 11940 35698
rect 11612 35556 11664 35562
rect 11612 35498 11664 35504
rect 11624 35170 11652 35498
rect 11716 35290 11744 35686
rect 11888 35634 11940 35640
rect 12360 35494 12388 38830
rect 12544 38350 12572 39238
rect 13004 39030 13032 40870
rect 13268 40588 13320 40594
rect 13268 40530 13320 40536
rect 13176 40384 13228 40390
rect 13176 40326 13228 40332
rect 13188 39030 13216 40326
rect 13280 40050 13308 40530
rect 13268 40044 13320 40050
rect 13268 39986 13320 39992
rect 13360 39840 13412 39846
rect 13280 39800 13360 39828
rect 12992 39024 13044 39030
rect 12992 38966 13044 38972
rect 13176 39024 13228 39030
rect 13176 38966 13228 38972
rect 13280 38894 13308 39800
rect 13360 39782 13412 39788
rect 13556 39642 13584 41006
rect 14096 40520 14148 40526
rect 14096 40462 14148 40468
rect 15108 40520 15160 40526
rect 15108 40462 15160 40468
rect 15936 40520 15988 40526
rect 15936 40462 15988 40468
rect 14108 40186 14136 40462
rect 14096 40180 14148 40186
rect 14096 40122 14148 40128
rect 13636 39976 13688 39982
rect 13636 39918 13688 39924
rect 13544 39636 13596 39642
rect 13544 39578 13596 39584
rect 13556 39030 13584 39578
rect 13544 39024 13596 39030
rect 13544 38966 13596 38972
rect 13268 38888 13320 38894
rect 13268 38830 13320 38836
rect 12624 38548 12676 38554
rect 12624 38490 12676 38496
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12636 37874 12664 38490
rect 12808 38208 12860 38214
rect 12808 38150 12860 38156
rect 12820 37874 12848 38150
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 12808 37868 12860 37874
rect 12808 37810 12860 37816
rect 12900 37460 12952 37466
rect 12900 37402 12952 37408
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12544 35834 12572 37062
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12636 35834 12664 36654
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 12532 35828 12584 35834
rect 12532 35770 12584 35776
rect 12624 35828 12676 35834
rect 12624 35770 12676 35776
rect 12716 35760 12768 35766
rect 12716 35702 12768 35708
rect 12348 35488 12400 35494
rect 12348 35430 12400 35436
rect 12728 35290 12756 35702
rect 12820 35562 12848 35974
rect 12808 35556 12860 35562
rect 12808 35498 12860 35504
rect 12820 35290 12848 35498
rect 11704 35284 11756 35290
rect 11704 35226 11756 35232
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 12624 35216 12676 35222
rect 11794 35184 11850 35193
rect 11624 35142 11794 35170
rect 12624 35158 12676 35164
rect 11794 35119 11850 35128
rect 11808 35086 11836 35119
rect 11796 35080 11848 35086
rect 11848 35040 11928 35068
rect 11796 35022 11848 35028
rect 11794 34640 11850 34649
rect 11794 34575 11850 34584
rect 11808 34542 11836 34575
rect 11796 34536 11848 34542
rect 11796 34478 11848 34484
rect 11900 34116 11928 35040
rect 12256 35012 12308 35018
rect 12256 34954 12308 34960
rect 12070 34776 12126 34785
rect 11992 34746 12070 34762
rect 11980 34740 12070 34746
rect 12032 34734 12070 34740
rect 12070 34711 12126 34720
rect 11980 34682 12032 34688
rect 12162 34640 12218 34649
rect 12162 34575 12164 34584
rect 12216 34575 12218 34584
rect 12164 34546 12216 34552
rect 12268 34202 12296 34954
rect 12440 34400 12492 34406
rect 12492 34360 12572 34388
rect 12440 34342 12492 34348
rect 12256 34196 12308 34202
rect 12256 34138 12308 34144
rect 11702 34096 11758 34105
rect 11900 34088 12020 34116
rect 11758 34040 11928 34048
rect 11702 34031 11704 34040
rect 11756 34020 11928 34040
rect 11704 34002 11756 34008
rect 11244 33798 11296 33804
rect 11440 33816 11560 33844
rect 11060 33652 11112 33658
rect 11060 33594 11112 33600
rect 11256 33522 11284 33798
rect 11334 33552 11390 33561
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10692 33516 10744 33522
rect 10692 33458 10744 33464
rect 11244 33516 11296 33522
rect 11334 33487 11390 33496
rect 11244 33458 11296 33464
rect 10612 33114 10640 33458
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10520 32366 10548 33050
rect 10704 32774 10732 33458
rect 11060 33448 11112 33454
rect 11060 33390 11112 33396
rect 10968 33380 11020 33386
rect 10968 33322 11020 33328
rect 10876 33312 10928 33318
rect 10980 33289 11008 33322
rect 10876 33254 10928 33260
rect 10966 33280 11022 33289
rect 10692 32768 10744 32774
rect 10692 32710 10744 32716
rect 10508 32360 10560 32366
rect 10508 32302 10560 32308
rect 10888 32280 10916 33254
rect 10966 33215 11022 33224
rect 11072 32910 11100 33390
rect 11256 33046 11284 33458
rect 11348 33454 11376 33487
rect 11336 33448 11388 33454
rect 11336 33390 11388 33396
rect 11244 33040 11296 33046
rect 11244 32982 11296 32988
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 11152 32564 11204 32570
rect 11152 32506 11204 32512
rect 10968 32292 11020 32298
rect 10888 32252 10968 32280
rect 10968 32234 11020 32240
rect 10428 32184 10548 32212
rect 10324 32166 10376 32172
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9678 31784 9734 31793
rect 9496 31680 9548 31686
rect 9496 31622 9548 31628
rect 9508 30818 9536 31622
rect 9600 31346 9628 31758
rect 9678 31719 9734 31728
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 9508 30790 9628 30818
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9508 30190 9536 30670
rect 9600 30394 9628 30790
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 30184 9548 30190
rect 9496 30126 9548 30132
rect 9508 29306 9536 30126
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9494 29200 9550 29209
rect 9494 29135 9496 29144
rect 9548 29135 9550 29144
rect 9496 29106 9548 29112
rect 9692 29050 9720 31719
rect 10048 31680 10100 31686
rect 10048 31622 10100 31628
rect 10336 31634 10364 32166
rect 10520 31754 10548 32184
rect 10980 31822 11008 32234
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10520 31726 10732 31754
rect 10598 31648 10654 31657
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9876 30938 9904 31214
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 10060 30734 10088 31622
rect 10336 31606 10598 31634
rect 10598 31583 10654 31592
rect 10140 31476 10192 31482
rect 10140 31418 10192 31424
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 10060 30433 10088 30670
rect 10046 30424 10102 30433
rect 9864 30388 9916 30394
rect 10046 30359 10102 30368
rect 9864 30330 9916 30336
rect 9876 29345 9904 30330
rect 9956 30252 10008 30258
rect 9956 30194 10008 30200
rect 9968 29646 9996 30194
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9862 29336 9918 29345
rect 9862 29271 9918 29280
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9508 29022 9720 29050
rect 9508 27946 9536 29022
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9496 27940 9548 27946
rect 9496 27882 9548 27888
rect 9508 27130 9536 27882
rect 9600 27713 9628 28562
rect 9680 28484 9732 28490
rect 9784 28472 9812 29106
rect 9876 28642 9904 29271
rect 9968 28762 9996 29582
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 9876 28614 9996 28642
rect 9732 28444 9812 28472
rect 9680 28426 9732 28432
rect 9692 27946 9720 28426
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9586 27704 9642 27713
rect 9876 27674 9904 28018
rect 9586 27639 9642 27648
rect 9864 27668 9916 27674
rect 9600 27470 9628 27639
rect 9864 27610 9916 27616
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9692 26790 9720 27270
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9220 26376 9272 26382
rect 9140 26336 9220 26364
rect 9220 26318 9272 26324
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 8852 26308 8904 26314
rect 9036 26308 9088 26314
rect 8904 26268 8984 26296
rect 8852 26250 8904 26256
rect 8760 25764 8812 25770
rect 8760 25706 8812 25712
rect 8760 25492 8812 25498
rect 8680 25452 8760 25480
rect 8760 25434 8812 25440
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8392 25220 8444 25226
rect 8668 25220 8720 25226
rect 8444 25180 8524 25208
rect 8392 25162 8444 25168
rect 8390 24576 8446 24585
rect 8390 24511 8446 24520
rect 8404 24138 8432 24511
rect 8496 24138 8524 25180
rect 8668 25162 8720 25168
rect 8680 24954 8708 25162
rect 8668 24948 8720 24954
rect 8720 24908 8892 24936
rect 8668 24890 8720 24896
rect 8760 24812 8812 24818
rect 8588 24772 8760 24800
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8484 24132 8536 24138
rect 8484 24074 8536 24080
rect 8260 23480 8340 23508
rect 8208 23462 8260 23468
rect 8220 22982 8248 23462
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 7944 21962 7972 22170
rect 8036 22098 8064 22646
rect 8128 22234 8156 22918
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 7932 21956 7984 21962
rect 7932 21898 7984 21904
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21554 7880 21830
rect 7944 21729 7972 21898
rect 7930 21720 7986 21729
rect 7930 21655 7986 21664
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 7930 21584 7986 21593
rect 7840 21548 7892 21554
rect 7930 21519 7986 21528
rect 7840 21490 7892 21496
rect 7944 21146 7972 21519
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7654 20088 7710 20097
rect 7654 20023 7710 20032
rect 7760 19961 7788 20946
rect 7746 19952 7802 19961
rect 7746 19887 7802 19896
rect 7746 19816 7802 19825
rect 7576 19774 7746 19802
rect 7470 19751 7526 19760
rect 7746 19751 7802 19760
rect 7286 19479 7342 19488
rect 7380 19508 7432 19514
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7300 19242 7328 19479
rect 7380 19450 7432 19456
rect 7378 19408 7434 19417
rect 7378 19343 7434 19352
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 6974 19094 7052 19122
rect 7194 19136 7250 19145
rect 6918 19071 6974 19080
rect 7194 19071 7250 19080
rect 6552 18702 6604 18708
rect 6656 18686 6776 18714
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6564 18329 6592 18566
rect 6550 18320 6606 18329
rect 6550 18255 6606 18264
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6472 17814 6500 18158
rect 6460 17808 6512 17814
rect 6460 17750 6512 17756
rect 6368 17672 6420 17678
rect 6564 17660 6592 18255
rect 6656 17814 6684 18686
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6748 18154 6776 18566
rect 6932 18358 6960 18566
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6840 17882 6868 18158
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6368 17614 6420 17620
rect 6472 17632 6592 17660
rect 6380 17338 6408 17614
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6472 17202 6500 17632
rect 6656 17610 6684 17750
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6564 16590 6592 17478
rect 6656 17184 6684 17546
rect 6840 17338 6868 17818
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 17196 6788 17202
rect 6656 17156 6736 17184
rect 6736 17138 6788 17144
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6458 16144 6514 16153
rect 6458 16079 6460 16088
rect 6512 16079 6514 16088
rect 6460 16050 6512 16056
rect 6748 15094 6776 17138
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6644 14476 6696 14482
rect 6748 14464 6776 15030
rect 6840 14958 6868 15302
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6932 14618 6960 18158
rect 7024 17649 7052 18702
rect 7208 18086 7236 19071
rect 7392 18630 7420 19343
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7286 18320 7342 18329
rect 7286 18255 7288 18264
rect 7340 18255 7342 18264
rect 7288 18226 7340 18232
rect 7196 18080 7248 18086
rect 7102 18048 7158 18057
rect 7196 18022 7248 18028
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7102 17983 7158 17992
rect 7010 17640 7066 17649
rect 7010 17575 7066 17584
rect 7116 17270 7144 17983
rect 7194 17912 7250 17921
rect 7194 17847 7250 17856
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 7208 17202 7236 17847
rect 7300 17746 7328 18022
rect 7392 17746 7420 18362
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7286 17504 7342 17513
rect 7286 17439 7342 17448
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7024 16658 7052 16934
rect 7208 16726 7236 17138
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6696 14436 6776 14464
rect 6644 14418 6696 14424
rect 6748 13802 6776 14436
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 1216 12300 1268 12306
rect 1216 12242 1268 12248
rect 1228 12073 1256 12242
rect 6840 12238 6868 14010
rect 6932 14006 6960 14554
rect 7024 14414 7052 14758
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7116 14074 7144 15846
rect 7300 15706 7328 17439
rect 7484 16590 7512 19751
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7668 18630 7696 19178
rect 7852 18970 7880 21082
rect 8036 21010 8064 21626
rect 8128 21185 8156 21898
rect 8220 21894 8248 22918
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8390 22400 8446 22409
rect 8312 22273 8340 22374
rect 8390 22335 8446 22344
rect 8298 22264 8354 22273
rect 8298 22199 8354 22208
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8312 21622 8340 22034
rect 8404 22030 8432 22335
rect 8496 22030 8524 22578
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8404 21865 8432 21966
rect 8390 21856 8446 21865
rect 8588 21842 8616 24772
rect 8760 24754 8812 24760
rect 8668 24336 8720 24342
rect 8668 24278 8720 24284
rect 8680 23866 8708 24278
rect 8760 24132 8812 24138
rect 8760 24074 8812 24080
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8680 22030 8708 23190
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8390 21791 8446 21800
rect 8496 21814 8616 21842
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8114 21176 8170 21185
rect 8114 21111 8170 21120
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 8220 20913 8248 21490
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 8300 20936 8352 20942
rect 8022 20904 8078 20913
rect 8022 20839 8024 20848
rect 8076 20839 8078 20848
rect 8206 20904 8262 20913
rect 8300 20878 8352 20884
rect 8206 20839 8262 20848
rect 8024 20810 8076 20816
rect 8312 20641 8340 20878
rect 8404 20874 8432 21354
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8298 20632 8354 20641
rect 7932 20596 7984 20602
rect 8298 20567 8354 20576
rect 7932 20538 7984 20544
rect 7944 20505 7972 20538
rect 8392 20528 8444 20534
rect 7930 20496 7986 20505
rect 7930 20431 7986 20440
rect 8390 20496 8392 20505
rect 8444 20496 8446 20505
rect 8496 20466 8524 21814
rect 8574 21720 8630 21729
rect 8574 21655 8630 21664
rect 8390 20431 8446 20440
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8208 20392 8260 20398
rect 7944 20352 8208 20380
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7944 18698 7972 20352
rect 8208 20334 8260 20340
rect 8392 20392 8444 20398
rect 8496 20369 8524 20402
rect 8392 20334 8444 20340
rect 8482 20360 8538 20369
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8036 20058 8064 20198
rect 8206 20088 8262 20097
rect 8024 20052 8076 20058
rect 8206 20023 8262 20032
rect 8024 19994 8076 20000
rect 8220 19854 8248 20023
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8114 19544 8170 19553
rect 8114 19479 8170 19488
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7576 18290 7604 18566
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7472 16584 7524 16590
rect 7378 16552 7434 16561
rect 7472 16526 7524 16532
rect 7378 16487 7434 16496
rect 7392 16114 7420 16487
rect 7484 16130 7512 16526
rect 7576 16250 7604 17070
rect 7668 16697 7696 18566
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7748 18080 7800 18086
rect 7746 18048 7748 18057
rect 7800 18048 7802 18057
rect 7746 17983 7802 17992
rect 7944 17882 7972 18362
rect 8128 18306 8156 19479
rect 8220 18766 8248 19790
rect 8312 19514 8340 20198
rect 8404 19718 8432 20334
rect 8482 20295 8538 20304
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8496 19514 8524 19722
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8390 19000 8446 19009
rect 8390 18935 8392 18944
rect 8444 18935 8446 18944
rect 8392 18906 8444 18912
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18358 8248 18566
rect 8036 18278 8156 18306
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7760 17338 7788 17546
rect 7852 17338 7880 17614
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7944 17270 7972 17478
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7654 16688 7710 16697
rect 7654 16623 7710 16632
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7380 16108 7432 16114
rect 7484 16102 7604 16130
rect 7380 16050 7432 16056
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 15026 7420 15302
rect 7484 15162 7512 15982
rect 7576 15162 7604 16102
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13734 6960 13806
rect 7392 13734 7420 14758
rect 7576 14414 7604 15098
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7668 14278 7696 16623
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 14958 7788 15846
rect 8036 15706 8064 18278
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17814 8156 18158
rect 8206 17912 8262 17921
rect 8206 17847 8262 17856
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8128 17270 8156 17750
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8220 16114 8248 17847
rect 8312 17746 8340 18838
rect 8392 18624 8444 18630
rect 8390 18592 8392 18601
rect 8444 18592 8446 18601
rect 8390 18527 8446 18536
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 18057 8432 18226
rect 8390 18048 8446 18057
rect 8390 17983 8446 17992
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17066 8340 17682
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16522 8340 17002
rect 8404 16590 8432 17478
rect 8496 17338 8524 18362
rect 8588 17542 8616 21655
rect 8680 21554 8708 21966
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8772 21434 8800 24074
rect 8864 23322 8892 24908
rect 8956 24290 8984 26268
rect 9036 26250 9088 26256
rect 9048 26042 9076 26250
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9048 24954 9076 25842
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9324 25294 9352 25638
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 9034 24848 9090 24857
rect 9034 24783 9036 24792
rect 9088 24783 9090 24792
rect 9128 24812 9180 24818
rect 9036 24754 9088 24760
rect 9128 24754 9180 24760
rect 9140 24410 9168 24754
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 8956 24262 9168 24290
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8956 23866 8984 24142
rect 9048 24041 9076 24142
rect 9034 24032 9090 24041
rect 9034 23967 9090 23976
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 9036 23656 9088 23662
rect 8956 23604 9036 23610
rect 8956 23598 9088 23604
rect 8956 23582 9076 23598
rect 9140 23594 9168 24262
rect 9232 23662 9260 25230
rect 9416 24834 9444 26318
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9508 25294 9536 25978
rect 9770 25800 9826 25809
rect 9770 25735 9826 25744
rect 9586 25392 9642 25401
rect 9586 25327 9642 25336
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9324 24818 9444 24834
rect 9312 24812 9444 24818
rect 9364 24806 9444 24812
rect 9312 24754 9364 24760
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 24274 9352 24550
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9128 23588 9180 23594
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 22166 8892 22578
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8864 21690 8892 21830
rect 8956 21729 8984 23582
rect 9128 23530 9180 23536
rect 9034 22672 9090 22681
rect 9034 22607 9036 22616
rect 9088 22607 9090 22616
rect 9128 22636 9180 22642
rect 9036 22578 9088 22584
rect 9128 22578 9180 22584
rect 9140 22522 9168 22578
rect 9048 22494 9168 22522
rect 9048 22030 9076 22494
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22098 9168 22374
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 9036 22024 9088 22030
rect 9324 21978 9352 24074
rect 9416 23474 9444 24806
rect 9496 24812 9548 24818
rect 9600 24800 9628 25327
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9548 24772 9628 24800
rect 9496 24754 9548 24760
rect 9494 24440 9550 24449
rect 9692 24426 9720 24822
rect 9784 24614 9812 25735
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 25129 9904 25230
rect 9862 25120 9918 25129
rect 9862 25055 9918 25064
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9876 24818 9904 24890
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9550 24398 9720 24426
rect 9494 24375 9550 24384
rect 9692 24206 9720 24398
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9770 24032 9826 24041
rect 9508 23798 9536 24006
rect 9770 23967 9826 23976
rect 9784 23866 9812 23967
rect 9876 23866 9904 24550
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9496 23792 9548 23798
rect 9496 23734 9548 23740
rect 9968 23526 9996 28614
rect 10152 27614 10180 31418
rect 10612 30938 10640 31583
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10612 30802 10640 30874
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10612 30394 10640 30738
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10230 29744 10286 29753
rect 10230 29679 10286 29688
rect 10244 29510 10272 29679
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10336 29306 10364 29446
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 10336 28762 10364 29242
rect 10428 29238 10456 30194
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10520 29238 10548 29786
rect 10416 29232 10468 29238
rect 10416 29174 10468 29180
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 10508 28688 10560 28694
rect 10508 28630 10560 28636
rect 10520 28150 10548 28630
rect 10612 28218 10640 28902
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 10324 28008 10376 28014
rect 10324 27950 10376 27956
rect 10416 28008 10468 28014
rect 10416 27950 10468 27956
rect 10232 27940 10284 27946
rect 10232 27882 10284 27888
rect 10060 27586 10180 27614
rect 10060 26042 10088 27586
rect 10244 27538 10272 27882
rect 10336 27674 10364 27950
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10428 27554 10456 27950
rect 10704 27614 10732 31726
rect 10980 31142 11008 31758
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10796 30802 10824 31078
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10796 30394 10824 30738
rect 10876 30660 10928 30666
rect 10876 30602 10928 30608
rect 10784 30388 10836 30394
rect 10784 30330 10836 30336
rect 10888 30258 10916 30602
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10796 28558 10824 29582
rect 10874 29200 10930 29209
rect 10874 29135 10876 29144
rect 10928 29135 10930 29144
rect 10876 29106 10928 29112
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10796 28218 10824 28494
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10704 27586 10916 27614
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10336 27526 10456 27554
rect 10140 27464 10192 27470
rect 10336 27418 10364 27526
rect 10140 27406 10192 27412
rect 10152 27130 10180 27406
rect 10244 27390 10364 27418
rect 10414 27432 10470 27441
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 10244 25430 10272 27390
rect 10414 27367 10416 27376
rect 10468 27367 10470 27376
rect 10692 27396 10744 27402
rect 10416 27338 10468 27344
rect 10692 27338 10744 27344
rect 10428 26976 10456 27338
rect 10704 27130 10732 27338
rect 10782 27160 10838 27169
rect 10692 27124 10744 27130
rect 10782 27095 10838 27104
rect 10692 27066 10744 27072
rect 10600 26988 10652 26994
rect 10428 26948 10600 26976
rect 10600 26930 10652 26936
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10324 26240 10376 26246
rect 10324 26182 10376 26188
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10336 26042 10364 26182
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10336 25294 10364 25978
rect 10520 25906 10548 26182
rect 10508 25900 10560 25906
rect 10508 25842 10560 25848
rect 10324 25288 10376 25294
rect 10244 25248 10324 25276
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 9956 23520 10008 23526
rect 9416 23446 9812 23474
rect 9956 23462 10008 23468
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9586 22944 9642 22953
rect 9416 22902 9586 22930
rect 9416 22642 9444 22902
rect 9586 22879 9642 22888
rect 9692 22658 9720 23258
rect 9508 22642 9720 22658
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9496 22636 9720 22642
rect 9548 22630 9720 22636
rect 9784 22658 9812 23446
rect 9784 22630 9904 22658
rect 9496 22578 9548 22584
rect 9416 22234 9444 22578
rect 9772 22568 9824 22574
rect 9494 22536 9550 22545
rect 9772 22510 9824 22516
rect 9494 22471 9550 22480
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9402 22128 9458 22137
rect 9508 22098 9536 22471
rect 9680 22432 9732 22438
rect 9600 22392 9680 22420
rect 9402 22063 9458 22072
rect 9496 22092 9548 22098
rect 9416 22030 9444 22063
rect 9496 22034 9548 22040
rect 9036 21966 9088 21972
rect 8942 21720 8998 21729
rect 8852 21684 8904 21690
rect 8942 21655 8998 21664
rect 8852 21626 8904 21632
rect 8942 21584 8998 21593
rect 8864 21542 8942 21570
rect 8864 21486 8892 21542
rect 8942 21519 8998 21528
rect 8680 21406 8800 21434
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 21412 8996 21418
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8680 17202 8708 21406
rect 8944 21354 8996 21360
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8864 20942 8892 21286
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8772 19825 8800 20266
rect 8758 19816 8814 19825
rect 8864 19786 8892 20402
rect 8758 19751 8814 19760
rect 8852 19780 8904 19786
rect 8772 19514 8800 19751
rect 8852 19722 8904 19728
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8772 18970 8800 19178
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8864 18698 8892 19110
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 17882 8800 18158
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8864 17746 8892 18090
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16590 8524 17070
rect 8680 16794 8708 17138
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8496 16250 8524 16526
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7838 15192 7894 15201
rect 8036 15162 8064 15642
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7838 15127 7894 15136
rect 8024 15156 8076 15162
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 6932 12986 6960 13670
rect 7392 13462 7420 13670
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 1214 12064 1270 12073
rect 1214 11999 1270 12008
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10985 1900 11154
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 1216 10124 1268 10130
rect 1216 10066 1268 10072
rect 1228 9897 1256 10066
rect 1214 9888 1270 9897
rect 1214 9823 1270 9832
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1228 8809 1256 8978
rect 3146 8936 3202 8945
rect 3146 8871 3202 8880
rect 1214 8800 1270 8809
rect 1214 8735 1270 8744
rect 1216 7948 1268 7954
rect 1216 7890 1268 7896
rect 1228 7721 1256 7890
rect 1214 7712 1270 7721
rect 1214 7647 1270 7656
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1228 6633 1256 6802
rect 1214 6624 1270 6633
rect 1214 6559 1270 6568
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5545 1900 5714
rect 1858 5536 1914 5545
rect 1858 5471 1914 5480
rect 3160 4826 3188 8871
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 11698
rect 7760 11150 7788 14894
rect 7852 14074 7880 15127
rect 8024 15098 8076 15104
rect 8128 14618 8156 15506
rect 8496 15026 8524 15846
rect 8772 15706 8800 15982
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8956 15502 8984 21354
rect 9048 21350 9076 21966
rect 9140 21950 9352 21978
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9496 21956 9548 21962
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 9048 20602 9076 20878
rect 9036 20596 9088 20602
rect 9036 20538 9088 20544
rect 9048 20058 9076 20538
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9048 19242 9076 19994
rect 9140 19922 9168 21950
rect 9496 21898 9548 21904
rect 9404 21888 9456 21894
rect 9310 21856 9366 21865
rect 9404 21830 9456 21836
rect 9310 21791 9366 21800
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9232 20398 9260 21626
rect 9324 21554 9352 21791
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9416 21457 9444 21830
rect 9508 21690 9536 21898
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9496 21480 9548 21486
rect 9402 21448 9458 21457
rect 9496 21422 9548 21428
rect 9402 21383 9458 21392
rect 9402 21040 9458 21049
rect 9402 20975 9458 20984
rect 9416 20942 9444 20975
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9508 20874 9536 21422
rect 9600 21010 9628 22392
rect 9680 22374 9732 22380
rect 9784 22234 9812 22510
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9680 21888 9732 21894
rect 9876 21842 9904 22630
rect 9968 22438 9996 23462
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9732 21836 9904 21842
rect 9680 21830 9904 21836
rect 9692 21814 9904 21830
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9496 20528 9548 20534
rect 9402 20496 9458 20505
rect 9312 20460 9364 20466
rect 9496 20470 9548 20476
rect 9402 20431 9404 20440
rect 9312 20402 9364 20408
rect 9456 20431 9458 20440
rect 9404 20402 9456 20408
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9128 19372 9180 19378
rect 9232 19360 9260 20334
rect 9324 20233 9352 20402
rect 9310 20224 9366 20233
rect 9310 20159 9366 20168
rect 9416 19514 9444 20402
rect 9508 19514 9536 20470
rect 9600 19689 9628 20742
rect 9692 19854 9720 21814
rect 9770 21720 9826 21729
rect 9770 21655 9826 21664
rect 9784 21350 9812 21655
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 20806 9812 21286
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9770 20496 9826 20505
rect 9770 20431 9772 20440
rect 9824 20431 9826 20440
rect 9772 20402 9824 20408
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9784 19922 9812 20266
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9586 19680 9642 19689
rect 9586 19615 9642 19624
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9312 19372 9364 19378
rect 9232 19332 9312 19360
rect 9128 19314 9180 19320
rect 9312 19314 9364 19320
rect 9140 19242 9168 19314
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 9876 18873 9904 20878
rect 9862 18864 9918 18873
rect 9862 18799 9918 18808
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9126 18592 9182 18601
rect 9048 18426 9076 18566
rect 9182 18550 9260 18578
rect 9126 18527 9182 18536
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9232 18290 9260 18550
rect 9416 18290 9444 18702
rect 9968 18612 9996 22102
rect 10060 21622 10088 22646
rect 10152 22137 10180 25162
rect 10244 24857 10272 25248
rect 10324 25230 10376 25236
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10230 24848 10286 24857
rect 10230 24783 10286 24792
rect 10244 24342 10272 24783
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10336 22778 10364 22986
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10232 22500 10284 22506
rect 10232 22442 10284 22448
rect 10138 22128 10194 22137
rect 10138 22063 10194 22072
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10152 21865 10180 21898
rect 10138 21856 10194 21865
rect 10138 21791 10194 21800
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 10060 20942 10088 21558
rect 10244 21146 10272 22442
rect 10324 22432 10376 22438
rect 10428 22409 10456 25094
rect 10520 24682 10548 25842
rect 10612 25294 10640 26386
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10508 24676 10560 24682
rect 10508 24618 10560 24624
rect 10520 24342 10548 24618
rect 10612 24426 10640 25094
rect 10704 24614 10732 25910
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10690 24440 10746 24449
rect 10612 24398 10690 24426
rect 10690 24375 10746 24384
rect 10508 24336 10560 24342
rect 10508 24278 10560 24284
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10324 22374 10376 22380
rect 10414 22400 10470 22409
rect 10336 21146 10364 22374
rect 10414 22335 10470 22344
rect 10520 22080 10548 23598
rect 10704 23526 10732 24142
rect 10796 23730 10824 27095
rect 10888 26450 10916 27586
rect 10980 26466 11008 31078
rect 11164 30274 11192 32506
rect 11334 30288 11390 30297
rect 11164 30246 11334 30274
rect 11334 30223 11336 30232
rect 11388 30223 11390 30232
rect 11336 30194 11388 30200
rect 11336 30116 11388 30122
rect 11336 30058 11388 30064
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 11152 29572 11204 29578
rect 11152 29514 11204 29520
rect 11058 29200 11114 29209
rect 11164 29170 11192 29514
rect 11256 29306 11284 29650
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11348 29238 11376 30058
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 11058 29135 11060 29144
rect 11112 29135 11114 29144
rect 11152 29164 11204 29170
rect 11060 29106 11112 29112
rect 11152 29106 11204 29112
rect 11072 28966 11100 29106
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11164 28762 11192 29106
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 11164 28472 11192 28698
rect 11244 28484 11296 28490
rect 11164 28444 11244 28472
rect 11244 28426 11296 28432
rect 11244 28144 11296 28150
rect 11244 28086 11296 28092
rect 11060 28008 11112 28014
rect 11112 27968 11192 27996
rect 11060 27950 11112 27956
rect 11058 27704 11114 27713
rect 11164 27674 11192 27968
rect 11058 27639 11114 27648
rect 11152 27668 11204 27674
rect 11072 27470 11100 27639
rect 11152 27610 11204 27616
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11164 26994 11192 27610
rect 11256 27470 11284 28086
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11256 27130 11284 27406
rect 11348 27334 11376 28018
rect 11440 27418 11468 33816
rect 11520 33652 11572 33658
rect 11520 33594 11572 33600
rect 11532 32842 11560 33594
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11716 33425 11744 33458
rect 11702 33416 11758 33425
rect 11702 33351 11758 33360
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11520 32836 11572 32842
rect 11520 32778 11572 32784
rect 11624 31958 11652 32846
rect 11716 32570 11744 33050
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 11808 32026 11836 32846
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11612 31952 11664 31958
rect 11900 31906 11928 34020
rect 11612 31894 11664 31900
rect 11716 31878 11928 31906
rect 11716 31770 11744 31878
rect 11992 31804 12020 34088
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 12164 33992 12216 33998
rect 12440 33992 12492 33998
rect 12164 33934 12216 33940
rect 12438 33960 12440 33969
rect 12492 33960 12494 33969
rect 12084 33504 12112 33934
rect 12176 33658 12204 33934
rect 12438 33895 12494 33904
rect 12544 33810 12572 34360
rect 12636 34134 12664 35158
rect 12808 34944 12860 34950
rect 12808 34886 12860 34892
rect 12820 34610 12848 34886
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12808 34468 12860 34474
rect 12808 34410 12860 34416
rect 12624 34128 12676 34134
rect 12624 34070 12676 34076
rect 12820 33998 12848 34410
rect 12912 34048 12940 37402
rect 13280 37398 13308 38830
rect 13360 38752 13412 38758
rect 13360 38694 13412 38700
rect 13268 37392 13320 37398
rect 13268 37334 13320 37340
rect 13176 37256 13228 37262
rect 13176 37198 13228 37204
rect 13188 37126 13216 37198
rect 12992 37120 13044 37126
rect 12992 37062 13044 37068
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13004 36922 13032 37062
rect 12992 36916 13044 36922
rect 12992 36858 13044 36864
rect 13188 36666 13216 37062
rect 13096 36638 13216 36666
rect 13096 36038 13124 36638
rect 13176 36576 13228 36582
rect 13176 36518 13228 36524
rect 13084 36032 13136 36038
rect 13084 35974 13136 35980
rect 12992 35488 13044 35494
rect 12992 35430 13044 35436
rect 13004 35290 13032 35430
rect 12992 35284 13044 35290
rect 12992 35226 13044 35232
rect 13096 35068 13124 35974
rect 13188 35834 13216 36518
rect 13176 35828 13228 35834
rect 13176 35770 13228 35776
rect 13280 35630 13308 37334
rect 13372 37262 13400 38694
rect 13648 38554 13676 39918
rect 13820 39840 13872 39846
rect 13820 39782 13872 39788
rect 13832 39098 13860 39782
rect 14108 39098 14136 40122
rect 14740 40044 14792 40050
rect 14740 39986 14792 39992
rect 14648 39432 14700 39438
rect 14648 39374 14700 39380
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 14096 39092 14148 39098
rect 14096 39034 14148 39040
rect 14660 38962 14688 39374
rect 14648 38956 14700 38962
rect 14648 38898 14700 38904
rect 14280 38888 14332 38894
rect 14280 38830 14332 38836
rect 13636 38548 13688 38554
rect 13636 38490 13688 38496
rect 14188 38412 14240 38418
rect 14188 38354 14240 38360
rect 13820 38344 13872 38350
rect 13820 38286 13872 38292
rect 13636 37664 13688 37670
rect 13636 37606 13688 37612
rect 13648 37330 13676 37606
rect 13636 37324 13688 37330
rect 13636 37266 13688 37272
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 13372 36378 13400 36722
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 13268 35624 13320 35630
rect 13266 35592 13268 35601
rect 13320 35592 13322 35601
rect 13266 35527 13322 35536
rect 13372 35222 13400 36314
rect 13452 36032 13504 36038
rect 13452 35974 13504 35980
rect 13360 35216 13412 35222
rect 13360 35158 13412 35164
rect 13464 35154 13492 35974
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13176 35080 13228 35086
rect 13096 35040 13176 35068
rect 13176 35022 13228 35028
rect 13084 34740 13136 34746
rect 13084 34682 13136 34688
rect 13096 34542 13124 34682
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 12992 34400 13044 34406
rect 13044 34360 13492 34388
rect 12992 34342 13044 34348
rect 13266 34096 13322 34105
rect 12912 34020 13032 34048
rect 13266 34031 13268 34040
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 12452 33782 12572 33810
rect 12164 33652 12216 33658
rect 12164 33594 12216 33600
rect 12254 33552 12310 33561
rect 12164 33516 12216 33522
rect 12084 33476 12164 33504
rect 12254 33487 12256 33496
rect 12164 33458 12216 33464
rect 12308 33487 12310 33496
rect 12348 33516 12400 33522
rect 12256 33458 12308 33464
rect 12452 33504 12480 33782
rect 12532 33652 12584 33658
rect 12728 33640 12756 33866
rect 12584 33612 12756 33640
rect 12532 33594 12584 33600
rect 12716 33516 12768 33522
rect 12452 33476 12664 33504
rect 12348 33458 12400 33464
rect 12176 33318 12204 33458
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12256 32972 12308 32978
rect 12360 32960 12388 33458
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 12308 32932 12388 32960
rect 12256 32914 12308 32920
rect 12164 32904 12216 32910
rect 12216 32852 12388 32858
rect 12164 32846 12388 32852
rect 12176 32842 12388 32846
rect 12544 32842 12572 33322
rect 12176 32836 12400 32842
rect 12176 32830 12348 32836
rect 12348 32778 12400 32784
rect 12532 32836 12584 32842
rect 12532 32778 12584 32784
rect 12072 32768 12124 32774
rect 12072 32710 12124 32716
rect 12084 32230 12112 32710
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 12256 32020 12308 32026
rect 12256 31962 12308 31968
rect 11532 31742 11744 31770
rect 11808 31776 12020 31804
rect 11532 31482 11560 31742
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 11612 31340 11664 31346
rect 11612 31282 11664 31288
rect 11624 30938 11652 31282
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 11532 29170 11560 30194
rect 11624 29850 11652 30194
rect 11612 29844 11664 29850
rect 11612 29786 11664 29792
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11532 28762 11560 29106
rect 11624 28966 11652 29242
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11520 28756 11572 28762
rect 11520 28698 11572 28704
rect 11716 28608 11744 31078
rect 11532 28580 11744 28608
rect 11532 27826 11560 28580
rect 11808 28506 11836 31776
rect 12072 31680 12124 31686
rect 12268 31657 12296 31962
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12072 31622 12124 31628
rect 12254 31648 12310 31657
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11900 30394 11928 30738
rect 12084 30666 12112 31622
rect 12254 31583 12310 31592
rect 12360 31124 12388 31758
rect 12636 31754 12664 33476
rect 12820 33504 12848 33934
rect 12768 33476 12848 33504
rect 12900 33516 12952 33522
rect 12716 33458 12768 33464
rect 12900 33458 12952 33464
rect 12714 33416 12770 33425
rect 12714 33351 12770 33360
rect 12808 33380 12860 33386
rect 12728 33114 12756 33351
rect 12808 33322 12860 33328
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12820 32774 12848 33322
rect 12912 32978 12940 33458
rect 12900 32972 12952 32978
rect 12900 32914 12952 32920
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 13004 32201 13032 34020
rect 13320 34031 13322 34040
rect 13268 34002 13320 34008
rect 13084 33992 13136 33998
rect 13084 33934 13136 33940
rect 13096 33658 13124 33934
rect 13174 33688 13230 33697
rect 13084 33652 13136 33658
rect 13174 33623 13176 33632
rect 13084 33594 13136 33600
rect 13228 33623 13230 33632
rect 13176 33594 13228 33600
rect 13266 33416 13322 33425
rect 13266 33351 13322 33360
rect 13280 32978 13308 33351
rect 13360 33312 13412 33318
rect 13360 33254 13412 33260
rect 13372 33114 13400 33254
rect 13360 33108 13412 33114
rect 13360 33050 13412 33056
rect 13268 32972 13320 32978
rect 13268 32914 13320 32920
rect 12990 32192 13046 32201
rect 12990 32127 13046 32136
rect 13004 31958 13032 32127
rect 12992 31952 13044 31958
rect 12992 31894 13044 31900
rect 12636 31726 12940 31754
rect 12440 31136 12492 31142
rect 12360 31096 12440 31124
rect 12440 31078 12492 31084
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11886 29880 11942 29889
rect 11886 29815 11888 29824
rect 11940 29815 11942 29824
rect 11888 29786 11940 29792
rect 11886 29744 11942 29753
rect 11886 29679 11942 29688
rect 11900 29646 11928 29679
rect 11992 29646 12020 30194
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 11992 29481 12020 29582
rect 11978 29472 12034 29481
rect 12084 29458 12112 30602
rect 12176 30394 12204 30670
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12164 30388 12216 30394
rect 12164 30330 12216 30336
rect 12268 30376 12296 30602
rect 12348 30388 12400 30394
rect 12268 30348 12348 30376
rect 12268 30274 12296 30348
rect 12348 30330 12400 30336
rect 12176 30246 12296 30274
rect 12176 29578 12204 30246
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12268 29714 12296 29990
rect 12452 29850 12480 30126
rect 12532 30116 12584 30122
rect 12532 30058 12584 30064
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12164 29572 12216 29578
rect 12164 29514 12216 29520
rect 12348 29572 12400 29578
rect 12544 29560 12572 30058
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12400 29532 12572 29560
rect 12348 29514 12400 29520
rect 12084 29430 12287 29458
rect 11978 29407 12034 29416
rect 12164 29300 12216 29306
rect 12259 29288 12287 29430
rect 12544 29306 12572 29532
rect 12636 29306 12664 29990
rect 12728 29714 12756 30670
rect 12808 29776 12860 29782
rect 12808 29718 12860 29724
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12716 29504 12768 29510
rect 12714 29472 12716 29481
rect 12768 29472 12770 29481
rect 12714 29407 12770 29416
rect 12532 29300 12584 29306
rect 12259 29260 12296 29288
rect 12164 29242 12216 29248
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 11992 28762 12020 29106
rect 12072 28960 12124 28966
rect 12072 28902 12124 28908
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 11716 28478 11836 28506
rect 11888 28484 11940 28490
rect 11612 28416 11664 28422
rect 11612 28358 11664 28364
rect 11624 27946 11652 28358
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11532 27798 11652 27826
rect 11440 27390 11560 27418
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11428 27328 11480 27334
rect 11428 27270 11480 27276
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 11242 27024 11298 27033
rect 11152 26988 11204 26994
rect 11242 26959 11298 26968
rect 11152 26930 11204 26936
rect 11256 26586 11284 26959
rect 11348 26926 11376 27270
rect 11440 27062 11468 27270
rect 11532 27130 11560 27390
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11428 27056 11480 27062
rect 11428 26998 11480 27004
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 10876 26444 10928 26450
rect 10980 26438 11100 26466
rect 10876 26386 10928 26392
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10980 25974 11008 26318
rect 11072 26246 11100 26438
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11060 26240 11112 26246
rect 11060 26182 11112 26188
rect 11058 26072 11114 26081
rect 11058 26007 11114 26016
rect 11072 25974 11100 26007
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 11060 25968 11112 25974
rect 11164 25945 11192 26386
rect 11060 25910 11112 25916
rect 11150 25936 11206 25945
rect 10876 25900 10928 25906
rect 11150 25871 11206 25880
rect 10876 25842 10928 25848
rect 10888 25129 10916 25842
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11072 25294 11100 25638
rect 11060 25288 11112 25294
rect 11152 25288 11204 25294
rect 11060 25230 11112 25236
rect 11150 25256 11152 25265
rect 11204 25256 11206 25265
rect 10968 25220 11020 25226
rect 11150 25191 11206 25200
rect 10968 25162 11020 25168
rect 10874 25120 10930 25129
rect 10874 25055 10930 25064
rect 10980 24954 11008 25162
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11164 24834 11192 25094
rect 11256 24954 11284 26386
rect 11348 25770 11376 26862
rect 11532 26450 11560 27066
rect 11624 26926 11652 27798
rect 11716 27554 11744 28478
rect 11888 28426 11940 28432
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11808 27674 11836 28358
rect 11900 28150 11928 28426
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 12084 28014 12112 28902
rect 12176 28626 12204 29242
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 12176 27606 12204 27814
rect 12164 27600 12216 27606
rect 11716 27526 11836 27554
rect 12164 27542 12216 27548
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11612 26920 11664 26926
rect 11612 26862 11664 26868
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11426 26072 11482 26081
rect 11716 26058 11744 26930
rect 11808 26382 11836 27526
rect 11978 27024 12034 27033
rect 11978 26959 11980 26968
rect 12032 26959 12034 26968
rect 12164 26988 12216 26994
rect 11980 26930 12032 26936
rect 12164 26930 12216 26936
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11624 26042 11744 26058
rect 11426 26007 11482 26016
rect 11612 26036 11744 26042
rect 11336 25764 11388 25770
rect 11336 25706 11388 25712
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 10980 24818 11192 24834
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10968 24812 11192 24818
rect 11020 24806 11192 24812
rect 10968 24754 11020 24760
rect 10888 24698 10916 24754
rect 11152 24744 11204 24750
rect 10888 24670 11100 24698
rect 11152 24686 11204 24692
rect 11072 24206 11100 24670
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10876 23588 10928 23594
rect 10876 23530 10928 23536
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10612 23338 10640 23462
rect 10612 23310 10732 23338
rect 10888 23322 10916 23530
rect 10704 23254 10732 23310
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10692 23248 10744 23254
rect 10598 23216 10654 23225
rect 10692 23190 10744 23196
rect 10598 23151 10654 23160
rect 10612 23118 10640 23151
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10598 22944 10654 22953
rect 10598 22879 10654 22888
rect 10612 22506 10640 22879
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10600 22092 10652 22098
rect 10520 22052 10600 22080
rect 10520 22001 10548 22052
rect 10600 22034 10652 22040
rect 10506 21992 10562 22001
rect 10506 21927 10562 21936
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10428 21350 10456 21830
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10244 20992 10272 21082
rect 10324 21004 10376 21010
rect 10244 20964 10324 20992
rect 10324 20946 10376 20952
rect 10048 20936 10100 20942
rect 10046 20904 10048 20913
rect 10100 20904 10102 20913
rect 10046 20839 10102 20848
rect 10232 20868 10284 20874
rect 10428 20856 10456 21082
rect 10284 20828 10456 20856
rect 10232 20810 10284 20816
rect 10520 20714 10548 21830
rect 10612 21690 10640 21898
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10612 21418 10640 21626
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10520 20686 10640 20714
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10322 20496 10378 20505
rect 10322 20431 10378 20440
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10152 19446 10180 19654
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10060 18970 10088 19246
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9876 18584 9996 18612
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9600 18193 9628 18226
rect 9586 18184 9642 18193
rect 9220 18148 9272 18154
rect 9586 18119 9642 18128
rect 9220 18090 9272 18096
rect 9036 18080 9088 18086
rect 9128 18080 9180 18086
rect 9036 18022 9088 18028
rect 9126 18048 9128 18057
rect 9180 18048 9182 18057
rect 9048 17814 9076 18022
rect 9126 17983 9182 17992
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9048 16794 9076 17750
rect 9140 17678 9168 17983
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9232 15570 9260 18090
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9416 17202 9444 17478
rect 9784 17202 9812 17478
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9416 16590 9444 17138
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9692 16250 9720 17138
rect 9876 16250 9904 18584
rect 9956 18420 10008 18426
rect 10152 18408 10180 19246
rect 10244 18766 10272 20198
rect 10336 19718 10364 20431
rect 10428 20097 10456 20538
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10414 20088 10470 20097
rect 10414 20023 10470 20032
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10336 19378 10364 19654
rect 10428 19394 10456 19790
rect 10520 19514 10548 20470
rect 10612 20398 10640 20686
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10704 20233 10732 23190
rect 10784 22976 10836 22982
rect 10980 22964 11008 24142
rect 11072 23905 11100 24142
rect 11058 23896 11114 23905
rect 11058 23831 11114 23840
rect 11164 23202 11192 24686
rect 11256 24290 11284 24890
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11348 24410 11376 24754
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 11256 24262 11376 24290
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11256 23730 11284 24142
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11348 23322 11376 24262
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11164 23174 11376 23202
rect 11440 23186 11468 26007
rect 11664 26030 11744 26036
rect 11612 25978 11664 25984
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11532 25498 11560 25910
rect 12176 25838 12204 26930
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 11980 25696 12032 25702
rect 11886 25664 11942 25673
rect 11808 25622 11886 25650
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11518 25392 11574 25401
rect 11518 25327 11574 25336
rect 11532 25294 11560 25327
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11060 23112 11112 23118
rect 11058 23080 11060 23089
rect 11244 23112 11296 23118
rect 11112 23080 11114 23089
rect 11244 23054 11296 23060
rect 11058 23015 11114 23024
rect 10836 22936 11008 22964
rect 10784 22918 10836 22924
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10782 22672 10838 22681
rect 10782 22607 10784 22616
rect 10836 22607 10838 22616
rect 10784 22578 10836 22584
rect 10888 22545 10916 22714
rect 10980 22574 11008 22936
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 11072 22778 11100 22918
rect 11256 22817 11284 23054
rect 11242 22808 11298 22817
rect 11060 22772 11112 22778
rect 11242 22743 11298 22752
rect 11060 22714 11112 22720
rect 10968 22568 11020 22574
rect 10874 22536 10930 22545
rect 10968 22510 11020 22516
rect 10874 22471 10930 22480
rect 10782 22400 10838 22409
rect 10782 22335 10838 22344
rect 10796 21622 10824 22335
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10796 21146 10824 21558
rect 10888 21554 10916 22471
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10980 20924 11008 22102
rect 11072 21554 11100 22714
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11164 22234 11192 22578
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11164 21690 11192 22170
rect 11256 22098 11284 22646
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11058 21448 11114 21457
rect 11348 21400 11376 23174
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11426 22400 11482 22409
rect 11426 22335 11482 22344
rect 11440 22030 11468 22335
rect 11532 22234 11560 25230
rect 11624 24410 11652 25230
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11716 24818 11744 24890
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11702 24440 11758 24449
rect 11612 24404 11664 24410
rect 11702 24375 11758 24384
rect 11612 24346 11664 24352
rect 11612 24200 11664 24206
rect 11716 24188 11744 24375
rect 11664 24160 11744 24188
rect 11612 24142 11664 24148
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11624 23118 11652 23462
rect 11612 23112 11664 23118
rect 11610 23080 11612 23089
rect 11664 23080 11666 23089
rect 11610 23015 11666 23024
rect 11612 22568 11664 22574
rect 11610 22536 11612 22545
rect 11664 22536 11666 22545
rect 11610 22471 11666 22480
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11426 21856 11482 21865
rect 11426 21791 11482 21800
rect 11440 21690 11468 21791
rect 11532 21690 11560 21898
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11532 21593 11560 21626
rect 11518 21584 11574 21593
rect 11518 21519 11574 21528
rect 11058 21383 11114 21392
rect 11072 20942 11100 21383
rect 11256 21372 11376 21400
rect 11150 21176 11206 21185
rect 11150 21111 11206 21120
rect 11164 21078 11192 21111
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 10893 20896 11008 20924
rect 11060 20936 11112 20942
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10796 20777 10824 20810
rect 10893 20788 10921 20896
rect 11060 20878 11112 20884
rect 10782 20768 10838 20777
rect 10782 20703 10838 20712
rect 10888 20760 10921 20788
rect 10968 20800 11020 20806
rect 10888 20618 10916 20760
rect 11060 20800 11112 20806
rect 10968 20742 11020 20748
rect 11058 20768 11060 20777
rect 11112 20768 11114 20777
rect 10796 20590 10916 20618
rect 10796 20466 10824 20590
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10690 20224 10746 20233
rect 10690 20159 10746 20168
rect 10796 19854 10824 20402
rect 10888 20369 10916 20402
rect 10980 20398 11008 20742
rect 11058 20703 11114 20712
rect 10968 20392 11020 20398
rect 10874 20360 10930 20369
rect 11152 20392 11204 20398
rect 10968 20334 11020 20340
rect 11072 20352 11152 20380
rect 10874 20295 10930 20304
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10888 20097 10916 20198
rect 10874 20088 10930 20097
rect 10874 20023 10930 20032
rect 10980 19990 11008 20334
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19514 10732 19722
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10324 19372 10376 19378
rect 10428 19366 10640 19394
rect 10324 19314 10376 19320
rect 10336 18766 10364 19314
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10324 18760 10376 18766
rect 10520 18737 10548 19178
rect 10324 18702 10376 18708
rect 10506 18728 10562 18737
rect 10416 18692 10468 18698
rect 10506 18663 10508 18672
rect 10416 18634 10468 18640
rect 10560 18663 10562 18672
rect 10508 18634 10560 18640
rect 10008 18380 10180 18408
rect 9956 18362 10008 18368
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 9416 15366 9444 15846
rect 9968 15570 9996 18226
rect 10060 16250 10088 18380
rect 10428 18290 10456 18634
rect 10416 18284 10468 18290
rect 10336 18244 10416 18272
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10244 17814 10272 18022
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10336 17678 10364 18244
rect 10416 18226 10468 18232
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10428 17678 10456 18090
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10244 17270 10272 17614
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10336 16726 10364 17614
rect 10520 17610 10548 18634
rect 10612 18358 10640 19366
rect 10874 19000 10930 19009
rect 10874 18935 10930 18944
rect 10782 18864 10838 18873
rect 10782 18799 10838 18808
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10520 17338 10548 17546
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10796 17202 10824 18799
rect 10888 18766 10916 18935
rect 10980 18834 11008 19926
rect 11072 19145 11100 20352
rect 11152 20334 11204 20340
rect 11152 20256 11204 20262
rect 11150 20224 11152 20233
rect 11204 20224 11206 20233
rect 11150 20159 11206 20168
rect 11256 19922 11284 21372
rect 11334 21312 11390 21321
rect 11334 21247 11390 21256
rect 11348 19961 11376 21247
rect 11624 21026 11652 22374
rect 11532 20998 11652 21026
rect 11532 20890 11560 20998
rect 11440 20862 11560 20890
rect 11334 19952 11390 19961
rect 11244 19916 11296 19922
rect 11334 19887 11390 19896
rect 11244 19858 11296 19864
rect 11348 19514 11376 19887
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11058 19136 11114 19145
rect 11058 19071 11114 19080
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18426 11008 18566
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11164 18358 11192 18634
rect 11440 18578 11468 20862
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11532 20466 11560 20742
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11532 19854 11560 20402
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11532 18902 11560 19246
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11348 18550 11468 18578
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10888 17746 10916 18090
rect 10966 17912 11022 17921
rect 10966 17847 11022 17856
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17338 10916 17546
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10704 16590 10732 16934
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10796 16250 10824 16662
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 14074 8156 14214
rect 8220 14074 8248 14962
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7852 13394 7880 13738
rect 8496 13530 8524 14554
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 9416 10062 9444 15302
rect 9784 14550 9812 15506
rect 9968 15162 9996 15506
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10060 14618 10088 16186
rect 10796 15162 10824 16186
rect 10980 16114 11008 17847
rect 11348 17338 11376 18550
rect 11624 18442 11652 20742
rect 11716 19922 11744 24160
rect 11808 23730 11836 25622
rect 12268 25684 12296 29260
rect 12532 29242 12584 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 12544 29102 12572 29242
rect 12820 29170 12848 29718
rect 12912 29458 12940 31726
rect 12992 30796 13044 30802
rect 12992 30738 13044 30744
rect 13004 30394 13032 30738
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 13084 30116 13136 30122
rect 13084 30058 13136 30064
rect 12990 29880 13046 29889
rect 12990 29815 13046 29824
rect 13004 29646 13032 29815
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 13096 29492 13124 30058
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 13176 29640 13228 29646
rect 13174 29608 13176 29617
rect 13228 29608 13230 29617
rect 13174 29543 13230 29552
rect 13096 29464 13216 29492
rect 12912 29430 13032 29458
rect 12900 29232 12952 29238
rect 12900 29174 12952 29180
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12348 28960 12400 28966
rect 12532 28960 12584 28966
rect 12400 28920 12480 28948
rect 12348 28902 12400 28908
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12360 27946 12388 28698
rect 12452 27946 12480 28920
rect 12532 28902 12584 28908
rect 12544 28490 12572 28902
rect 12820 28778 12848 29106
rect 12728 28762 12848 28778
rect 12716 28756 12848 28762
rect 12768 28750 12848 28756
rect 12716 28698 12768 28704
rect 12624 28620 12676 28626
rect 12676 28580 12756 28608
rect 12624 28562 12676 28568
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12348 27940 12400 27946
rect 12348 27882 12400 27888
rect 12440 27940 12492 27946
rect 12440 27882 12492 27888
rect 12348 27668 12400 27674
rect 12348 27610 12400 27616
rect 12360 26314 12388 27610
rect 12624 27464 12676 27470
rect 12622 27432 12624 27441
rect 12676 27432 12678 27441
rect 12622 27367 12678 27376
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12348 26308 12400 26314
rect 12348 26250 12400 26256
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 12452 26042 12480 26250
rect 12440 26036 12492 26042
rect 11980 25638 12032 25644
rect 12176 25656 12296 25684
rect 12360 25996 12440 26024
rect 11886 25599 11942 25608
rect 11992 25498 12020 25638
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11992 25294 12020 25434
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11886 24984 11942 24993
rect 11886 24919 11942 24928
rect 12072 24948 12124 24954
rect 11900 24818 11928 24919
rect 12072 24890 12124 24896
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11900 24274 11928 24550
rect 11992 24410 12020 24754
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 11900 23730 11928 24210
rect 11992 23798 12020 24346
rect 12084 24138 12112 24890
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 12084 23633 12112 24074
rect 12070 23624 12126 23633
rect 12070 23559 12126 23568
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11808 22098 11836 22374
rect 11900 22273 11928 23190
rect 12176 23066 12204 25656
rect 12254 25120 12310 25129
rect 12254 25055 12310 25064
rect 12268 24818 12296 25055
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12254 23896 12310 23905
rect 12254 23831 12310 23840
rect 12268 23594 12296 23831
rect 12256 23588 12308 23594
rect 12256 23530 12308 23536
rect 11992 23050 12296 23066
rect 11992 23044 12308 23050
rect 11992 23038 12256 23044
rect 11992 22681 12020 23038
rect 12256 22986 12308 22992
rect 12072 22976 12124 22982
rect 12360 22930 12388 25996
rect 12440 25978 12492 25984
rect 12544 25770 12572 26318
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 12544 25294 12572 25706
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12544 23508 12572 25230
rect 12636 24954 12664 26862
rect 12728 25820 12756 28580
rect 12912 27690 12940 29174
rect 13004 28966 13032 29430
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 13096 29209 13124 29242
rect 13082 29200 13138 29209
rect 13082 29135 13138 29144
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 13004 28218 13032 28358
rect 13096 28218 13124 29135
rect 13188 29073 13216 29464
rect 13268 29096 13320 29102
rect 13174 29064 13230 29073
rect 13268 29038 13320 29044
rect 13372 29050 13400 29650
rect 13464 29170 13492 34360
rect 13556 34202 13584 36858
rect 13636 36644 13688 36650
rect 13636 36586 13688 36592
rect 13648 35086 13676 36586
rect 13832 36174 13860 38286
rect 14096 37664 14148 37670
rect 14096 37606 14148 37612
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 13912 37392 13964 37398
rect 13912 37334 13964 37340
rect 13924 36854 13952 37334
rect 13912 36848 13964 36854
rect 13912 36790 13964 36796
rect 13912 36576 13964 36582
rect 13912 36518 13964 36524
rect 13924 36378 13952 36518
rect 13912 36372 13964 36378
rect 13912 36314 13964 36320
rect 13820 36168 13872 36174
rect 13820 36110 13872 36116
rect 13728 36100 13780 36106
rect 13728 36042 13780 36048
rect 13740 35834 13768 36042
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13832 35834 13860 35974
rect 14016 35850 14044 37402
rect 14108 36786 14136 37606
rect 14200 37330 14228 38354
rect 14292 37466 14320 38830
rect 14372 38276 14424 38282
rect 14372 38218 14424 38224
rect 14280 37460 14332 37466
rect 14280 37402 14332 37408
rect 14188 37324 14240 37330
rect 14188 37266 14240 37272
rect 14292 36825 14320 37402
rect 14278 36816 14334 36825
rect 14096 36780 14148 36786
rect 14278 36751 14334 36760
rect 14096 36722 14148 36728
rect 14292 36122 14320 36751
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 13820 35828 13872 35834
rect 13820 35770 13872 35776
rect 13924 35822 14044 35850
rect 14200 36094 14320 36122
rect 13820 35556 13872 35562
rect 13820 35498 13872 35504
rect 13636 35080 13688 35086
rect 13636 35022 13688 35028
rect 13832 34610 13860 35498
rect 13924 35086 13952 35822
rect 14004 35692 14056 35698
rect 14004 35634 14056 35640
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 13912 34740 13964 34746
rect 13912 34682 13964 34688
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13924 34066 13952 34682
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13556 32502 13584 33934
rect 13820 33856 13872 33862
rect 13820 33798 13872 33804
rect 13636 33516 13688 33522
rect 13636 33458 13688 33464
rect 13648 33289 13676 33458
rect 13728 33312 13780 33318
rect 13634 33280 13690 33289
rect 13728 33254 13780 33260
rect 13634 33215 13690 33224
rect 13634 33144 13690 33153
rect 13740 33130 13768 33254
rect 13690 33102 13768 33130
rect 13634 33079 13636 33088
rect 13688 33079 13690 33088
rect 13636 33050 13688 33056
rect 13634 32600 13690 32609
rect 13634 32535 13636 32544
rect 13688 32535 13690 32544
rect 13636 32506 13688 32512
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13542 32328 13598 32337
rect 13542 32263 13598 32272
rect 13556 31958 13584 32263
rect 13728 32224 13780 32230
rect 13728 32166 13780 32172
rect 13544 31952 13596 31958
rect 13544 31894 13596 31900
rect 13740 31686 13768 32166
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13556 31482 13584 31622
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13634 31376 13690 31385
rect 13634 31311 13690 31320
rect 13728 31340 13780 31346
rect 13648 30870 13676 31311
rect 13728 31282 13780 31288
rect 13740 30938 13768 31282
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13636 30864 13688 30870
rect 13636 30806 13688 30812
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13542 29744 13598 29753
rect 13542 29679 13598 29688
rect 13556 29510 13584 29679
rect 13740 29617 13768 30534
rect 13726 29608 13782 29617
rect 13726 29543 13782 29552
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13648 29050 13676 29106
rect 13174 28999 13230 29008
rect 13280 28762 13308 29038
rect 13372 29022 13676 29050
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13268 28756 13320 28762
rect 13268 28698 13320 28704
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13372 28642 13400 28698
rect 13280 28614 13400 28642
rect 13464 28626 13492 28902
rect 13452 28620 13504 28626
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 12820 27662 12940 27690
rect 12820 27606 12848 27662
rect 12808 27600 12860 27606
rect 12808 27542 12860 27548
rect 12900 27600 12952 27606
rect 13004 27588 13032 27950
rect 13096 27713 13124 28018
rect 13082 27704 13138 27713
rect 13188 27674 13216 28154
rect 13082 27639 13138 27648
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 12952 27560 13032 27588
rect 12900 27542 12952 27548
rect 12820 27130 12848 27542
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12912 26994 12940 27542
rect 13280 27470 13308 28614
rect 13452 28562 13504 28568
rect 13452 28484 13504 28490
rect 13556 28472 13584 28902
rect 13504 28444 13584 28472
rect 13452 28426 13504 28432
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13188 27130 13216 27406
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 12900 26988 12952 26994
rect 12900 26930 12952 26936
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 12808 25832 12860 25838
rect 12728 25792 12808 25820
rect 12808 25774 12860 25780
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12820 24614 12848 25774
rect 12912 25362 12940 26930
rect 13004 26586 13032 26930
rect 13280 26738 13308 27270
rect 13096 26710 13308 26738
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 12990 25392 13046 25401
rect 12900 25356 12952 25362
rect 12990 25327 13046 25336
rect 12900 25298 12952 25304
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12714 24304 12770 24313
rect 12714 24239 12716 24248
rect 12768 24239 12770 24248
rect 12716 24210 12768 24216
rect 12912 24206 12940 25094
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12622 23760 12678 23769
rect 13004 23730 13032 25327
rect 13096 23866 13124 26710
rect 13266 25800 13322 25809
rect 13266 25735 13268 25744
rect 13320 25735 13322 25744
rect 13268 25706 13320 25712
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 12622 23695 12624 23704
rect 12676 23695 12678 23704
rect 12992 23724 13044 23730
rect 12624 23666 12676 23672
rect 12992 23666 13044 23672
rect 12624 23520 12676 23526
rect 12544 23480 12624 23508
rect 12624 23462 12676 23468
rect 12636 23118 12664 23462
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12072 22918 12124 22924
rect 11978 22672 12034 22681
rect 11978 22607 12034 22616
rect 11886 22264 11942 22273
rect 11886 22199 11942 22208
rect 11900 22148 11928 22199
rect 11980 22160 12032 22166
rect 11900 22120 11980 22148
rect 11980 22102 12032 22108
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 18970 11744 19314
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11440 18414 11652 18442
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11440 16590 11468 18414
rect 11716 18222 11744 18702
rect 11808 18630 11836 21898
rect 11900 21690 11928 21966
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11900 21554 11928 21626
rect 12084 21554 12112 22918
rect 12268 22902 12388 22930
rect 12268 21894 12296 22902
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12360 22506 12388 22714
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12360 22098 12388 22170
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12452 22030 12480 23054
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12544 22545 12572 22918
rect 12820 22710 12848 22986
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 12716 22568 12768 22574
rect 12530 22536 12586 22545
rect 12716 22510 12768 22516
rect 12530 22471 12586 22480
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 21418 12112 21490
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11900 20233 11928 20538
rect 11886 20224 11942 20233
rect 11886 20159 11942 20168
rect 11992 19990 12020 21354
rect 12268 21146 12296 21830
rect 12452 21350 12480 21966
rect 12624 21888 12676 21894
rect 12544 21848 12624 21876
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12544 21162 12572 21848
rect 12624 21830 12676 21836
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12452 21134 12572 21162
rect 12636 21146 12664 21490
rect 12728 21418 12756 22510
rect 12820 21622 12848 22646
rect 12912 22522 12940 22986
rect 12912 22494 13032 22522
rect 13096 22506 13124 23054
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12900 21480 12952 21486
rect 12898 21448 12900 21457
rect 12952 21448 12954 21457
rect 12716 21412 12768 21418
rect 12898 21383 12954 21392
rect 12716 21354 12768 21360
rect 12624 21140 12676 21146
rect 12070 21040 12126 21049
rect 12070 20975 12126 20984
rect 12084 20806 12112 20975
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12176 20618 12204 20742
rect 12084 20590 12204 20618
rect 12084 20466 12112 20590
rect 12162 20496 12218 20505
rect 12072 20460 12124 20466
rect 12162 20431 12218 20440
rect 12072 20402 12124 20408
rect 12176 20398 12204 20431
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12072 20256 12124 20262
rect 12124 20204 12204 20210
rect 12072 20198 12204 20204
rect 12084 20182 12204 20198
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11520 18148 11572 18154
rect 11520 18090 11572 18096
rect 11532 17746 11560 18090
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11624 17746 11652 18022
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11532 16794 11560 17070
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11072 15366 11100 16390
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 15706 11376 15846
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11532 15434 11560 16730
rect 11716 16697 11744 17274
rect 11808 16998 11836 18226
rect 11900 17678 11928 19858
rect 12070 19680 12126 19689
rect 12070 19615 12126 19624
rect 12084 19446 12112 19615
rect 12176 19446 12204 20182
rect 12072 19440 12124 19446
rect 11978 19408 12034 19417
rect 12072 19382 12124 19388
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11978 19343 11980 19352
rect 12032 19343 12034 19352
rect 11980 19314 12032 19320
rect 12176 19122 12204 19382
rect 12268 19378 12296 21082
rect 12452 21049 12480 21134
rect 12624 21082 12676 21088
rect 12438 21040 12494 21049
rect 12438 20975 12494 20984
rect 12636 20942 12664 21082
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12728 20806 12756 21354
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12346 20088 12402 20097
rect 12346 20023 12402 20032
rect 12360 19922 12388 20023
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 12360 19514 12388 19722
rect 12544 19514 12572 20198
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19514 12664 19790
rect 12728 19514 12756 20742
rect 12820 19718 12848 21286
rect 13004 21162 13032 22494
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 13096 21690 13124 22442
rect 13188 22166 13216 24754
rect 13266 24440 13322 24449
rect 13266 24375 13322 24384
rect 13280 23730 13308 24375
rect 13372 24342 13400 28154
rect 13464 26042 13492 28426
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13556 27878 13584 28018
rect 13648 27946 13676 29022
rect 13740 28558 13768 29038
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13832 28218 13860 33798
rect 14016 33658 14044 35634
rect 14200 35562 14228 36094
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 14188 35556 14240 35562
rect 14188 35498 14240 35504
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 14108 34746 14136 34886
rect 14096 34740 14148 34746
rect 14096 34682 14148 34688
rect 14200 34678 14228 34886
rect 14188 34672 14240 34678
rect 14188 34614 14240 34620
rect 14096 34604 14148 34610
rect 14096 34546 14148 34552
rect 14108 33998 14136 34546
rect 14292 34542 14320 35974
rect 14384 35290 14412 38218
rect 14660 37942 14688 38898
rect 14648 37936 14700 37942
rect 14648 37878 14700 37884
rect 14464 37732 14516 37738
rect 14464 37674 14516 37680
rect 14476 37466 14504 37674
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 14372 35284 14424 35290
rect 14372 35226 14424 35232
rect 14476 34678 14504 37402
rect 14660 37330 14688 37878
rect 14648 37324 14700 37330
rect 14648 37266 14700 37272
rect 14556 37188 14608 37194
rect 14556 37130 14608 37136
rect 14568 36922 14596 37130
rect 14556 36916 14608 36922
rect 14556 36858 14608 36864
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14464 34672 14516 34678
rect 14464 34614 14516 34620
rect 14568 34542 14596 36654
rect 14660 35766 14688 37266
rect 14752 36242 14780 39986
rect 15016 39840 15068 39846
rect 15016 39782 15068 39788
rect 15028 39030 15056 39782
rect 15016 39024 15068 39030
rect 15016 38966 15068 38972
rect 15120 38554 15148 40462
rect 15752 40384 15804 40390
rect 15752 40326 15804 40332
rect 15292 39976 15344 39982
rect 15292 39918 15344 39924
rect 15108 38548 15160 38554
rect 15108 38490 15160 38496
rect 14832 38276 14884 38282
rect 14832 38218 14884 38224
rect 14844 37126 14872 38218
rect 15304 38214 15332 39918
rect 15568 39840 15620 39846
rect 15568 39782 15620 39788
rect 15476 38412 15528 38418
rect 15476 38354 15528 38360
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 15292 38208 15344 38214
rect 15292 38150 15344 38156
rect 15120 37942 15148 38150
rect 15108 37936 15160 37942
rect 15108 37878 15160 37884
rect 14924 37868 14976 37874
rect 14924 37810 14976 37816
rect 14936 37777 14964 37810
rect 14922 37768 14978 37777
rect 14922 37703 14978 37712
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 14936 37262 14964 37606
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 14922 36816 14978 36825
rect 14922 36751 14978 36760
rect 14936 36718 14964 36751
rect 14924 36712 14976 36718
rect 14924 36654 14976 36660
rect 14936 36582 14964 36654
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 14740 36236 14792 36242
rect 14740 36178 14792 36184
rect 14752 36145 14780 36178
rect 14738 36136 14794 36145
rect 14738 36071 14794 36080
rect 14648 35760 14700 35766
rect 14648 35702 14700 35708
rect 14660 35086 14688 35702
rect 14832 35692 14884 35698
rect 14832 35634 14884 35640
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14568 33998 14596 34478
rect 14844 34066 14872 35634
rect 14924 35012 14976 35018
rect 14924 34954 14976 34960
rect 14936 34746 14964 34954
rect 15014 34776 15070 34785
rect 14924 34740 14976 34746
rect 15070 34746 15148 34762
rect 15070 34740 15160 34746
rect 15070 34734 15108 34740
rect 15014 34711 15070 34720
rect 14924 34682 14976 34688
rect 15108 34682 15160 34688
rect 15108 34468 15160 34474
rect 15108 34410 15160 34416
rect 14922 34232 14978 34241
rect 14922 34167 14978 34176
rect 14832 34060 14884 34066
rect 14832 34002 14884 34008
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 14556 33992 14608 33998
rect 14608 33952 14688 33980
rect 14556 33934 14608 33940
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 14464 33584 14516 33590
rect 14464 33526 14516 33532
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 13924 32434 13952 32846
rect 14002 32464 14058 32473
rect 13912 32428 13964 32434
rect 14002 32399 14004 32408
rect 13912 32370 13964 32376
rect 14056 32399 14058 32408
rect 14004 32370 14056 32376
rect 13924 30598 13952 32370
rect 14016 30598 14044 32370
rect 13912 30592 13964 30598
rect 13912 30534 13964 30540
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14016 30394 14044 30534
rect 14004 30388 14056 30394
rect 14004 30330 14056 30336
rect 14004 30048 14056 30054
rect 14004 29990 14056 29996
rect 14016 29850 14044 29990
rect 14004 29844 14056 29850
rect 14004 29786 14056 29792
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 13728 28144 13780 28150
rect 13728 28086 13780 28092
rect 13636 27940 13688 27946
rect 13636 27882 13688 27888
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13556 27690 13584 27814
rect 13556 27662 13676 27690
rect 13542 27568 13598 27577
rect 13542 27503 13598 27512
rect 13556 27130 13584 27503
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13648 26926 13676 27662
rect 13740 27606 13768 28086
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 13832 27713 13860 28018
rect 14016 27826 14044 29786
rect 14108 28506 14136 32846
rect 14200 32026 14228 33390
rect 14476 32434 14504 33526
rect 14660 33522 14688 33952
rect 14740 33924 14792 33930
rect 14740 33866 14792 33872
rect 14648 33516 14700 33522
rect 14648 33458 14700 33464
rect 14752 33386 14780 33866
rect 14936 33538 14964 34167
rect 15120 34134 15148 34410
rect 15212 34202 15240 37606
rect 15304 34626 15332 38150
rect 15384 37868 15436 37874
rect 15384 37810 15436 37816
rect 15396 37670 15424 37810
rect 15384 37664 15436 37670
rect 15384 37606 15436 37612
rect 15384 36100 15436 36106
rect 15384 36042 15436 36048
rect 15396 35290 15424 36042
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15488 34746 15516 38354
rect 15580 35306 15608 39782
rect 15764 39370 15792 40326
rect 15752 39364 15804 39370
rect 15752 39306 15804 39312
rect 15948 39098 15976 40462
rect 16488 40384 16540 40390
rect 16488 40326 16540 40332
rect 16500 40186 16528 40326
rect 16488 40180 16540 40186
rect 16488 40122 16540 40128
rect 16856 39976 16908 39982
rect 16856 39918 16908 39924
rect 16028 39296 16080 39302
rect 16028 39238 16080 39244
rect 16396 39296 16448 39302
rect 16396 39238 16448 39244
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 15660 38752 15712 38758
rect 15660 38694 15712 38700
rect 15844 38752 15896 38758
rect 15844 38694 15896 38700
rect 15672 36650 15700 38694
rect 15752 37800 15804 37806
rect 15752 37742 15804 37748
rect 15764 36786 15792 37742
rect 15856 37097 15884 38694
rect 15948 37874 15976 39034
rect 16040 38418 16068 39238
rect 16408 38758 16436 39238
rect 16396 38752 16448 38758
rect 16396 38694 16448 38700
rect 16868 38554 16896 39918
rect 17224 39840 17276 39846
rect 17224 39782 17276 39788
rect 17236 39438 17264 39782
rect 17132 39432 17184 39438
rect 17132 39374 17184 39380
rect 17224 39432 17276 39438
rect 17224 39374 17276 39380
rect 16856 38548 16908 38554
rect 16856 38490 16908 38496
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 16040 38010 16068 38354
rect 16856 38276 16908 38282
rect 16856 38218 16908 38224
rect 16028 38004 16080 38010
rect 16028 37946 16080 37952
rect 16212 38004 16264 38010
rect 16212 37946 16264 37952
rect 16224 37874 16252 37946
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 15842 37088 15898 37097
rect 15842 37023 15898 37032
rect 15856 36786 15884 37023
rect 15752 36780 15804 36786
rect 15752 36722 15804 36728
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 15660 36644 15712 36650
rect 15660 36586 15712 36592
rect 15672 36242 15700 36586
rect 15660 36236 15712 36242
rect 15660 36178 15712 36184
rect 15580 35278 15700 35306
rect 15568 35216 15620 35222
rect 15568 35158 15620 35164
rect 15476 34740 15528 34746
rect 15476 34682 15528 34688
rect 15304 34598 15516 34626
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 15382 34504 15438 34513
rect 15200 34196 15252 34202
rect 15200 34138 15252 34144
rect 15108 34128 15160 34134
rect 15108 34070 15160 34076
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 14844 33510 14964 33538
rect 14740 33380 14792 33386
rect 14740 33322 14792 33328
rect 14648 33312 14700 33318
rect 14648 33254 14700 33260
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14292 32026 14320 32370
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14384 31929 14412 32370
rect 14568 32065 14596 32370
rect 14554 32056 14610 32065
rect 14554 31991 14610 32000
rect 14370 31920 14426 31929
rect 14370 31855 14426 31864
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14188 31680 14240 31686
rect 14188 31622 14240 31628
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14200 30190 14228 31622
rect 14280 31272 14332 31278
rect 14280 31214 14332 31220
rect 14292 30394 14320 31214
rect 14476 30598 14504 31622
rect 14568 31142 14596 31826
rect 14556 31136 14608 31142
rect 14556 31078 14608 31084
rect 14568 30938 14596 31078
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14200 28762 14228 30126
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 14292 30025 14320 30058
rect 14278 30016 14334 30025
rect 14278 29951 14334 29960
rect 14292 29646 14320 29951
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14188 28756 14240 28762
rect 14188 28698 14240 28704
rect 14108 28478 14228 28506
rect 14384 28490 14412 30534
rect 14476 30433 14504 30534
rect 14462 30424 14518 30433
rect 14462 30359 14518 30368
rect 14462 29744 14518 29753
rect 14462 29679 14464 29688
rect 14516 29679 14518 29688
rect 14464 29650 14516 29656
rect 14568 28994 14596 30874
rect 14660 30569 14688 33254
rect 14844 32450 14872 33510
rect 14924 33448 14976 33454
rect 14924 33390 14976 33396
rect 14936 32570 14964 33390
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 14844 32422 14964 32450
rect 14740 32360 14792 32366
rect 14844 32337 14872 32422
rect 14740 32302 14792 32308
rect 14830 32328 14886 32337
rect 14752 31124 14780 32302
rect 14830 32263 14886 32272
rect 14832 31136 14884 31142
rect 14752 31096 14832 31124
rect 14832 31078 14884 31084
rect 14844 30870 14872 31078
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14936 30802 14964 32422
rect 15028 30938 15056 33934
rect 15120 33590 15148 33934
rect 15108 33584 15160 33590
rect 15108 33526 15160 33532
rect 15212 33522 15240 34138
rect 15304 33590 15332 34478
rect 15488 34474 15516 34598
rect 15382 34439 15438 34448
rect 15476 34468 15528 34474
rect 15396 33998 15424 34439
rect 15476 34410 15528 34416
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15292 33584 15344 33590
rect 15292 33526 15344 33532
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15580 33402 15608 35158
rect 15672 33522 15700 35278
rect 15764 35154 15792 36722
rect 15752 35148 15804 35154
rect 15752 35090 15804 35096
rect 15856 34610 15884 36722
rect 16224 36378 16252 37810
rect 16396 37800 16448 37806
rect 16868 37754 16896 38218
rect 17144 37874 17172 39374
rect 17040 37868 17092 37874
rect 17040 37810 17092 37816
rect 17132 37868 17184 37874
rect 17132 37810 17184 37816
rect 16396 37742 16448 37748
rect 16304 37120 16356 37126
rect 16304 37062 16356 37068
rect 16316 36718 16344 37062
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 16212 36372 16264 36378
rect 16212 36314 16264 36320
rect 16120 36168 16172 36174
rect 16120 36110 16172 36116
rect 16132 35494 16160 36110
rect 16212 36032 16264 36038
rect 16212 35974 16264 35980
rect 16224 35766 16252 35974
rect 16408 35834 16436 37742
rect 16776 37726 16896 37754
rect 16948 37800 17000 37806
rect 16948 37742 17000 37748
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16672 37664 16724 37670
rect 16672 37606 16724 37612
rect 16500 37330 16528 37606
rect 16488 37324 16540 37330
rect 16488 37266 16540 37272
rect 16488 37120 16540 37126
rect 16488 37062 16540 37068
rect 16500 36786 16528 37062
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16396 35828 16448 35834
rect 16396 35770 16448 35776
rect 16212 35760 16264 35766
rect 16212 35702 16264 35708
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 15844 34604 15896 34610
rect 15844 34546 15896 34552
rect 16028 34128 16080 34134
rect 16028 34070 16080 34076
rect 15844 34060 15896 34066
rect 15844 34002 15896 34008
rect 15660 33516 15712 33522
rect 15660 33458 15712 33464
rect 15672 33425 15700 33458
rect 15304 33374 15608 33402
rect 15658 33416 15714 33425
rect 15304 31754 15332 33374
rect 15658 33351 15714 33360
rect 15568 33312 15620 33318
rect 15382 33280 15438 33289
rect 15438 33238 15516 33266
rect 15568 33254 15620 33260
rect 15382 33215 15438 33224
rect 15382 32600 15438 32609
rect 15382 32535 15438 32544
rect 15212 31726 15332 31754
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 15108 30864 15160 30870
rect 15108 30806 15160 30812
rect 14924 30796 14976 30802
rect 14924 30738 14976 30744
rect 14646 30560 14702 30569
rect 14646 30495 14702 30504
rect 14832 30320 14884 30326
rect 14832 30262 14884 30268
rect 14844 29866 14872 30262
rect 15120 30258 15148 30806
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 15212 30190 15240 31726
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 14844 29838 14964 29866
rect 14648 29708 14700 29714
rect 14648 29650 14700 29656
rect 14832 29708 14884 29714
rect 14832 29650 14884 29656
rect 14660 29170 14688 29650
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14476 28966 14596 28994
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 13924 27798 14044 27826
rect 13818 27704 13874 27713
rect 13818 27639 13874 27648
rect 13728 27600 13780 27606
rect 13728 27542 13780 27548
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13740 26382 13768 27542
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13832 26382 13860 26726
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 13556 24818 13584 25162
rect 13648 24954 13676 25842
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13740 24993 13768 25230
rect 13726 24984 13782 24993
rect 13636 24948 13688 24954
rect 13726 24919 13782 24928
rect 13636 24890 13688 24896
rect 13726 24848 13782 24857
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13544 24812 13596 24818
rect 13726 24783 13728 24792
rect 13544 24754 13596 24760
rect 13780 24783 13782 24792
rect 13728 24754 13780 24760
rect 13464 24698 13492 24754
rect 13464 24670 13676 24698
rect 13464 24614 13492 24670
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13360 24336 13412 24342
rect 13412 24284 13584 24290
rect 13360 24278 13584 24284
rect 13372 24262 13584 24278
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 13464 23866 13492 24074
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13280 22778 13308 23054
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13372 22953 13400 22986
rect 13358 22944 13414 22953
rect 13358 22879 13414 22888
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 13372 22030 13400 22442
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13280 21690 13308 21966
rect 13464 21842 13492 22102
rect 13556 22030 13584 24262
rect 13648 23361 13676 24670
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13740 24206 13768 24346
rect 13832 24274 13860 25978
rect 13924 24818 13952 27798
rect 14108 27690 14136 28358
rect 14200 28218 14228 28478
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14200 28121 14228 28154
rect 14186 28112 14242 28121
rect 14186 28047 14242 28056
rect 14188 28008 14240 28014
rect 14188 27950 14240 27956
rect 14016 27662 14136 27690
rect 14016 27538 14044 27662
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 27305 14044 27474
rect 14002 27296 14058 27305
rect 14002 27231 14058 27240
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14016 26450 14044 26930
rect 14200 26772 14228 27950
rect 14372 27872 14424 27878
rect 14370 27840 14372 27849
rect 14424 27840 14426 27849
rect 14370 27775 14426 27784
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14292 26926 14320 27406
rect 14476 27282 14504 28966
rect 14660 28098 14688 29106
rect 14752 29034 14780 29106
rect 14844 29102 14872 29650
rect 14936 29646 14964 29838
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14936 29170 14964 29582
rect 14924 29164 14976 29170
rect 14924 29106 14976 29112
rect 14832 29096 14884 29102
rect 14832 29038 14884 29044
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14568 28070 14688 28098
rect 14568 27554 14596 28070
rect 14648 28008 14700 28014
rect 14752 27962 14780 28970
rect 15106 28928 15162 28937
rect 15106 28863 15162 28872
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14700 27956 14780 27962
rect 14648 27950 14780 27956
rect 14660 27934 14780 27950
rect 14568 27526 14688 27554
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14384 27254 14504 27282
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14200 26744 14320 26772
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14200 25294 14228 25842
rect 14292 25498 14320 26744
rect 14384 26450 14412 27254
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14384 26042 14412 26386
rect 14476 26330 14504 27066
rect 14568 26994 14596 27406
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14476 26314 14596 26330
rect 14476 26308 14608 26314
rect 14476 26302 14556 26308
rect 14556 26250 14608 26256
rect 14464 26240 14516 26246
rect 14464 26182 14516 26188
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14476 25702 14504 26182
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14280 25492 14332 25498
rect 14280 25434 14332 25440
rect 14372 25424 14424 25430
rect 14372 25366 14424 25372
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14004 25220 14056 25226
rect 14004 25162 14056 25168
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13910 24304 13966 24313
rect 13820 24268 13872 24274
rect 13910 24239 13966 24248
rect 13820 24210 13872 24216
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13634 23352 13690 23361
rect 13634 23287 13690 23296
rect 13832 22930 13860 24210
rect 13924 24206 13952 24239
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14016 23866 14044 25162
rect 14200 24886 14228 25230
rect 14292 24954 14320 25230
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14188 24880 14240 24886
rect 14188 24822 14240 24828
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 14094 24440 14150 24449
rect 14094 24375 14096 24384
rect 14148 24375 14150 24384
rect 14096 24346 14148 24352
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 14016 23050 14044 23462
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 13832 22902 14044 22930
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13464 21814 13584 21842
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13372 21185 13400 21626
rect 13556 21554 13584 21814
rect 13648 21729 13676 22510
rect 13740 22166 13768 22578
rect 13728 22160 13780 22166
rect 13728 22102 13780 22108
rect 13634 21720 13690 21729
rect 13634 21655 13690 21664
rect 13648 21622 13676 21655
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13358 21176 13414 21185
rect 13004 21134 13308 21162
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12900 20800 12952 20806
rect 12898 20768 12900 20777
rect 12952 20768 12954 20777
rect 12898 20703 12954 20712
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12912 20058 12940 20402
rect 13004 20233 13032 20878
rect 13096 20602 13124 20946
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13082 20496 13138 20505
rect 13188 20482 13216 20878
rect 13138 20454 13216 20482
rect 13082 20431 13138 20440
rect 13174 20360 13230 20369
rect 13280 20346 13308 21134
rect 13358 21111 13414 21120
rect 13280 20318 13400 20346
rect 13174 20295 13230 20304
rect 12990 20224 13046 20233
rect 12990 20159 13046 20168
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13004 19990 13032 20159
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 13004 19446 13032 19722
rect 13096 19718 13124 19790
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12256 19372 12308 19378
rect 13004 19334 13032 19382
rect 12256 19314 12308 19320
rect 12084 19094 12204 19122
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11992 18086 12020 18294
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12084 17338 12112 19094
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12176 18766 12204 18906
rect 12268 18766 12296 19314
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12912 19306 13032 19334
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12256 18760 12308 18766
rect 12636 18737 12664 19246
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18766 12756 19178
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12716 18760 12768 18766
rect 12256 18702 12308 18708
rect 12622 18728 12678 18737
rect 12716 18702 12768 18708
rect 12622 18663 12678 18672
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11702 16688 11758 16697
rect 12070 16688 12126 16697
rect 11992 16658 12070 16674
rect 11702 16623 11758 16632
rect 11980 16652 12070 16658
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11624 16250 11652 16526
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11716 16182 11744 16623
rect 12032 16646 12070 16652
rect 12070 16623 12126 16632
rect 12176 16640 12204 18566
rect 12544 18290 12572 18566
rect 12636 18358 12664 18663
rect 12820 18426 12848 19110
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12268 16794 12296 18158
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17338 12388 17478
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12544 17202 12572 18226
rect 12636 17785 12664 18294
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12622 17776 12678 17785
rect 12622 17711 12678 17720
rect 12728 17338 12756 18158
rect 12912 18086 12940 19306
rect 13096 18902 13124 19654
rect 13188 18902 13216 20295
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13280 19378 13308 20198
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12820 16658 12848 17682
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12912 17338 12940 17614
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12808 16652 12860 16658
rect 12176 16612 12296 16640
rect 11980 16594 12032 16600
rect 12072 16584 12124 16590
rect 12162 16552 12218 16561
rect 12124 16532 12162 16538
rect 12072 16526 12162 16532
rect 12084 16510 12162 16526
rect 12162 16487 12218 16496
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11992 16046 12020 16390
rect 12268 16114 12296 16612
rect 12808 16594 12860 16600
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10888 14822 10916 15302
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14618 10916 14758
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 10888 14074 10916 14554
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 11072 12434 11100 15302
rect 11532 15026 11560 15370
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14822 11836 14962
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11072 12406 11192 12434
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 11164 8974 11192 12406
rect 11992 11762 12020 15982
rect 12268 15502 12296 16050
rect 12820 15706 12848 16594
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12912 16250 12940 16390
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 13004 16046 13032 18362
rect 13280 18290 13308 18634
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17338 13124 18022
rect 13188 17921 13216 18158
rect 13174 17912 13230 17921
rect 13174 17847 13230 17856
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13188 17202 13216 17847
rect 13372 17746 13400 20318
rect 13556 19922 13584 21490
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13556 19825 13584 19858
rect 13542 19816 13598 19825
rect 13542 19751 13598 19760
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18290 13492 19178
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 18426 13584 18566
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13450 18184 13506 18193
rect 13450 18119 13452 18128
rect 13504 18119 13506 18128
rect 13452 18090 13504 18096
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13268 17536 13320 17542
rect 13320 17496 13400 17524
rect 13268 17478 13320 17484
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13280 16522 13308 17206
rect 13372 16726 13400 17496
rect 13464 17490 13492 17818
rect 13556 17814 13584 18022
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13648 17762 13676 21286
rect 13832 20942 13860 22714
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13924 22438 13952 22578
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13924 22001 13952 22170
rect 13910 21992 13966 22001
rect 13910 21927 13966 21936
rect 14016 21894 14044 22902
rect 14108 22030 14136 24210
rect 14200 24070 14228 24618
rect 14292 24585 14320 24686
rect 14278 24576 14334 24585
rect 14278 24511 14334 24520
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 20262 13860 20742
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13740 19009 13768 19178
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13726 19000 13782 19009
rect 13726 18935 13782 18944
rect 13832 18766 13860 19110
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13740 18154 13768 18566
rect 13832 18426 13860 18566
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13818 18320 13874 18329
rect 13818 18255 13874 18264
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13556 17678 13584 17750
rect 13648 17734 13768 17762
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13634 17640 13690 17649
rect 13634 17575 13636 17584
rect 13688 17575 13690 17584
rect 13636 17546 13688 17552
rect 13464 17462 13584 17490
rect 13450 17368 13506 17377
rect 13450 17303 13452 17312
rect 13504 17303 13506 17312
rect 13452 17274 13504 17280
rect 13556 17105 13584 17462
rect 13634 17232 13690 17241
rect 13634 17167 13690 17176
rect 13542 17096 13598 17105
rect 13542 17031 13598 17040
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15162 12572 15302
rect 13004 15162 13032 15982
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13188 15609 13216 15846
rect 13174 15600 13230 15609
rect 13174 15535 13176 15544
rect 13228 15535 13230 15544
rect 13176 15506 13228 15512
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13188 14550 13216 15506
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13372 14278 13400 16458
rect 13648 16454 13676 17167
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13740 15706 13768 17734
rect 13832 16998 13860 18255
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16794 13860 16934
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13924 16658 13952 21830
rect 14016 21554 14044 21830
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14004 21344 14056 21350
rect 14002 21312 14004 21321
rect 14056 21312 14058 21321
rect 14002 21247 14058 21256
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 19334 14044 20810
rect 14108 19961 14136 21966
rect 14200 21400 14228 23666
rect 14292 23662 14320 24511
rect 14384 24342 14412 25366
rect 14476 25294 14504 25638
rect 14660 25294 14688 27526
rect 14752 27402 14780 27934
rect 14740 27396 14792 27402
rect 14740 27338 14792 27344
rect 14752 26926 14780 27338
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14738 25664 14794 25673
rect 14738 25599 14794 25608
rect 14752 25498 14780 25599
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14660 24993 14688 25230
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14646 24984 14702 24993
rect 14646 24919 14702 24928
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14292 21554 14320 22170
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14200 21372 14320 21400
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14200 20398 14228 20810
rect 14292 20602 14320 21372
rect 14384 21350 14412 24278
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14476 20874 14504 24754
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14568 23798 14596 24074
rect 14752 23866 14780 25162
rect 14740 23860 14792 23866
rect 14660 23820 14740 23848
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14660 22642 14688 23820
rect 14740 23802 14792 23808
rect 14844 23798 14872 28698
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 15028 27878 15056 28154
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14844 23322 14872 23734
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14740 23248 14792 23254
rect 14936 23225 14964 27406
rect 15028 27305 15056 27542
rect 15014 27296 15070 27305
rect 15014 27231 15070 27240
rect 15120 27169 15148 28863
rect 15212 27946 15240 30126
rect 15396 28994 15424 32535
rect 15488 32280 15516 33238
rect 15580 32570 15608 33254
rect 15660 32904 15712 32910
rect 15712 32852 15792 32858
rect 15660 32846 15792 32852
rect 15672 32830 15792 32846
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15672 32570 15700 32710
rect 15568 32564 15620 32570
rect 15568 32506 15620 32512
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15488 32252 15608 32280
rect 15474 32192 15530 32201
rect 15474 32127 15530 32136
rect 15488 31890 15516 32127
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15476 31748 15528 31754
rect 15476 31690 15528 31696
rect 15488 31414 15516 31690
rect 15580 31686 15608 32252
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15672 31414 15700 32370
rect 15764 31822 15792 32830
rect 15752 31816 15804 31822
rect 15856 31793 15884 34002
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 15948 33658 15976 33934
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 16040 33402 16068 34070
rect 16132 33522 16160 35430
rect 16408 34746 16436 35770
rect 16580 35556 16632 35562
rect 16580 35498 16632 35504
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16396 34740 16448 34746
rect 16396 34682 16448 34688
rect 16224 33658 16252 34682
rect 16500 34610 16528 35022
rect 16592 34950 16620 35498
rect 16580 34944 16632 34950
rect 16580 34886 16632 34892
rect 16684 34678 16712 37606
rect 16776 35222 16804 37726
rect 16856 37188 16908 37194
rect 16856 37130 16908 37136
rect 16868 36854 16896 37130
rect 16856 36848 16908 36854
rect 16856 36790 16908 36796
rect 16856 36372 16908 36378
rect 16856 36314 16908 36320
rect 16764 35216 16816 35222
rect 16764 35158 16816 35164
rect 16672 34672 16724 34678
rect 16764 34672 16816 34678
rect 16672 34614 16724 34620
rect 16762 34640 16764 34649
rect 16816 34640 16818 34649
rect 16488 34604 16540 34610
rect 16316 34564 16488 34592
rect 16316 33658 16344 34564
rect 16762 34575 16818 34584
rect 16488 34546 16540 34552
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 16396 33924 16448 33930
rect 16396 33866 16448 33872
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 16304 33652 16356 33658
rect 16304 33594 16356 33600
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 16212 33448 16264 33454
rect 16040 33374 16160 33402
rect 16212 33390 16264 33396
rect 15936 32904 15988 32910
rect 15936 32846 15988 32852
rect 15948 32570 15976 32846
rect 16026 32600 16082 32609
rect 15936 32564 15988 32570
rect 16026 32535 16082 32544
rect 15936 32506 15988 32512
rect 16040 32502 16068 32535
rect 16028 32496 16080 32502
rect 16028 32438 16080 32444
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15752 31758 15804 31764
rect 15842 31784 15898 31793
rect 15842 31719 15898 31728
rect 15752 31680 15804 31686
rect 15948 31668 15976 32370
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 15752 31622 15804 31628
rect 15856 31640 15976 31668
rect 15476 31408 15528 31414
rect 15476 31350 15528 31356
rect 15660 31408 15712 31414
rect 15660 31350 15712 31356
rect 15474 30968 15530 30977
rect 15474 30903 15476 30912
rect 15528 30903 15530 30912
rect 15476 30874 15528 30880
rect 15764 30802 15792 31622
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15672 30394 15700 30534
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15474 30288 15530 30297
rect 15474 30223 15476 30232
rect 15528 30223 15530 30232
rect 15660 30252 15712 30258
rect 15476 30194 15528 30200
rect 15660 30194 15712 30200
rect 15476 29776 15528 29782
rect 15474 29744 15476 29753
rect 15528 29744 15530 29753
rect 15474 29679 15530 29688
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15580 29170 15608 29582
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 15396 28966 15516 28994
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 28150 15332 28358
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15200 27940 15252 27946
rect 15200 27882 15252 27888
rect 15304 27334 15332 28086
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15106 27160 15162 27169
rect 15106 27095 15162 27104
rect 15396 27062 15424 28154
rect 15384 27056 15436 27062
rect 15384 26998 15436 27004
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15028 23662 15056 26862
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15120 26246 15148 26726
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15106 24576 15162 24585
rect 15106 24511 15162 24520
rect 15016 23656 15068 23662
rect 15016 23598 15068 23604
rect 14740 23190 14792 23196
rect 14922 23216 14978 23225
rect 14752 22642 14780 23190
rect 14922 23151 14978 23160
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14660 22234 14688 22578
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14292 20466 14320 20538
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14188 20392 14240 20398
rect 14240 20340 14412 20346
rect 14188 20334 14412 20340
rect 14200 20318 14412 20334
rect 14094 19952 14150 19961
rect 14094 19887 14150 19896
rect 14108 19446 14136 19887
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19553 14228 19654
rect 14186 19544 14242 19553
rect 14186 19479 14242 19488
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14016 19306 14228 19334
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 18290 14044 18566
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14016 17241 14044 18022
rect 14002 17232 14058 17241
rect 14002 17167 14004 17176
rect 14056 17167 14058 17176
rect 14004 17138 14056 17144
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16658 14044 17002
rect 14200 16697 14228 19306
rect 14280 18896 14332 18902
rect 14278 18864 14280 18873
rect 14332 18864 14334 18873
rect 14278 18799 14334 18808
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18329 14320 18702
rect 14278 18320 14334 18329
rect 14278 18255 14334 18264
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 17882 14320 18158
rect 14384 18086 14412 20318
rect 14476 20097 14504 20810
rect 14462 20088 14518 20097
rect 14462 20023 14518 20032
rect 14476 19786 14504 20023
rect 14568 19836 14596 21830
rect 14660 20466 14688 21966
rect 14752 21486 14780 22578
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 21690 14872 22374
rect 14936 22030 14964 23151
rect 15120 23118 15148 24511
rect 15212 23866 15240 26930
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15304 26042 15332 26318
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15304 25294 15332 25638
rect 15396 25430 15424 26318
rect 15488 25906 15516 28966
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15580 27130 15608 27950
rect 15568 27124 15620 27130
rect 15568 27066 15620 27072
rect 15672 26450 15700 30194
rect 15856 30138 15884 31640
rect 16040 31278 16068 31826
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 15934 30288 15990 30297
rect 15934 30223 15936 30232
rect 15988 30223 15990 30232
rect 15936 30194 15988 30200
rect 15856 30110 15976 30138
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15856 29102 15884 29582
rect 15948 29238 15976 30110
rect 16132 29832 16160 33374
rect 16224 32978 16252 33390
rect 16304 33108 16356 33114
rect 16304 33050 16356 33056
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16224 30326 16252 32914
rect 16316 32570 16344 33050
rect 16408 33046 16436 33866
rect 16592 33522 16620 34478
rect 16868 33980 16896 36314
rect 16960 36242 16988 37742
rect 17052 37466 17080 37810
rect 17222 37768 17278 37777
rect 17222 37703 17224 37712
rect 17276 37703 17278 37712
rect 17224 37674 17276 37680
rect 17040 37460 17092 37466
rect 17040 37402 17092 37408
rect 17224 37256 17276 37262
rect 17222 37224 17224 37233
rect 17276 37224 17278 37233
rect 17040 37188 17092 37194
rect 17222 37159 17278 37168
rect 17040 37130 17092 37136
rect 17052 37097 17080 37130
rect 17038 37088 17094 37097
rect 17038 37023 17094 37032
rect 17236 36718 17264 37159
rect 17224 36712 17276 36718
rect 17224 36654 17276 36660
rect 17132 36644 17184 36650
rect 17132 36586 17184 36592
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 17040 36100 17092 36106
rect 17040 36042 17092 36048
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 16960 34746 16988 35566
rect 17052 35222 17080 36042
rect 17144 35601 17172 36586
rect 17130 35592 17186 35601
rect 17130 35527 17186 35536
rect 17040 35216 17092 35222
rect 17040 35158 17092 35164
rect 17144 35154 17172 35527
rect 17236 35442 17264 36654
rect 17328 36378 17356 41386
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 23664 40588 23716 40594
rect 23664 40530 23716 40536
rect 23480 40520 23532 40526
rect 23480 40462 23532 40468
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 23492 39982 23520 40462
rect 17776 39976 17828 39982
rect 17776 39918 17828 39924
rect 23480 39976 23532 39982
rect 23480 39918 23532 39924
rect 17500 38956 17552 38962
rect 17500 38898 17552 38904
rect 17512 38570 17540 38898
rect 17684 38888 17736 38894
rect 17684 38830 17736 38836
rect 17512 38542 17632 38570
rect 17500 38412 17552 38418
rect 17500 38354 17552 38360
rect 17512 37398 17540 38354
rect 17500 37392 17552 37398
rect 17500 37334 17552 37340
rect 17408 37188 17460 37194
rect 17408 37130 17460 37136
rect 17420 36786 17448 37130
rect 17408 36780 17460 36786
rect 17408 36722 17460 36728
rect 17316 36372 17368 36378
rect 17316 36314 17368 36320
rect 17512 36145 17540 37334
rect 17604 37262 17632 38542
rect 17696 38214 17724 38830
rect 17788 38758 17816 39918
rect 18328 39840 18380 39846
rect 18328 39782 18380 39788
rect 23296 39840 23348 39846
rect 23296 39782 23348 39788
rect 18144 39432 18196 39438
rect 18144 39374 18196 39380
rect 17960 39296 18012 39302
rect 17960 39238 18012 39244
rect 17972 38962 18000 39238
rect 18156 39098 18184 39374
rect 18340 39098 18368 39782
rect 22376 39636 22428 39642
rect 22376 39578 22428 39584
rect 22100 39364 22152 39370
rect 22152 39324 22324 39352
rect 22100 39306 22152 39312
rect 18696 39296 18748 39302
rect 18696 39238 18748 39244
rect 21456 39296 21508 39302
rect 21456 39238 21508 39244
rect 18708 39098 18736 39238
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 18144 39092 18196 39098
rect 18144 39034 18196 39040
rect 18328 39092 18380 39098
rect 18328 39034 18380 39040
rect 18696 39092 18748 39098
rect 18696 39034 18748 39040
rect 17960 38956 18012 38962
rect 17960 38898 18012 38904
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 21364 38956 21416 38962
rect 21364 38898 21416 38904
rect 18788 38888 18840 38894
rect 18788 38830 18840 38836
rect 17776 38752 17828 38758
rect 17776 38694 17828 38700
rect 17684 38208 17736 38214
rect 17684 38150 17736 38156
rect 17592 37256 17644 37262
rect 17644 37216 17724 37244
rect 17592 37198 17644 37204
rect 17592 36916 17644 36922
rect 17592 36858 17644 36864
rect 17498 36136 17554 36145
rect 17498 36071 17500 36080
rect 17552 36071 17554 36080
rect 17500 36042 17552 36048
rect 17408 36032 17460 36038
rect 17408 35974 17460 35980
rect 17236 35414 17356 35442
rect 17224 35216 17276 35222
rect 17224 35158 17276 35164
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 16684 33952 16896 33980
rect 16580 33516 16632 33522
rect 16580 33458 16632 33464
rect 16684 33402 16712 33952
rect 17052 33930 17080 34342
rect 17144 34134 17172 34886
rect 17132 34128 17184 34134
rect 17132 34070 17184 34076
rect 17040 33924 17092 33930
rect 17040 33866 17092 33872
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 16592 33374 16712 33402
rect 16396 33040 16448 33046
rect 16396 32982 16448 32988
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16500 32570 16528 32846
rect 16304 32564 16356 32570
rect 16304 32506 16356 32512
rect 16488 32564 16540 32570
rect 16488 32506 16540 32512
rect 16592 32450 16620 33374
rect 16776 32502 16804 33594
rect 17236 33522 17264 35158
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 16856 33312 16908 33318
rect 16856 33254 16908 33260
rect 16868 33114 16896 33254
rect 16856 33108 16908 33114
rect 16856 33050 16908 33056
rect 16948 32768 17000 32774
rect 16948 32710 17000 32716
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 16764 32496 16816 32502
rect 16500 32422 16620 32450
rect 16762 32464 16764 32473
rect 16816 32464 16818 32473
rect 16396 32224 16448 32230
rect 16396 32166 16448 32172
rect 16408 31686 16436 32166
rect 16500 31906 16528 32422
rect 16762 32399 16818 32408
rect 16960 32366 16988 32710
rect 17052 32570 17080 32710
rect 17040 32564 17092 32570
rect 17040 32506 17092 32512
rect 17144 32450 17172 32710
rect 17052 32422 17172 32450
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16592 32026 16620 32302
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16500 31878 16620 31906
rect 16396 31680 16448 31686
rect 16396 31622 16448 31628
rect 16396 31272 16448 31278
rect 16396 31214 16448 31220
rect 16408 31142 16436 31214
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16212 30320 16264 30326
rect 16212 30262 16264 30268
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16224 29850 16252 30126
rect 16040 29804 16160 29832
rect 16212 29844 16264 29850
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15844 29096 15896 29102
rect 15844 29038 15896 29044
rect 15856 28694 15884 29038
rect 15844 28688 15896 28694
rect 15844 28630 15896 28636
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15948 28218 15976 28358
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 16040 27033 16068 29804
rect 16212 29786 16264 29792
rect 16118 29744 16174 29753
rect 16118 29679 16174 29688
rect 16132 29578 16160 29679
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16132 29170 16160 29514
rect 16302 29472 16358 29481
rect 16302 29407 16358 29416
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 16224 27402 16252 27814
rect 16212 27396 16264 27402
rect 16212 27338 16264 27344
rect 16210 27160 16266 27169
rect 16210 27095 16266 27104
rect 16026 27024 16082 27033
rect 16026 26959 16082 26968
rect 16120 26580 16172 26586
rect 16120 26522 16172 26528
rect 15752 26512 15804 26518
rect 15752 26454 15804 26460
rect 16026 26480 16082 26489
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15672 26217 15700 26386
rect 15658 26208 15714 26217
rect 15658 26143 15714 26152
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15672 25906 15700 25978
rect 15476 25900 15528 25906
rect 15660 25900 15712 25906
rect 15476 25842 15528 25848
rect 15580 25860 15660 25888
rect 15384 25424 15436 25430
rect 15384 25366 15436 25372
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15384 25152 15436 25158
rect 15382 25120 15384 25129
rect 15436 25120 15438 25129
rect 15382 25055 15438 25064
rect 15384 24880 15436 24886
rect 15384 24822 15436 24828
rect 15292 24676 15344 24682
rect 15292 24618 15344 24624
rect 15304 24138 15332 24618
rect 15396 24342 15424 24822
rect 15488 24410 15516 25842
rect 15580 24818 15608 25860
rect 15660 25842 15712 25848
rect 15764 25770 15792 26454
rect 16026 26415 16082 26424
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 15856 25906 15884 26182
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15660 25764 15712 25770
rect 15660 25706 15712 25712
rect 15752 25764 15804 25770
rect 15752 25706 15804 25712
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15212 22982 15240 23598
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15028 22409 15056 22578
rect 15014 22400 15070 22409
rect 15014 22335 15070 22344
rect 14924 22024 14976 22030
rect 15016 22024 15068 22030
rect 14924 21966 14976 21972
rect 15014 21992 15016 22001
rect 15068 21992 15070 22001
rect 15014 21927 15070 21936
rect 14922 21720 14978 21729
rect 14832 21684 14884 21690
rect 14978 21678 15056 21706
rect 14922 21655 14978 21664
rect 14832 21626 14884 21632
rect 14924 21616 14976 21622
rect 14844 21564 14924 21570
rect 14844 21558 14976 21564
rect 14844 21542 14964 21558
rect 15028 21554 15056 21678
rect 15120 21554 15148 22714
rect 15016 21548 15068 21554
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14740 21344 14792 21350
rect 14844 21321 14872 21542
rect 15016 21490 15068 21496
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15120 21457 15148 21490
rect 15106 21448 15162 21457
rect 15106 21383 15162 21392
rect 14924 21344 14976 21350
rect 14740 21286 14792 21292
rect 14830 21312 14886 21321
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14648 19848 14700 19854
rect 14568 19808 14648 19836
rect 14648 19790 14700 19796
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 14292 16794 14320 17546
rect 14384 17202 14412 17546
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14186 16688 14242 16697
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 14004 16652 14056 16658
rect 14186 16623 14242 16632
rect 14004 16594 14056 16600
rect 13818 16552 13874 16561
rect 13818 16487 13874 16496
rect 14004 16516 14056 16522
rect 13832 16182 13860 16487
rect 14200 16504 14228 16623
rect 14476 16590 14504 19314
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14568 18698 14596 18838
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14554 18456 14610 18465
rect 14660 18442 14688 19110
rect 14610 18414 14688 18442
rect 14752 18426 14780 21286
rect 14924 21286 14976 21292
rect 14830 21247 14886 21256
rect 14936 21078 14964 21286
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14844 20806 14872 20878
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14830 20360 14886 20369
rect 14936 20346 14964 20742
rect 15028 20534 15056 20742
rect 15120 20602 15148 21383
rect 15212 21350 15240 22918
rect 15304 22166 15332 23666
rect 15488 23202 15516 24346
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15580 24070 15608 24278
rect 15672 24206 15700 25706
rect 15856 25673 15884 25842
rect 15948 25770 15976 26318
rect 15936 25764 15988 25770
rect 15936 25706 15988 25712
rect 15842 25664 15898 25673
rect 15842 25599 15898 25608
rect 15934 25528 15990 25537
rect 15934 25463 15990 25472
rect 15948 25294 15976 25463
rect 16040 25362 16068 26415
rect 16132 26081 16160 26522
rect 16118 26072 16174 26081
rect 16118 26007 16174 26016
rect 16224 25786 16252 27095
rect 16132 25758 16252 25786
rect 16028 25356 16080 25362
rect 16028 25298 16080 25304
rect 15936 25288 15988 25294
rect 15988 25236 16068 25242
rect 15936 25230 16068 25236
rect 15948 25214 16068 25230
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15660 24200 15712 24206
rect 15764 24177 15792 24550
rect 15660 24142 15712 24148
rect 15750 24168 15806 24177
rect 15750 24103 15806 24112
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15396 23174 15516 23202
rect 15396 22778 15424 23174
rect 15580 23066 15608 23462
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15488 23038 15608 23066
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 21418 15332 21898
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15200 20936 15252 20942
rect 15396 20924 15424 22510
rect 15488 22438 15516 23038
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15580 22642 15608 22918
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15488 21690 15516 22374
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15252 20896 15424 20924
rect 15200 20878 15252 20884
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14886 20318 14964 20346
rect 14830 20295 14886 20304
rect 15212 20058 15240 20878
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 14740 18420 14792 18426
rect 14554 18391 14556 18400
rect 14608 18391 14610 18400
rect 14556 18362 14608 18368
rect 14740 18362 14792 18368
rect 14844 18290 14872 19790
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14648 18284 14700 18290
rect 14832 18284 14884 18290
rect 14700 18244 14780 18272
rect 14648 18226 14700 18232
rect 14646 18184 14702 18193
rect 14646 18119 14648 18128
rect 14700 18119 14702 18128
rect 14648 18090 14700 18096
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17728 14596 18022
rect 14752 17796 14780 18244
rect 14832 18226 14884 18232
rect 14936 18154 14964 19246
rect 15028 18970 15056 19654
rect 15120 19514 15148 19790
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15120 19145 15148 19450
rect 15304 19156 15332 19790
rect 15396 19446 15424 19790
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15384 19304 15436 19310
rect 15382 19272 15384 19281
rect 15436 19272 15438 19281
rect 15382 19207 15438 19216
rect 15384 19168 15436 19174
rect 15106 19136 15162 19145
rect 15304 19128 15384 19156
rect 15384 19110 15436 19116
rect 15106 19071 15162 19080
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15028 18766 15056 18906
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15028 18290 15056 18702
rect 15290 18320 15346 18329
rect 15016 18284 15068 18290
rect 15290 18255 15292 18264
rect 15016 18226 15068 18232
rect 15344 18255 15346 18264
rect 15292 18226 15344 18232
rect 15198 18184 15254 18193
rect 14924 18148 14976 18154
rect 15254 18154 15332 18170
rect 15254 18148 15344 18154
rect 15254 18142 15292 18148
rect 15198 18119 15254 18128
rect 14924 18090 14976 18096
rect 15292 18090 15344 18096
rect 14743 17768 14780 17796
rect 15292 17808 15344 17814
rect 14830 17776 14886 17785
rect 14648 17740 14700 17746
rect 14568 17700 14648 17728
rect 14568 17338 14596 17700
rect 14648 17682 14700 17688
rect 14743 17660 14771 17768
rect 14830 17711 14886 17720
rect 15290 17776 15292 17785
rect 15344 17776 15346 17785
rect 15290 17711 15346 17720
rect 14844 17678 14872 17711
rect 15396 17678 15424 19110
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15488 17678 15516 18158
rect 14832 17672 14884 17678
rect 14743 17632 14780 17660
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16590 14688 16934
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14056 16476 14228 16504
rect 14004 16458 14056 16464
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13924 15570 13952 15846
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 15026 13492 15302
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13924 14618 13952 15506
rect 14292 14618 14320 16118
rect 14476 16114 14504 16526
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14476 15026 14504 16050
rect 14752 15570 14780 17632
rect 14832 17614 14884 17620
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14936 17338 14964 17478
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15028 17066 15056 17614
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15120 17241 15148 17478
rect 15106 17232 15162 17241
rect 15304 17202 15332 17478
rect 15106 17167 15162 17176
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 15014 16960 15070 16969
rect 15014 16895 15070 16904
rect 15028 16794 15056 16895
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15396 16726 15424 17614
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15384 16584 15436 16590
rect 15382 16552 15384 16561
rect 15436 16552 15438 16561
rect 15382 16487 15438 16496
rect 15488 16182 15516 16934
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15580 15638 15608 21626
rect 15672 21185 15700 23258
rect 15856 22778 15884 25094
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 15948 24070 15976 24890
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 21418 15792 21830
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15658 21176 15714 21185
rect 15658 21111 15714 21120
rect 15672 19904 15700 21111
rect 15764 20913 15792 21354
rect 15750 20904 15806 20913
rect 15750 20839 15806 20848
rect 15856 20602 15884 22714
rect 15948 22545 15976 23666
rect 16040 22658 16068 25214
rect 16132 24290 16160 25758
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16224 25498 16252 25638
rect 16316 25498 16344 29407
rect 16408 28150 16436 31078
rect 16488 30184 16540 30190
rect 16486 30152 16488 30161
rect 16540 30152 16542 30161
rect 16486 30087 16542 30096
rect 16488 29504 16540 29510
rect 16488 29446 16540 29452
rect 16500 28490 16528 29446
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16396 28144 16448 28150
rect 16396 28086 16448 28092
rect 16486 28112 16542 28121
rect 16486 28047 16488 28056
rect 16540 28047 16542 28056
rect 16488 28018 16540 28024
rect 16394 26616 16450 26625
rect 16394 26551 16450 26560
rect 16408 26382 16436 26551
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16408 25974 16436 26182
rect 16500 26042 16528 26318
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16396 25968 16448 25974
rect 16396 25910 16448 25916
rect 16500 25838 16528 25978
rect 16592 25906 16620 31878
rect 16684 31754 16712 32166
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 16764 31748 16816 31754
rect 16764 31690 16816 31696
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16684 26382 16712 30670
rect 16776 29714 16804 31690
rect 17052 31226 17080 32422
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 17236 31482 17264 32302
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 16868 31198 17080 31226
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 16776 28558 16804 29650
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16776 28218 16804 28494
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16764 28008 16816 28014
rect 16762 27976 16764 27985
rect 16816 27976 16818 27985
rect 16762 27911 16818 27920
rect 16762 27568 16818 27577
rect 16762 27503 16818 27512
rect 16776 27305 16804 27503
rect 16762 27296 16818 27305
rect 16762 27231 16818 27240
rect 16776 26926 16804 27231
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 16684 26042 16712 26182
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16396 25832 16448 25838
rect 16394 25800 16396 25809
rect 16488 25832 16540 25838
rect 16448 25800 16450 25809
rect 16488 25774 16540 25780
rect 16394 25735 16450 25744
rect 16672 25764 16724 25770
rect 16672 25706 16724 25712
rect 16212 25492 16264 25498
rect 16212 25434 16264 25440
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16224 24954 16252 25434
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16316 24970 16344 25230
rect 16316 24954 16528 24970
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16304 24948 16528 24954
rect 16356 24942 16528 24948
rect 16304 24890 16356 24896
rect 16396 24880 16448 24886
rect 16396 24822 16448 24828
rect 16132 24262 16252 24290
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16132 22778 16160 24142
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16040 22630 16160 22658
rect 15934 22536 15990 22545
rect 15934 22471 15990 22480
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21690 15976 21830
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15672 19876 15884 19904
rect 15658 19816 15714 19825
rect 15658 19751 15660 19760
rect 15712 19751 15714 19760
rect 15660 19722 15712 19728
rect 15672 16794 15700 19722
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15764 18766 15792 19450
rect 15856 18970 15884 19876
rect 15948 19378 15976 20742
rect 16040 20602 16068 20878
rect 16132 20874 16160 22630
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16040 19922 16068 20402
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15948 18970 15976 19314
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15856 18834 15884 18906
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15856 18630 15884 18770
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15856 18290 15884 18566
rect 16040 18465 16068 19858
rect 16132 19009 16160 20810
rect 16224 20466 16252 24262
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23526 16344 24006
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16302 23352 16358 23361
rect 16302 23287 16358 23296
rect 16316 22420 16344 23287
rect 16408 22642 16436 24822
rect 16500 24290 16528 24942
rect 16592 24750 16620 25434
rect 16684 25362 16712 25706
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16776 25158 16804 26318
rect 16868 25430 16896 31198
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17144 30598 17172 31078
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 16948 30320 17000 30326
rect 16948 30262 17000 30268
rect 16960 29306 16988 30262
rect 17144 30258 17172 30534
rect 17236 30274 17264 31214
rect 17328 30938 17356 35414
rect 17420 34202 17448 35974
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17408 34196 17460 34202
rect 17408 34138 17460 34144
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17420 30977 17448 33798
rect 17512 33590 17540 34682
rect 17604 33998 17632 36858
rect 17696 35630 17724 37216
rect 17788 36174 17816 38694
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 17880 38282 17908 38490
rect 18420 38344 18472 38350
rect 18420 38286 18472 38292
rect 17868 38276 17920 38282
rect 17868 38218 17920 38224
rect 18328 38004 18380 38010
rect 18248 37964 18328 37992
rect 18052 37460 18104 37466
rect 18052 37402 18104 37408
rect 17868 37120 17920 37126
rect 17868 37062 17920 37068
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17880 35562 17908 37062
rect 17972 36922 18000 37062
rect 17960 36916 18012 36922
rect 17960 36858 18012 36864
rect 17960 36644 18012 36650
rect 17960 36586 18012 36592
rect 17972 36174 18000 36586
rect 17960 36168 18012 36174
rect 17960 36110 18012 36116
rect 17868 35556 17920 35562
rect 17868 35498 17920 35504
rect 17592 33992 17644 33998
rect 17592 33934 17644 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17788 32910 17816 33934
rect 17972 33930 18000 36110
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17880 32774 17908 33458
rect 17972 33454 18000 33866
rect 18064 33658 18092 37402
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 18156 35494 18184 35974
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 18156 33658 18184 35430
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 18144 33652 18196 33658
rect 18144 33594 18196 33600
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 18156 33046 18184 33594
rect 18144 33040 18196 33046
rect 18144 32982 18196 32988
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17406 30968 17462 30977
rect 17316 30932 17368 30938
rect 17604 30938 17632 31690
rect 17880 31482 17908 32506
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17972 32026 18000 32234
rect 17960 32020 18012 32026
rect 17960 31962 18012 31968
rect 18052 31952 18104 31958
rect 18050 31920 18052 31929
rect 18104 31920 18106 31929
rect 18156 31890 18184 32982
rect 18050 31855 18106 31864
rect 18144 31884 18196 31890
rect 18144 31826 18196 31832
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17696 31249 17724 31282
rect 17682 31240 17738 31249
rect 17682 31175 17738 31184
rect 17880 31142 17908 31282
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17406 30903 17462 30912
rect 17592 30932 17644 30938
rect 17316 30874 17368 30880
rect 17592 30874 17644 30880
rect 17316 30728 17368 30734
rect 17314 30696 17316 30705
rect 17776 30728 17828 30734
rect 17368 30696 17370 30705
rect 17776 30670 17828 30676
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17314 30631 17370 30640
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 17132 30252 17184 30258
rect 17236 30246 17448 30274
rect 17132 30194 17184 30200
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 17038 29336 17094 29345
rect 16948 29300 17000 29306
rect 17038 29271 17094 29280
rect 16948 29242 17000 29248
rect 17052 29238 17080 29271
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 27674 16988 28358
rect 17040 27940 17092 27946
rect 17040 27882 17092 27888
rect 16948 27668 17000 27674
rect 16948 27610 17000 27616
rect 17052 27305 17080 27882
rect 17038 27296 17094 27305
rect 17038 27231 17094 27240
rect 17144 27130 17172 30058
rect 17224 30048 17276 30054
rect 17224 29990 17276 29996
rect 17236 29850 17264 29990
rect 17224 29844 17276 29850
rect 17224 29786 17276 29792
rect 17420 29696 17448 30246
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17236 29668 17448 29696
rect 17236 27614 17264 29668
rect 17512 29170 17540 30194
rect 17604 29646 17632 30194
rect 17696 30054 17724 30602
rect 17788 30394 17816 30670
rect 17972 30433 18000 30670
rect 17958 30424 18014 30433
rect 17776 30388 17828 30394
rect 17958 30359 18014 30368
rect 17776 30330 17828 30336
rect 17684 30048 17736 30054
rect 17684 29990 17736 29996
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17328 28762 17356 29038
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17328 27985 17356 28494
rect 17314 27976 17370 27985
rect 17314 27911 17370 27920
rect 17236 27586 17356 27614
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 17236 27062 17264 27406
rect 17224 27056 17276 27062
rect 17224 26998 17276 27004
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 16948 26512 17000 26518
rect 16948 26454 17000 26460
rect 16960 26314 16988 26454
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 17236 26246 17264 26862
rect 17328 26790 17356 27586
rect 17420 27418 17448 29106
rect 17696 28966 17724 29990
rect 17788 29578 17816 30330
rect 17958 30288 18014 30297
rect 17958 30223 17960 30232
rect 18012 30223 18014 30232
rect 17960 30194 18012 30200
rect 17866 29880 17922 29889
rect 17866 29815 17922 29824
rect 17776 29572 17828 29578
rect 17776 29514 17828 29520
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 17684 28960 17736 28966
rect 17684 28902 17736 28908
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 28098 17540 28358
rect 17512 28082 17632 28098
rect 17512 28076 17644 28082
rect 17512 28070 17592 28076
rect 17592 28018 17644 28024
rect 17684 28008 17736 28014
rect 17604 27956 17684 27962
rect 17604 27950 17736 27956
rect 17604 27934 17724 27950
rect 17604 27878 17632 27934
rect 17788 27878 17816 29038
rect 17880 28994 17908 29815
rect 17880 28966 18000 28994
rect 17972 28762 18000 28966
rect 17960 28756 18012 28762
rect 17960 28698 18012 28704
rect 17868 28688 17920 28694
rect 17868 28630 17920 28636
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17776 27872 17828 27878
rect 17776 27814 17828 27820
rect 17774 27568 17830 27577
rect 17774 27503 17830 27512
rect 17420 27390 17540 27418
rect 17408 27328 17460 27334
rect 17406 27296 17408 27305
rect 17460 27296 17462 27305
rect 17406 27231 17462 27240
rect 17420 26994 17448 27231
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17406 26888 17462 26897
rect 17406 26823 17462 26832
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17314 26344 17370 26353
rect 17420 26330 17448 26823
rect 17370 26302 17448 26330
rect 17314 26279 17316 26288
rect 17368 26279 17370 26288
rect 17316 26250 17368 26256
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 16856 25424 16908 25430
rect 16856 25366 16908 25372
rect 17040 25220 17092 25226
rect 17040 25162 17092 25168
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16670 24984 16726 24993
rect 16670 24919 16726 24928
rect 16684 24800 16712 24919
rect 16764 24812 16816 24818
rect 16684 24772 16764 24800
rect 16764 24754 16816 24760
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16592 24410 16620 24686
rect 16764 24676 16816 24682
rect 16764 24618 16816 24624
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16672 24336 16724 24342
rect 16500 24262 16620 24290
rect 16672 24278 16724 24284
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16396 22432 16448 22438
rect 16316 22392 16396 22420
rect 16396 22374 16448 22380
rect 16408 22114 16436 22374
rect 16500 22234 16528 24142
rect 16592 23050 16620 24262
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16684 22506 16712 24278
rect 16776 23730 16804 24618
rect 16868 24313 16896 24754
rect 16854 24304 16910 24313
rect 16854 24239 16910 24248
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16776 23118 16804 23462
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16592 22234 16620 22374
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16486 22128 16542 22137
rect 16304 22092 16356 22098
rect 16408 22086 16486 22114
rect 16486 22063 16542 22072
rect 16304 22034 16356 22040
rect 16316 21690 16344 22034
rect 16580 22024 16632 22030
rect 16500 21984 16580 22012
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16408 21690 16436 21830
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16316 20874 16344 21422
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16408 20602 16436 21490
rect 16500 21321 16528 21984
rect 16580 21966 16632 21972
rect 16578 21584 16634 21593
rect 16578 21519 16580 21528
rect 16632 21519 16634 21528
rect 16580 21490 16632 21496
rect 16486 21312 16542 21321
rect 16486 21247 16542 21256
rect 16592 20913 16620 21490
rect 16684 21350 16712 22442
rect 16776 21554 16804 22510
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16762 21448 16818 21457
rect 16762 21383 16818 21392
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16578 20904 16634 20913
rect 16488 20868 16540 20874
rect 16578 20839 16634 20848
rect 16488 20810 16540 20816
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16212 19984 16264 19990
rect 16408 19961 16436 20198
rect 16212 19926 16264 19932
rect 16394 19952 16450 19961
rect 16118 19000 16174 19009
rect 16118 18935 16120 18944
rect 16172 18935 16174 18944
rect 16120 18906 16172 18912
rect 16118 18864 16174 18873
rect 16118 18799 16174 18808
rect 16132 18766 16160 18799
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16026 18456 16082 18465
rect 15936 18420 15988 18426
rect 16026 18391 16082 18400
rect 15936 18362 15988 18368
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15764 17105 15792 17682
rect 15856 17678 15884 18226
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15948 17270 15976 18362
rect 16040 18222 16068 18391
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15948 16726 15976 17206
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16040 15638 16068 18158
rect 16132 16250 16160 18702
rect 16224 17649 16252 19926
rect 16394 19887 16450 19896
rect 16500 19334 16528 20810
rect 16580 20800 16632 20806
rect 16578 20768 16580 20777
rect 16632 20768 16634 20777
rect 16578 20703 16634 20712
rect 16408 19306 16528 19334
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18068 16344 18702
rect 16408 18193 16436 19306
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18465 16528 18702
rect 16486 18456 16542 18465
rect 16486 18391 16488 18400
rect 16540 18391 16542 18400
rect 16488 18362 16540 18368
rect 16592 18358 16620 20703
rect 16684 19514 16712 21286
rect 16776 19990 16804 21383
rect 16868 20398 16896 24239
rect 16960 24206 16988 25094
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 17052 23474 17080 25162
rect 17144 23594 17172 25434
rect 17236 24993 17264 26182
rect 17512 25702 17540 27390
rect 17590 27296 17646 27305
rect 17590 27231 17646 27240
rect 17604 26364 17632 27231
rect 17684 26852 17736 26858
rect 17684 26794 17736 26800
rect 17696 26586 17724 26794
rect 17788 26586 17816 27503
rect 17880 27470 17908 28630
rect 18064 28404 18092 31214
rect 18156 30938 18184 31826
rect 18144 30932 18196 30938
rect 18144 30874 18196 30880
rect 18142 29608 18198 29617
rect 18142 29543 18198 29552
rect 18156 29306 18184 29543
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18156 28490 18184 29106
rect 18248 28994 18276 37964
rect 18432 37992 18460 38286
rect 18604 38208 18656 38214
rect 18604 38150 18656 38156
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 18432 37964 18552 37992
rect 18328 37946 18380 37952
rect 18420 37800 18472 37806
rect 18420 37742 18472 37748
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 18340 35834 18368 37674
rect 18432 36922 18460 37742
rect 18524 37670 18552 37964
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 18420 36916 18472 36922
rect 18420 36858 18472 36864
rect 18616 36718 18644 38150
rect 18708 37942 18736 38150
rect 18696 37936 18748 37942
rect 18696 37878 18748 37884
rect 18800 37754 18828 38830
rect 19616 38752 19668 38758
rect 19616 38694 19668 38700
rect 19628 38350 19656 38694
rect 19616 38344 19668 38350
rect 19616 38286 19668 38292
rect 19996 38282 20024 38898
rect 20260 38752 20312 38758
rect 20260 38694 20312 38700
rect 20444 38752 20496 38758
rect 20444 38694 20496 38700
rect 21272 38752 21324 38758
rect 21272 38694 21324 38700
rect 20168 38548 20220 38554
rect 20168 38490 20220 38496
rect 19984 38276 20036 38282
rect 19984 38218 20036 38224
rect 20076 38208 20128 38214
rect 20076 38150 20128 38156
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 20088 37942 20116 38150
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 19248 37868 19300 37874
rect 19248 37810 19300 37816
rect 18708 37726 18828 37754
rect 18880 37800 18932 37806
rect 18880 37742 18932 37748
rect 18708 36718 18736 37726
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 18800 37262 18828 37606
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 18604 36712 18656 36718
rect 18604 36654 18656 36660
rect 18696 36712 18748 36718
rect 18696 36654 18748 36660
rect 18512 36576 18564 36582
rect 18432 36536 18512 36564
rect 18328 35828 18380 35834
rect 18328 35770 18380 35776
rect 18328 35692 18380 35698
rect 18328 35634 18380 35640
rect 18340 35290 18368 35634
rect 18328 35284 18380 35290
rect 18328 35226 18380 35232
rect 18432 34184 18460 36536
rect 18512 36518 18564 36524
rect 18616 36174 18644 36654
rect 18512 36168 18564 36174
rect 18512 36110 18564 36116
rect 18604 36168 18656 36174
rect 18604 36110 18656 36116
rect 18524 35834 18552 36110
rect 18512 35828 18564 35834
rect 18512 35770 18564 35776
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18524 34649 18552 35022
rect 18616 34950 18644 36110
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 18604 34944 18656 34950
rect 18604 34886 18656 34892
rect 18510 34640 18566 34649
rect 18510 34575 18566 34584
rect 18340 34156 18460 34184
rect 18340 31414 18368 34156
rect 18524 33454 18552 34575
rect 18708 34542 18736 35158
rect 18696 34536 18748 34542
rect 18696 34478 18748 34484
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18512 33448 18564 33454
rect 18512 33390 18564 33396
rect 18616 33046 18644 34002
rect 18788 33992 18840 33998
rect 18788 33934 18840 33940
rect 18800 33862 18828 33934
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18604 33040 18656 33046
rect 18604 32982 18656 32988
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18432 31482 18460 32846
rect 18512 32836 18564 32842
rect 18512 32778 18564 32784
rect 18524 32745 18552 32778
rect 18510 32736 18566 32745
rect 18510 32671 18566 32680
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18524 32026 18552 32370
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18616 31872 18644 32166
rect 18694 32056 18750 32065
rect 18694 31991 18750 32000
rect 18524 31844 18644 31872
rect 18420 31476 18472 31482
rect 18420 31418 18472 31424
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 18524 31346 18552 31844
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18420 31136 18472 31142
rect 18616 31113 18644 31418
rect 18420 31078 18472 31084
rect 18602 31104 18658 31113
rect 18432 30734 18460 31078
rect 18602 31039 18658 31048
rect 18510 30968 18566 30977
rect 18708 30938 18736 31991
rect 18800 31754 18828 33798
rect 18892 33318 18920 37742
rect 19260 37330 19288 37810
rect 19248 37324 19300 37330
rect 19248 37266 19300 37272
rect 19246 37224 19302 37233
rect 19246 37159 19248 37168
rect 19300 37159 19302 37168
rect 19248 37130 19300 37136
rect 19156 37120 19208 37126
rect 19156 37062 19208 37068
rect 19168 36922 19196 37062
rect 19156 36916 19208 36922
rect 19156 36858 19208 36864
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19156 36644 19208 36650
rect 19156 36586 19208 36592
rect 19168 35494 19196 36586
rect 19260 36378 19288 36654
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19248 36372 19300 36378
rect 19248 36314 19300 36320
rect 19352 35698 19380 36518
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19156 35488 19208 35494
rect 19156 35430 19208 35436
rect 19444 35222 19472 37878
rect 20180 37874 20208 38490
rect 20272 38486 20300 38694
rect 20260 38480 20312 38486
rect 20260 38422 20312 38428
rect 20352 38208 20404 38214
rect 20352 38150 20404 38156
rect 20364 37992 20392 38150
rect 20272 37964 20392 37992
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 19812 37262 19840 37402
rect 19800 37256 19852 37262
rect 19800 37198 19852 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20180 36122 20208 37810
rect 20272 36378 20300 37964
rect 20456 37330 20484 38694
rect 21178 38584 21234 38593
rect 21178 38519 21180 38528
rect 21232 38519 21234 38528
rect 21180 38490 21232 38496
rect 20536 38480 20588 38486
rect 20536 38422 20588 38428
rect 20718 38448 20774 38457
rect 20548 37874 20576 38422
rect 20718 38383 20720 38392
rect 20772 38383 20774 38392
rect 20720 38354 20772 38360
rect 21284 38282 21312 38694
rect 21376 38350 21404 38898
rect 21364 38344 21416 38350
rect 21364 38286 21416 38292
rect 21272 38276 21324 38282
rect 21272 38218 21324 38224
rect 21284 38185 21312 38218
rect 21270 38176 21326 38185
rect 21270 38111 21326 38120
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20732 37874 20760 37946
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20548 37754 20576 37810
rect 20548 37726 20668 37754
rect 20640 37720 20668 37726
rect 20812 37732 20864 37738
rect 20640 37692 20812 37720
rect 20812 37674 20864 37680
rect 21284 37670 21312 38111
rect 21376 37806 21404 38286
rect 21468 38214 21496 39238
rect 21916 38956 21968 38962
rect 21916 38898 21968 38904
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 21640 38752 21692 38758
rect 21640 38694 21692 38700
rect 21548 38480 21600 38486
rect 21652 38457 21680 38694
rect 21548 38422 21600 38428
rect 21638 38448 21694 38457
rect 21456 38208 21508 38214
rect 21456 38150 21508 38156
rect 21364 37800 21416 37806
rect 21364 37742 21416 37748
rect 20536 37664 20588 37670
rect 20536 37606 20588 37612
rect 21272 37664 21324 37670
rect 21272 37606 21324 37612
rect 20444 37324 20496 37330
rect 20444 37266 20496 37272
rect 20352 36576 20404 36582
rect 20352 36518 20404 36524
rect 20260 36372 20312 36378
rect 20260 36314 20312 36320
rect 20088 36094 20208 36122
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20088 35222 20116 36094
rect 20168 36032 20220 36038
rect 20168 35974 20220 35980
rect 20180 35698 20208 35974
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 19432 35216 19484 35222
rect 19432 35158 19484 35164
rect 20076 35216 20128 35222
rect 20076 35158 20128 35164
rect 20076 35080 20128 35086
rect 20076 35022 20128 35028
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 19982 34912 20038 34921
rect 19076 34610 19104 34886
rect 19574 34844 19882 34853
rect 19982 34847 20038 34856
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 19064 34604 19116 34610
rect 19064 34546 19116 34552
rect 19156 34536 19208 34542
rect 19156 34478 19208 34484
rect 18972 33992 19024 33998
rect 18972 33934 19024 33940
rect 18984 33658 19012 33934
rect 18972 33652 19024 33658
rect 18972 33594 19024 33600
rect 19168 33522 19196 34478
rect 19444 33522 19472 34614
rect 19892 34604 19944 34610
rect 19996 34592 20024 34847
rect 20088 34746 20116 35022
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19944 34564 20024 34592
rect 19892 34546 19944 34552
rect 19708 34536 19760 34542
rect 19708 34478 19760 34484
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19628 33998 19656 34138
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19720 33980 19748 34478
rect 20364 34134 20392 36518
rect 20548 35766 20576 37606
rect 20812 37120 20864 37126
rect 20812 37062 20864 37068
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20824 36922 20852 37062
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20628 36576 20680 36582
rect 20628 36518 20680 36524
rect 20640 36106 20668 36518
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 20536 35760 20588 35766
rect 20536 35702 20588 35708
rect 21008 35222 21036 37062
rect 20996 35216 21048 35222
rect 20996 35158 21048 35164
rect 20904 35012 20956 35018
rect 20904 34954 20956 34960
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20732 34746 20760 34886
rect 20916 34746 20944 34954
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20352 34128 20404 34134
rect 20352 34070 20404 34076
rect 19892 33992 19944 33998
rect 19720 33952 19892 33980
rect 19720 33862 19748 33952
rect 19892 33934 19944 33940
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 19708 33856 19760 33862
rect 19708 33798 19760 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 19156 33516 19208 33522
rect 19156 33458 19208 33464
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 19076 32910 19104 33458
rect 19168 32910 19196 33458
rect 19064 32904 19116 32910
rect 18878 32872 18934 32881
rect 19064 32846 19116 32852
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 18878 32807 18934 32816
rect 18892 32212 18920 32807
rect 19064 32768 19116 32774
rect 19064 32710 19116 32716
rect 18972 32224 19024 32230
rect 18892 32184 18972 32212
rect 18972 32166 19024 32172
rect 18800 31726 18920 31754
rect 18788 31408 18840 31414
rect 18788 31350 18840 31356
rect 18510 30903 18566 30912
rect 18604 30932 18656 30938
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18340 30569 18368 30670
rect 18524 30666 18552 30903
rect 18604 30874 18656 30880
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18616 30666 18644 30874
rect 18696 30796 18748 30802
rect 18696 30738 18748 30744
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18604 30660 18656 30666
rect 18604 30602 18656 30608
rect 18326 30560 18382 30569
rect 18326 30495 18382 30504
rect 18604 30320 18656 30326
rect 18604 30262 18656 30268
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18340 29510 18368 29990
rect 18512 29572 18564 29578
rect 18512 29514 18564 29520
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18524 29306 18552 29514
rect 18616 29481 18644 30262
rect 18602 29472 18658 29481
rect 18602 29407 18658 29416
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18420 29232 18472 29238
rect 18420 29174 18472 29180
rect 18248 28966 18368 28994
rect 18144 28484 18196 28490
rect 18144 28426 18196 28432
rect 17972 28376 18092 28404
rect 17972 27674 18000 28376
rect 18142 28248 18198 28257
rect 18142 28183 18198 28192
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 18064 27130 18092 27338
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17776 26376 17828 26382
rect 17604 26336 17776 26364
rect 17776 26318 17828 26324
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17512 25498 17540 25638
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17408 25288 17460 25294
rect 17512 25265 17540 25298
rect 17408 25230 17460 25236
rect 17498 25256 17554 25265
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17222 24984 17278 24993
rect 17222 24919 17278 24928
rect 17328 24818 17356 25094
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17328 24342 17356 24754
rect 17224 24336 17276 24342
rect 17222 24304 17224 24313
rect 17316 24336 17368 24342
rect 17276 24304 17278 24313
rect 17316 24278 17368 24284
rect 17222 24239 17278 24248
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17132 23588 17184 23594
rect 17132 23530 17184 23536
rect 16960 23446 17080 23474
rect 16960 22234 16988 23446
rect 17040 23316 17092 23322
rect 17144 23304 17172 23530
rect 17236 23322 17264 24142
rect 17328 24138 17356 24278
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 17314 23760 17370 23769
rect 17314 23695 17370 23704
rect 17092 23276 17172 23304
rect 17224 23316 17276 23322
rect 17040 23258 17092 23264
rect 17224 23258 17276 23264
rect 17328 23254 17356 23695
rect 17316 23248 17368 23254
rect 17038 23216 17094 23225
rect 17038 23151 17094 23160
rect 17222 23216 17278 23225
rect 17316 23190 17368 23196
rect 17222 23151 17278 23160
rect 17052 23050 17080 23151
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16946 22128 17002 22137
rect 16946 22063 17002 22072
rect 16960 21962 16988 22063
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 17052 21842 17080 22986
rect 17236 22681 17264 23151
rect 17328 23089 17356 23190
rect 17314 23080 17370 23089
rect 17314 23015 17370 23024
rect 17316 22976 17368 22982
rect 17314 22944 17316 22953
rect 17368 22944 17370 22953
rect 17314 22879 17370 22888
rect 17222 22672 17278 22681
rect 17222 22607 17224 22616
rect 17276 22607 17278 22616
rect 17224 22578 17276 22584
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 16960 21814 17080 21842
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16868 19990 16896 20334
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16776 19514 16804 19790
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16684 18426 16712 19450
rect 16762 18864 16818 18873
rect 16960 18850 16988 21814
rect 17144 21554 17172 22374
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17130 21448 17186 21457
rect 17040 21412 17092 21418
rect 17130 21383 17132 21392
rect 17040 21354 17092 21360
rect 17184 21383 17186 21392
rect 17132 21354 17184 21360
rect 17052 20330 17080 21354
rect 17144 20466 17172 21354
rect 17236 21078 17264 22578
rect 17316 22568 17368 22574
rect 17420 22545 17448 25230
rect 17498 25191 17554 25200
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17512 24614 17540 25094
rect 17604 24750 17632 25162
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 23798 17540 24550
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17604 23100 17632 23598
rect 17696 23497 17724 24754
rect 17788 24070 17816 25434
rect 17776 24064 17828 24070
rect 17880 24041 17908 26726
rect 17972 26586 18000 26726
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 18050 26344 18106 26353
rect 18050 26279 18106 26288
rect 17960 25968 18012 25974
rect 17960 25910 18012 25916
rect 17972 24410 18000 25910
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 18064 24274 18092 26279
rect 18156 25809 18184 28183
rect 18234 27840 18290 27849
rect 18234 27775 18290 27784
rect 18248 26382 18276 27775
rect 18340 27130 18368 28966
rect 18432 28150 18460 29174
rect 18604 28688 18656 28694
rect 18602 28656 18604 28665
rect 18656 28656 18658 28665
rect 18602 28591 18658 28600
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 18420 27872 18472 27878
rect 18616 27849 18644 28494
rect 18420 27814 18472 27820
rect 18602 27840 18658 27849
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18432 26994 18460 27814
rect 18602 27775 18658 27784
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18616 26926 18644 27066
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18326 26616 18382 26625
rect 18326 26551 18382 26560
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18142 25800 18198 25809
rect 18142 25735 18198 25744
rect 18236 25764 18288 25770
rect 18236 25706 18288 25712
rect 18248 25430 18276 25706
rect 18236 25424 18288 25430
rect 18236 25366 18288 25372
rect 18340 24818 18368 26551
rect 18420 26444 18472 26450
rect 18420 26386 18472 26392
rect 18432 25498 18460 26386
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18524 25401 18552 25638
rect 18510 25392 18566 25401
rect 18510 25327 18566 25336
rect 18512 25288 18564 25294
rect 18432 25248 18512 25276
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17776 24006 17828 24012
rect 17866 24032 17922 24041
rect 17866 23967 17922 23976
rect 17972 23798 18000 24142
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17682 23488 17738 23497
rect 17682 23423 17738 23432
rect 17788 23225 17816 23666
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17774 23216 17830 23225
rect 17774 23151 17830 23160
rect 17776 23112 17828 23118
rect 17604 23072 17776 23100
rect 17776 23054 17828 23060
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17316 22510 17368 22516
rect 17406 22536 17462 22545
rect 17328 22166 17356 22510
rect 17406 22471 17462 22480
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17420 22030 17448 22471
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20466 17264 20878
rect 17328 20641 17356 21286
rect 17314 20632 17370 20641
rect 17314 20567 17370 20576
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17052 19310 17080 19790
rect 17236 19378 17264 20402
rect 17328 19786 17356 20402
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16818 18822 16988 18850
rect 16762 18799 16818 18808
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16394 18184 16450 18193
rect 16394 18119 16450 18128
rect 16316 18040 16528 18068
rect 16302 17912 16358 17921
rect 16302 17847 16358 17856
rect 16210 17640 16266 17649
rect 16210 17575 16266 17584
rect 16316 17542 16344 17847
rect 16500 17610 16528 18040
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16224 17048 16252 17478
rect 16316 17270 16344 17478
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 16304 17060 16356 17066
rect 16224 17020 16304 17048
rect 16304 17002 16356 17008
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16316 15638 16344 16594
rect 16500 16454 16528 17546
rect 16592 16969 16620 17614
rect 16578 16960 16634 16969
rect 16578 16895 16634 16904
rect 16776 16794 16804 18702
rect 17144 18630 17172 19314
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 18290 17172 18566
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17052 17882 17080 18090
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16960 17678 16988 17750
rect 16856 17672 16908 17678
rect 16854 17640 16856 17649
rect 16948 17672 17000 17678
rect 16908 17640 16910 17649
rect 16948 17614 17000 17620
rect 16854 17575 16910 17584
rect 17052 16794 17080 17818
rect 17236 17134 17264 19314
rect 17314 19272 17370 19281
rect 17314 19207 17370 19216
rect 17328 18902 17356 19207
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17420 18222 17448 21966
rect 17512 21962 17540 22918
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17592 22432 17644 22438
rect 17590 22400 17592 22409
rect 17644 22400 17646 22409
rect 17590 22335 17646 22344
rect 17696 22098 17724 22578
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17498 21856 17554 21865
rect 17498 21791 17554 21800
rect 17512 21690 17540 21791
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17498 21448 17554 21457
rect 17498 21383 17554 21392
rect 17512 21350 17540 21383
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17512 21146 17540 21286
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17512 20262 17540 21082
rect 17604 21010 17632 21966
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17696 21554 17724 21898
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 20534 17632 20742
rect 17696 20602 17724 21490
rect 17788 21026 17816 23054
rect 17880 21865 17908 23598
rect 18156 23594 18184 24550
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 18064 23225 18092 23462
rect 18050 23216 18106 23225
rect 18050 23151 18106 23160
rect 18064 22982 18092 23151
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18064 22778 18092 22918
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17972 22438 18000 22646
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17866 21856 17922 21865
rect 17866 21791 17922 21800
rect 17972 21350 18000 22374
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18064 21622 18092 21830
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 21350 18092 21422
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18050 21040 18106 21049
rect 17788 20998 17908 21026
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 19854 17632 20198
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17590 19272 17646 19281
rect 17500 19236 17552 19242
rect 17590 19207 17646 19216
rect 17500 19178 17552 19184
rect 17512 18290 17540 19178
rect 17604 18329 17632 19207
rect 17590 18320 17646 18329
rect 17500 18284 17552 18290
rect 17696 18290 17724 19994
rect 17788 19854 17816 20402
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17788 19446 17816 19790
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17880 18970 17908 20998
rect 18050 20975 18052 20984
rect 18104 20975 18106 20984
rect 18052 20946 18104 20952
rect 18156 20874 18184 23530
rect 18248 22386 18276 24754
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18340 23322 18368 24006
rect 18432 23594 18460 25248
rect 18512 25230 18564 25236
rect 18616 24750 18644 25842
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18512 24336 18564 24342
rect 18512 24278 18564 24284
rect 18524 23798 18552 24278
rect 18604 24200 18656 24206
rect 18602 24168 18604 24177
rect 18656 24168 18658 24177
rect 18602 24103 18658 24112
rect 18512 23792 18564 23798
rect 18564 23752 18644 23780
rect 18512 23734 18564 23740
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18510 23352 18566 23361
rect 18328 23316 18380 23322
rect 18510 23287 18566 23296
rect 18328 23258 18380 23264
rect 18420 23112 18472 23118
rect 18326 23080 18382 23089
rect 18420 23054 18472 23060
rect 18326 23015 18328 23024
rect 18380 23015 18382 23024
rect 18328 22986 18380 22992
rect 18432 22642 18460 23054
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18524 22574 18552 23287
rect 18512 22568 18564 22574
rect 18512 22510 18564 22516
rect 18420 22432 18472 22438
rect 18248 22358 18368 22386
rect 18420 22374 18472 22380
rect 18340 22273 18368 22358
rect 18326 22264 18382 22273
rect 18236 22228 18288 22234
rect 18326 22199 18382 22208
rect 18236 22170 18288 22176
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17972 18766 18000 20538
rect 18064 19281 18092 20810
rect 18156 20602 18184 20810
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18050 19272 18106 19281
rect 18156 19242 18184 20402
rect 18248 19938 18276 22170
rect 18432 22094 18460 22374
rect 18510 22264 18566 22273
rect 18510 22199 18566 22208
rect 18340 22066 18460 22094
rect 18340 20466 18368 22066
rect 18420 22024 18472 22030
rect 18524 22012 18552 22199
rect 18472 21984 18552 22012
rect 18420 21966 18472 21972
rect 18432 20806 18460 21966
rect 18616 21944 18644 23752
rect 18708 22438 18736 30738
rect 18800 30666 18828 31350
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18892 30138 18920 31726
rect 18984 31260 19012 32166
rect 19076 32026 19104 32710
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 19168 31958 19196 32846
rect 19444 32502 19472 33458
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19996 33114 20024 33254
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 20076 33108 20128 33114
rect 20076 33050 20128 33056
rect 19984 32972 20036 32978
rect 20088 32960 20116 33050
rect 20036 32932 20116 32960
rect 20168 32972 20220 32978
rect 19984 32914 20036 32920
rect 20364 32960 20392 33934
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20220 32932 20392 32960
rect 20168 32914 20220 32920
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 20076 32768 20128 32774
rect 20076 32710 20128 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19156 31952 19208 31958
rect 19156 31894 19208 31900
rect 19260 31482 19288 32370
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19248 31476 19300 31482
rect 19248 31418 19300 31424
rect 19154 31376 19210 31385
rect 19154 31311 19156 31320
rect 19208 31311 19210 31320
rect 19156 31282 19208 31288
rect 19064 31272 19116 31278
rect 18984 31232 19064 31260
rect 19064 31214 19116 31220
rect 19154 31240 19210 31249
rect 19154 31175 19156 31184
rect 19208 31175 19210 31184
rect 19248 31204 19300 31210
rect 19156 31146 19208 31152
rect 19248 31146 19300 31152
rect 19168 30682 19196 31146
rect 19260 30734 19288 31146
rect 19352 30802 19380 32302
rect 19444 31890 19472 32438
rect 19996 32434 20024 32710
rect 20088 32570 20116 32710
rect 20076 32564 20128 32570
rect 20076 32506 20128 32512
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 19616 32020 19668 32026
rect 19616 31962 19668 31968
rect 19432 31884 19484 31890
rect 19432 31826 19484 31832
rect 19524 31680 19576 31686
rect 19511 31628 19524 31668
rect 19628 31668 19656 31962
rect 19892 31816 19944 31822
rect 19944 31776 20024 31804
rect 19892 31758 19944 31764
rect 19576 31640 19656 31668
rect 19511 31622 19576 31628
rect 19423 31476 19475 31482
rect 19511 31464 19539 31622
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31482 20024 31776
rect 19984 31476 20036 31482
rect 19511 31436 19748 31464
rect 19423 31418 19475 31424
rect 19444 31362 19472 31418
rect 19444 31334 19656 31362
rect 19720 31346 19748 31436
rect 19984 31418 20036 31424
rect 20088 31346 20116 32166
rect 20272 32026 20300 32932
rect 20456 32570 20484 33458
rect 20536 33312 20588 33318
rect 20536 33254 20588 33260
rect 20548 32978 20576 33254
rect 20536 32972 20588 32978
rect 20536 32914 20588 32920
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20444 32428 20496 32434
rect 20496 32388 20576 32416
rect 20444 32370 20496 32376
rect 20352 32224 20404 32230
rect 20352 32166 20404 32172
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20260 31748 20312 31754
rect 20260 31690 20312 31696
rect 20166 31376 20222 31385
rect 19522 30832 19578 30841
rect 19340 30796 19392 30802
rect 19392 30776 19522 30784
rect 19392 30767 19578 30776
rect 19392 30756 19564 30767
rect 19340 30738 19392 30744
rect 18800 30110 18920 30138
rect 18984 30654 19196 30682
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 19340 30660 19392 30666
rect 18800 26790 18828 30110
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18892 29306 18920 29990
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18984 28694 19012 30654
rect 19392 30620 19472 30648
rect 19340 30602 19392 30608
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19168 30297 19196 30534
rect 19154 30288 19210 30297
rect 19154 30223 19210 30232
rect 19064 30116 19116 30122
rect 19064 30058 19116 30064
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19076 29850 19104 30058
rect 19168 30025 19196 30058
rect 19154 30016 19210 30025
rect 19154 29951 19210 29960
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 19260 29306 19288 30534
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19168 28966 19196 29106
rect 19352 29102 19380 29990
rect 19444 29288 19472 30620
rect 19628 30580 19656 31334
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 20076 31340 20128 31346
rect 20166 31311 20222 31320
rect 20076 31282 20128 31288
rect 19511 30552 19656 30580
rect 19511 30376 19539 30552
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19511 30348 19564 30376
rect 19536 30122 19564 30348
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19524 30116 19576 30122
rect 19524 30058 19576 30064
rect 19812 29646 19840 30126
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19616 29300 19668 29306
rect 19444 29260 19564 29288
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 19064 28960 19116 28966
rect 19064 28902 19116 28908
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19076 28778 19104 28902
rect 19076 28750 19196 28778
rect 18972 28688 19024 28694
rect 18892 28648 18972 28676
rect 18892 27554 18920 28648
rect 18972 28630 19024 28636
rect 19168 28558 19196 28750
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 19156 28552 19208 28558
rect 19156 28494 19208 28500
rect 19338 28520 19394 28529
rect 18984 28014 19012 28494
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 18984 27674 19012 27950
rect 18972 27668 19024 27674
rect 18972 27610 19024 27616
rect 18892 27526 19012 27554
rect 18878 27024 18934 27033
rect 18878 26959 18934 26968
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18800 26518 18828 26726
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18892 26450 18920 26959
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 18786 25528 18842 25537
rect 18984 25514 19012 27526
rect 19076 27305 19104 28494
rect 19338 28455 19394 28464
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19168 27849 19196 28358
rect 19352 28082 19380 28455
rect 19423 28416 19475 28422
rect 19536 28404 19564 29260
rect 19616 29242 19668 29248
rect 19628 29102 19656 29242
rect 19996 29170 20024 31282
rect 20076 30592 20128 30598
rect 20180 30569 20208 31311
rect 20076 30534 20128 30540
rect 20166 30560 20222 30569
rect 20088 30054 20116 30534
rect 20166 30495 20222 30504
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20166 29472 20222 29481
rect 20088 29430 20166 29458
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19800 28688 19852 28694
rect 19892 28688 19944 28694
rect 19800 28630 19852 28636
rect 19890 28656 19892 28665
rect 19944 28656 19946 28665
rect 20088 28642 20116 29430
rect 20166 29407 20222 29416
rect 20168 28756 20220 28762
rect 20168 28698 20220 28704
rect 20180 28665 20208 28698
rect 19812 28529 19840 28630
rect 19890 28591 19946 28600
rect 19996 28614 20116 28642
rect 20166 28656 20222 28665
rect 19798 28520 19854 28529
rect 19798 28455 19854 28464
rect 19423 28358 19475 28364
rect 19511 28376 19564 28404
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19154 27840 19210 27849
rect 19154 27775 19210 27784
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19248 27328 19300 27334
rect 19062 27296 19118 27305
rect 19248 27270 19300 27276
rect 19062 27231 19118 27240
rect 19260 26761 19288 27270
rect 19246 26752 19302 26761
rect 19246 26687 19302 26696
rect 19156 26444 19208 26450
rect 19156 26386 19208 26392
rect 19062 26208 19118 26217
rect 19062 26143 19118 26152
rect 19076 25906 19104 26143
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 18842 25486 19012 25514
rect 18786 25463 18842 25472
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18800 24410 18828 24754
rect 18984 24721 19012 25366
rect 19076 24750 19104 25842
rect 19168 25702 19196 26386
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19064 24744 19116 24750
rect 18970 24712 19026 24721
rect 19064 24686 19116 24692
rect 18970 24647 19026 24656
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18800 23118 18828 24346
rect 18892 24206 18920 24550
rect 19062 24440 19118 24449
rect 19062 24375 19118 24384
rect 18972 24336 19024 24342
rect 18972 24278 19024 24284
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18892 23526 18920 24142
rect 18984 23730 19012 24278
rect 19076 24206 19104 24375
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19062 24032 19118 24041
rect 19062 23967 19118 23976
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18786 22944 18842 22953
rect 18786 22879 18842 22888
rect 18800 22624 18828 22879
rect 18892 22817 18920 23462
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 18878 22808 18934 22817
rect 18878 22743 18934 22752
rect 18984 22642 19012 23258
rect 19076 22778 19104 23967
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18972 22636 19024 22642
rect 18800 22596 18920 22624
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18616 21916 18736 21944
rect 18510 21720 18566 21729
rect 18708 21672 18736 21916
rect 18510 21655 18566 21664
rect 18524 21350 18552 21655
rect 18616 21644 18736 21672
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18512 21072 18564 21078
rect 18616 21060 18644 21644
rect 18800 21554 18828 22374
rect 18892 22030 18920 22596
rect 18972 22578 19024 22584
rect 18970 22400 19026 22409
rect 19076 22386 19104 22714
rect 19026 22358 19104 22386
rect 18970 22335 19026 22344
rect 18970 22264 19026 22273
rect 18970 22199 19026 22208
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18708 21146 18736 21490
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18564 21032 18644 21060
rect 18512 21014 18564 21020
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18418 20632 18474 20641
rect 18418 20567 18420 20576
rect 18472 20567 18474 20576
rect 18420 20538 18472 20544
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18326 19952 18382 19961
rect 18248 19910 18326 19938
rect 18326 19887 18382 19896
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 19310 18276 19654
rect 18340 19378 18368 19790
rect 18432 19718 18460 20402
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18050 19207 18106 19216
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18248 18766 18276 19246
rect 18340 18766 18368 19314
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18432 19009 18460 19246
rect 18418 19000 18474 19009
rect 18418 18935 18474 18944
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 17972 18426 18000 18702
rect 18340 18426 18368 18702
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18432 18601 18460 18634
rect 18418 18592 18474 18601
rect 18418 18527 18474 18536
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 17590 18255 17646 18264
rect 17684 18284 17736 18290
rect 17500 18226 17552 18232
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17604 18154 17632 18255
rect 17684 18226 17736 18232
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17406 18048 17462 18057
rect 17406 17983 17462 17992
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 17377 17356 17614
rect 17314 17368 17370 17377
rect 17314 17303 17370 17312
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16776 16250 16804 16730
rect 17328 16726 17356 17303
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 17420 16114 17448 17983
rect 17592 17808 17644 17814
rect 17590 17776 17592 17785
rect 17644 17776 17646 17785
rect 17590 17711 17646 17720
rect 17696 17678 17724 18226
rect 17972 17882 18000 18362
rect 18052 18284 18104 18290
rect 18524 18272 18552 21014
rect 18788 20936 18840 20942
rect 18694 20904 18750 20913
rect 18604 20868 18656 20874
rect 18788 20878 18840 20884
rect 18694 20839 18750 20848
rect 18604 20810 18656 20816
rect 18616 20058 18644 20810
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18616 19689 18644 19858
rect 18602 19680 18658 19689
rect 18602 19615 18658 19624
rect 18616 18834 18644 19615
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18104 18244 18552 18272
rect 18052 18226 18104 18232
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18064 17746 18092 18090
rect 18432 17746 18460 18244
rect 18708 18170 18736 20839
rect 18800 20505 18828 20878
rect 18892 20602 18920 21966
rect 18984 21865 19012 22199
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18970 21856 19026 21865
rect 18970 21791 19026 21800
rect 18970 21720 19026 21729
rect 18970 21655 19026 21664
rect 18984 21554 19012 21655
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 19076 21434 19104 21966
rect 19168 21962 19196 25638
rect 19260 24954 19288 25706
rect 19352 25294 19380 27610
rect 19444 27538 19472 28358
rect 19511 28200 19539 28376
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19511 28172 19564 28200
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19432 27328 19484 27334
rect 19536 27316 19564 28172
rect 19800 28144 19852 28150
rect 19800 28086 19852 28092
rect 19812 27441 19840 28086
rect 19798 27432 19854 27441
rect 19798 27367 19854 27376
rect 19484 27288 19564 27316
rect 19432 27270 19484 27276
rect 19444 27112 19472 27270
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27112 20024 28614
rect 20166 28591 20222 28600
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20088 27674 20116 28494
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19444 27084 19656 27112
rect 19432 26784 19484 26790
rect 19628 26761 19656 27084
rect 19720 27084 20024 27112
rect 19432 26726 19484 26732
rect 19614 26752 19670 26761
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19248 24948 19300 24954
rect 19444 24936 19472 26726
rect 19614 26687 19670 26696
rect 19720 26228 19748 27084
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19904 26364 19932 26726
rect 20088 26586 20116 27406
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19965 26376 20017 26382
rect 19904 26336 19965 26364
rect 20076 26376 20128 26382
rect 20017 26324 20024 26364
rect 19965 26318 20024 26324
rect 20076 26318 20128 26324
rect 19511 26200 19748 26228
rect 19511 26024 19539 26200
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 26042 20024 26318
rect 20088 26042 20116 26318
rect 19984 26036 20036 26042
rect 19511 25996 19564 26024
rect 19536 25498 19564 25996
rect 19984 25978 20036 25984
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19904 25430 19932 25638
rect 20180 25498 20208 28494
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 19892 25424 19944 25430
rect 19798 25392 19854 25401
rect 19892 25366 19944 25372
rect 19798 25327 19854 25336
rect 19812 25158 19840 25327
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 19800 25152 19852 25158
rect 19800 25094 19852 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19444 24908 19656 24936
rect 19248 24890 19300 24896
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19260 23730 19288 24754
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19352 24041 19380 24686
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19444 24206 19472 24618
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19338 24032 19394 24041
rect 19338 23967 19394 23976
rect 19444 23905 19472 24142
rect 19628 24052 19656 24908
rect 19800 24744 19852 24750
rect 19706 24712 19762 24721
rect 19800 24686 19852 24692
rect 19706 24647 19762 24656
rect 19720 24206 19748 24647
rect 19812 24206 19840 24686
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19904 24410 19932 24550
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19996 24138 20024 25230
rect 20076 25152 20128 25158
rect 20180 25129 20208 25230
rect 20076 25094 20128 25100
rect 20166 25120 20222 25129
rect 20088 24993 20116 25094
rect 20166 25055 20222 25064
rect 20074 24984 20130 24993
rect 20074 24919 20130 24928
rect 20088 24818 20116 24919
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24342 20116 24754
rect 20272 24682 20300 31690
rect 20364 30802 20392 32166
rect 20548 31754 20576 32388
rect 20640 32366 20668 34546
rect 21008 34406 21036 35158
rect 21376 35086 21404 37742
rect 21560 37670 21588 38422
rect 21638 38383 21694 38392
rect 21548 37664 21600 37670
rect 21548 37606 21600 37612
rect 21560 37330 21588 37606
rect 21548 37324 21600 37330
rect 21548 37266 21600 37272
rect 21652 36854 21680 38383
rect 21836 37806 21864 38830
rect 21928 38593 21956 38898
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 21914 38584 21970 38593
rect 21914 38519 21970 38528
rect 21916 38344 21968 38350
rect 22112 38332 22140 38694
rect 22296 38418 22324 39324
rect 22284 38412 22336 38418
rect 22284 38354 22336 38360
rect 21968 38304 22140 38332
rect 22192 38344 22244 38350
rect 21916 38286 21968 38292
rect 22192 38286 22244 38292
rect 22204 37856 22232 38286
rect 22388 38010 22416 39578
rect 23204 39296 23256 39302
rect 23204 39238 23256 39244
rect 23216 38758 23244 39238
rect 23204 38752 23256 38758
rect 23204 38694 23256 38700
rect 23216 38350 23244 38694
rect 23308 38486 23336 39782
rect 23388 39296 23440 39302
rect 23388 39238 23440 39244
rect 23400 38894 23428 39238
rect 23492 39030 23520 39918
rect 23676 39846 23704 40530
rect 23952 40050 23980 42026
rect 24492 42016 24544 42022
rect 24492 41958 24544 41964
rect 27344 42016 27396 42022
rect 27344 41958 27396 41964
rect 27896 42016 27948 42022
rect 27896 41958 27948 41964
rect 29092 42016 29144 42022
rect 29092 41958 29144 41964
rect 31024 42016 31076 42022
rect 31024 41958 31076 41964
rect 31484 42016 31536 42022
rect 31484 41958 31536 41964
rect 32680 42016 32732 42022
rect 32680 41958 32732 41964
rect 32772 42016 32824 42022
rect 32772 41958 32824 41964
rect 36452 42016 36504 42022
rect 36452 41958 36504 41964
rect 37648 42016 37700 42022
rect 37648 41958 37700 41964
rect 24504 41414 24532 41958
rect 27356 41414 27384 41958
rect 24504 41386 24624 41414
rect 27356 41386 27476 41414
rect 24596 40526 24624 41386
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 25056 40594 25084 40870
rect 25044 40588 25096 40594
rect 25044 40530 25096 40536
rect 27448 40526 27476 41386
rect 27804 41064 27856 41070
rect 27804 41006 27856 41012
rect 27712 40996 27764 41002
rect 27712 40938 27764 40944
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 27436 40520 27488 40526
rect 27436 40462 27488 40468
rect 24216 40452 24268 40458
rect 24216 40394 24268 40400
rect 26240 40452 26292 40458
rect 26240 40394 26292 40400
rect 24228 40118 24256 40394
rect 24768 40384 24820 40390
rect 24768 40326 24820 40332
rect 24780 40118 24808 40326
rect 24216 40112 24268 40118
rect 24216 40054 24268 40060
rect 24768 40112 24820 40118
rect 24768 40054 24820 40060
rect 23940 40044 23992 40050
rect 23940 39986 23992 39992
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 24124 39840 24176 39846
rect 24124 39782 24176 39788
rect 23480 39024 23532 39030
rect 23480 38966 23532 38972
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23480 38752 23532 38758
rect 23480 38694 23532 38700
rect 23296 38480 23348 38486
rect 23296 38422 23348 38428
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22560 37868 22612 37874
rect 22204 37828 22324 37856
rect 21824 37800 21876 37806
rect 21824 37742 21876 37748
rect 22100 37800 22152 37806
rect 22100 37742 22152 37748
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 21640 36848 21692 36854
rect 21640 36790 21692 36796
rect 21456 36712 21508 36718
rect 21456 36654 21508 36660
rect 21468 36174 21496 36654
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21468 35698 21496 36110
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21088 35080 21140 35086
rect 21364 35080 21416 35086
rect 21140 35040 21220 35068
rect 21088 35022 21140 35028
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20996 34400 21048 34406
rect 20996 34342 21048 34348
rect 20732 32570 20760 34342
rect 20812 33652 20864 33658
rect 20812 33594 20864 33600
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20824 32434 20852 33594
rect 21100 33522 21128 34886
rect 21192 33833 21220 35040
rect 21364 35022 21416 35028
rect 21270 34640 21326 34649
rect 21270 34575 21272 34584
rect 21324 34575 21326 34584
rect 21272 34546 21324 34552
rect 21272 34400 21324 34406
rect 21272 34342 21324 34348
rect 21178 33824 21234 33833
rect 21178 33759 21234 33768
rect 21088 33516 21140 33522
rect 21140 33476 21220 33504
rect 21088 33458 21140 33464
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20916 32910 20944 33390
rect 20904 32904 20956 32910
rect 20904 32846 20956 32852
rect 20916 32502 20944 32846
rect 20904 32496 20956 32502
rect 20904 32438 20956 32444
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20916 31890 20944 32438
rect 20996 32360 21048 32366
rect 20996 32302 21048 32308
rect 21008 31958 21036 32302
rect 20996 31952 21048 31958
rect 20996 31894 21048 31900
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20536 31476 20588 31482
rect 20536 31418 20588 31424
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 20456 30870 20484 31214
rect 20548 31142 20576 31418
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20444 30864 20496 30870
rect 20444 30806 20496 30812
rect 20352 30796 20404 30802
rect 20352 30738 20404 30744
rect 20364 30326 20392 30738
rect 20640 30682 20668 31282
rect 20812 31204 20864 31210
rect 20812 31146 20864 31152
rect 20718 30832 20774 30841
rect 20718 30767 20720 30776
rect 20772 30767 20774 30776
rect 20720 30738 20772 30744
rect 20456 30654 20668 30682
rect 20720 30660 20772 30666
rect 20456 30598 20484 30654
rect 20720 30602 20772 30608
rect 20444 30592 20496 30598
rect 20536 30592 20588 30598
rect 20444 30534 20496 30540
rect 20534 30560 20536 30569
rect 20588 30560 20590 30569
rect 20534 30495 20590 30504
rect 20732 30394 20760 30602
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20352 30320 20404 30326
rect 20444 30320 20496 30326
rect 20352 30262 20404 30268
rect 20442 30288 20444 30297
rect 20824 30297 20852 31146
rect 20916 30802 20944 31826
rect 21088 31680 21140 31686
rect 21088 31622 21140 31628
rect 21100 31414 21128 31622
rect 21192 31414 21220 33476
rect 21284 32230 21312 34342
rect 21376 33998 21404 35022
rect 21652 33998 21680 36790
rect 21744 36038 21772 37062
rect 22112 36242 22140 37742
rect 22192 37732 22244 37738
rect 22192 37674 22244 37680
rect 22204 36922 22232 37674
rect 22296 37262 22324 37828
rect 22560 37810 22612 37816
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22296 37126 22324 37198
rect 22468 37188 22520 37194
rect 22468 37130 22520 37136
rect 22284 37120 22336 37126
rect 22284 37062 22336 37068
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 22480 36378 22508 37130
rect 22572 37126 22600 37810
rect 23216 37210 23244 38286
rect 23308 37330 23336 38422
rect 23492 38350 23520 38694
rect 23676 38418 23704 39782
rect 24136 39370 24164 39782
rect 24124 39364 24176 39370
rect 24124 39306 24176 39312
rect 24228 38894 24256 40054
rect 24492 39840 24544 39846
rect 24492 39782 24544 39788
rect 25320 39840 25372 39846
rect 25320 39782 25372 39788
rect 24504 39438 24532 39782
rect 25332 39438 25360 39782
rect 26252 39642 26280 40394
rect 26608 40384 26660 40390
rect 26608 40326 26660 40332
rect 26700 40384 26752 40390
rect 26700 40326 26752 40332
rect 27160 40384 27212 40390
rect 27160 40326 27212 40332
rect 27620 40384 27672 40390
rect 27620 40326 27672 40332
rect 26620 40050 26648 40326
rect 26712 40118 26740 40326
rect 26700 40112 26752 40118
rect 26700 40054 26752 40060
rect 26608 40044 26660 40050
rect 26608 39986 26660 39992
rect 26240 39636 26292 39642
rect 26240 39578 26292 39584
rect 26332 39636 26384 39642
rect 26332 39578 26384 39584
rect 25964 39500 26016 39506
rect 25964 39442 26016 39448
rect 24400 39432 24452 39438
rect 24400 39374 24452 39380
rect 24492 39432 24544 39438
rect 24492 39374 24544 39380
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24320 39030 24348 39238
rect 24412 39098 24440 39374
rect 24400 39092 24452 39098
rect 24400 39034 24452 39040
rect 24504 39030 24532 39374
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24308 39024 24360 39030
rect 24308 38966 24360 38972
rect 24492 39024 24544 39030
rect 24492 38966 24544 38972
rect 23940 38888 23992 38894
rect 23940 38830 23992 38836
rect 24216 38888 24268 38894
rect 24216 38830 24268 38836
rect 23664 38412 23716 38418
rect 23664 38354 23716 38360
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23756 37664 23808 37670
rect 23756 37606 23808 37612
rect 23296 37324 23348 37330
rect 23296 37266 23348 37272
rect 22836 37188 22888 37194
rect 23216 37182 23428 37210
rect 22836 37130 22888 37136
rect 22560 37120 22612 37126
rect 22560 37062 22612 37068
rect 22848 36922 22876 37130
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 23400 37074 23428 37182
rect 23572 37120 23624 37126
rect 22836 36916 22888 36922
rect 22836 36858 22888 36864
rect 23124 36786 23152 37062
rect 23400 37046 23520 37074
rect 23572 37062 23624 37068
rect 23112 36780 23164 36786
rect 23112 36722 23164 36728
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23124 36689 23152 36722
rect 23110 36680 23166 36689
rect 23110 36615 23166 36624
rect 22468 36372 22520 36378
rect 22468 36314 22520 36320
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 21824 36168 21876 36174
rect 21824 36110 21876 36116
rect 21732 36032 21784 36038
rect 21732 35974 21784 35980
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21364 33856 21416 33862
rect 21364 33798 21416 33804
rect 21376 33658 21404 33798
rect 21364 33652 21416 33658
rect 21364 33594 21416 33600
rect 21548 33516 21600 33522
rect 21548 33458 21600 33464
rect 21560 33289 21588 33458
rect 21546 33280 21602 33289
rect 21546 33215 21602 33224
rect 21362 33008 21418 33017
rect 21362 32943 21418 32952
rect 21272 32224 21324 32230
rect 21272 32166 21324 32172
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21088 31408 21140 31414
rect 21088 31350 21140 31356
rect 21180 31408 21232 31414
rect 21180 31350 21232 31356
rect 20996 31272 21048 31278
rect 20996 31214 21048 31220
rect 20904 30796 20956 30802
rect 20904 30738 20956 30744
rect 21008 30682 21036 31214
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 20916 30654 21036 30682
rect 20916 30598 20944 30654
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20496 30288 20498 30297
rect 20364 29617 20392 30262
rect 20442 30223 20498 30232
rect 20810 30288 20866 30297
rect 20810 30223 20866 30232
rect 20812 30184 20864 30190
rect 20732 30144 20812 30172
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20350 29608 20406 29617
rect 20350 29543 20406 29552
rect 20548 29170 20576 29650
rect 20732 29306 20760 30144
rect 20812 30126 20864 30132
rect 20812 29572 20864 29578
rect 20812 29514 20864 29520
rect 20824 29306 20852 29514
rect 20916 29510 20944 30534
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 20996 30116 21048 30122
rect 20996 30058 21048 30064
rect 21008 29646 21036 30058
rect 21100 29850 21128 30194
rect 21088 29844 21140 29850
rect 21088 29786 21140 29792
rect 21192 29646 21220 31078
rect 21284 30433 21312 31690
rect 21376 31249 21404 32943
rect 21456 31680 21508 31686
rect 21456 31622 21508 31628
rect 21548 31680 21600 31686
rect 21548 31622 21600 31628
rect 21362 31240 21418 31249
rect 21362 31175 21418 31184
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21270 30424 21326 30433
rect 21270 30359 21326 30368
rect 21376 30258 21404 31078
rect 21364 30252 21416 30258
rect 21364 30194 21416 30200
rect 21362 30152 21418 30161
rect 21468 30138 21496 31622
rect 21560 30161 21588 31622
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21652 30190 21680 31078
rect 21640 30184 21692 30190
rect 21418 30110 21496 30138
rect 21362 30087 21418 30096
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 21008 29306 21036 29582
rect 21468 29481 21496 30110
rect 21546 30152 21602 30161
rect 21640 30126 21692 30132
rect 21546 30087 21602 30096
rect 21744 29753 21772 35974
rect 21836 35834 21864 36110
rect 21824 35828 21876 35834
rect 21824 35770 21876 35776
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 22008 35012 22060 35018
rect 22008 34954 22060 34960
rect 21836 34746 21864 34954
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 21824 34604 21876 34610
rect 21824 34546 21876 34552
rect 21836 33114 21864 34546
rect 21916 33924 21968 33930
rect 21916 33866 21968 33872
rect 21928 33454 21956 33866
rect 22020 33590 22048 34954
rect 22204 34746 22232 35090
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22652 34944 22704 34950
rect 22652 34886 22704 34892
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22296 34610 22324 34886
rect 22664 34746 22692 34886
rect 22652 34740 22704 34746
rect 22652 34682 22704 34688
rect 23020 34740 23072 34746
rect 23020 34682 23072 34688
rect 23032 34649 23060 34682
rect 22374 34640 22430 34649
rect 22284 34604 22336 34610
rect 23018 34640 23074 34649
rect 22430 34598 22508 34626
rect 22374 34575 22430 34584
rect 22284 34546 22336 34552
rect 22376 34536 22428 34542
rect 22376 34478 22428 34484
rect 22388 34202 22416 34478
rect 22376 34196 22428 34202
rect 22376 34138 22428 34144
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 22008 33584 22060 33590
rect 22008 33526 22060 33532
rect 21916 33448 21968 33454
rect 21916 33390 21968 33396
rect 21824 33108 21876 33114
rect 21824 33050 21876 33056
rect 21836 31346 21864 33050
rect 22020 32230 22048 33526
rect 22204 33114 22232 34002
rect 22388 33658 22416 34138
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22388 32978 22416 33254
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22480 32570 22508 34598
rect 23018 34575 23074 34584
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 22652 34128 22704 34134
rect 22652 34070 22704 34076
rect 22664 33862 22692 34070
rect 22744 33992 22796 33998
rect 22744 33934 22796 33940
rect 22756 33862 22784 33934
rect 22928 33924 22980 33930
rect 22848 33884 22928 33912
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 22020 31770 22048 32166
rect 22112 31890 22140 32302
rect 22100 31884 22152 31890
rect 22100 31826 22152 31832
rect 22020 31742 22140 31770
rect 21916 31680 21968 31686
rect 21916 31622 21968 31628
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21928 31226 21956 31622
rect 21836 31198 21956 31226
rect 21836 30569 21864 31198
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 21822 30560 21878 30569
rect 21822 30495 21878 30504
rect 22020 30394 22048 30670
rect 22008 30388 22060 30394
rect 22008 30330 22060 30336
rect 21730 29744 21786 29753
rect 21730 29679 21786 29688
rect 21178 29472 21234 29481
rect 21178 29407 21234 29416
rect 21454 29472 21510 29481
rect 21454 29407 21510 29416
rect 21192 29306 21220 29407
rect 21454 29336 21510 29345
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 21180 29300 21232 29306
rect 21454 29271 21510 29280
rect 21180 29242 21232 29248
rect 21468 29170 21496 29271
rect 21744 29170 21772 29679
rect 22112 29345 22140 31742
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 22744 31340 22796 31346
rect 22744 31282 22796 31288
rect 22204 30122 22232 31282
rect 22560 31204 22612 31210
rect 22756 31192 22784 31282
rect 22612 31164 22784 31192
rect 22560 31146 22612 31152
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 22192 30116 22244 30122
rect 22192 30058 22244 30064
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22204 29646 22232 29786
rect 22296 29714 22324 31078
rect 22374 30968 22430 30977
rect 22374 30903 22430 30912
rect 22468 30932 22520 30938
rect 22388 30190 22416 30903
rect 22468 30874 22520 30880
rect 22480 30258 22508 30874
rect 22650 30696 22706 30705
rect 22650 30631 22706 30640
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22480 29782 22508 30194
rect 22664 30054 22692 30631
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22468 29776 22520 29782
rect 22468 29718 22520 29724
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22098 29336 22154 29345
rect 22098 29271 22154 29280
rect 22204 29220 22232 29582
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22204 29192 22324 29220
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 20442 29064 20498 29073
rect 20442 28999 20498 29008
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20364 27674 20392 28494
rect 20456 28422 20484 28999
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20548 28098 20576 28902
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20824 28121 20852 28562
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20916 28150 20944 28358
rect 20904 28144 20956 28150
rect 20456 28082 20576 28098
rect 20444 28076 20576 28082
rect 20496 28070 20576 28076
rect 20810 28112 20866 28121
rect 20904 28086 20956 28092
rect 20810 28047 20866 28056
rect 20444 28018 20496 28024
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 21088 27872 21140 27878
rect 21088 27814 21140 27820
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20364 26994 20392 27610
rect 20732 27538 20760 27814
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20732 27130 20760 27270
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 20548 26790 20576 26862
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20548 26489 20576 26726
rect 20640 26586 20668 27066
rect 20824 26926 20852 27814
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20534 26480 20590 26489
rect 20534 26415 20590 26424
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20364 25498 20392 26318
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20536 26240 20588 26246
rect 20536 26182 20588 26188
rect 20352 25492 20404 25498
rect 20456 25480 20484 26182
rect 20548 26042 20576 26182
rect 20536 26036 20588 26042
rect 20536 25978 20588 25984
rect 20640 25702 20668 26318
rect 20732 26314 20760 26726
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20718 25936 20774 25945
rect 20718 25871 20720 25880
rect 20772 25871 20774 25880
rect 20720 25842 20772 25848
rect 20824 25838 20852 26454
rect 20916 26024 20944 26930
rect 21008 26314 21036 27542
rect 21100 27470 21128 27814
rect 21192 27606 21220 29106
rect 21272 27872 21324 27878
rect 21270 27840 21272 27849
rect 21324 27840 21326 27849
rect 21270 27775 21326 27784
rect 21180 27600 21232 27606
rect 21180 27542 21232 27548
rect 21284 27470 21312 27775
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21192 26450 21220 26862
rect 21180 26444 21232 26450
rect 21180 26386 21232 26392
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 20916 25996 21036 26024
rect 20902 25936 20958 25945
rect 21008 25906 21036 25996
rect 20902 25871 20958 25880
rect 20996 25900 21048 25906
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20628 25696 20680 25702
rect 20916 25673 20944 25871
rect 20996 25842 21048 25848
rect 21100 25702 21128 26182
rect 21088 25696 21140 25702
rect 20628 25638 20680 25644
rect 20902 25664 20958 25673
rect 21088 25638 21140 25644
rect 20902 25599 20958 25608
rect 20536 25492 20588 25498
rect 20456 25452 20536 25480
rect 20352 25434 20404 25440
rect 21192 25480 21220 26386
rect 21272 25492 21324 25498
rect 21192 25452 21272 25480
rect 20536 25434 20588 25440
rect 21272 25434 21324 25440
rect 20364 25378 20392 25434
rect 20626 25392 20682 25401
rect 20364 25350 20626 25378
rect 20626 25327 20682 25336
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 20350 25120 20406 25129
rect 20350 25055 20406 25064
rect 20364 24818 20392 25055
rect 20456 24993 20484 25230
rect 20720 25220 20772 25226
rect 20720 25162 20772 25168
rect 20442 24984 20498 24993
rect 20442 24919 20498 24928
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20260 24676 20312 24682
rect 20444 24676 20496 24682
rect 20260 24618 20312 24624
rect 20364 24636 20444 24664
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20180 24342 20208 24550
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 20168 24336 20220 24342
rect 20168 24278 20220 24284
rect 20260 24268 20312 24274
rect 20260 24210 20312 24216
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19800 24064 19852 24070
rect 19628 24024 19800 24052
rect 20076 24064 20128 24070
rect 19800 24006 19852 24012
rect 19982 24032 20038 24041
rect 20076 24006 20128 24012
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19574 23964 19882 23973
rect 19982 23967 20038 23976
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19430 23896 19486 23905
rect 19574 23899 19882 23908
rect 19352 23854 19430 23882
rect 19352 23730 19380 23854
rect 19430 23831 19486 23840
rect 19800 23860 19852 23866
rect 19996 23848 20024 23967
rect 19852 23820 20024 23848
rect 19800 23802 19852 23808
rect 20088 23798 20116 24006
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19260 23322 19288 23666
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19524 23588 19576 23594
rect 19444 23548 19524 23576
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19340 23112 19392 23118
rect 19260 23072 19340 23100
rect 19260 22778 19288 23072
rect 19444 23066 19472 23548
rect 19524 23530 19576 23536
rect 19890 23352 19946 23361
rect 19890 23287 19892 23296
rect 19944 23287 19946 23296
rect 19892 23258 19944 23264
rect 19616 23248 19668 23254
rect 19996 23202 20024 23598
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 20088 23322 20116 23530
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19616 23190 19668 23196
rect 19340 23054 19392 23060
rect 19435 23038 19472 23066
rect 19435 22964 19463 23038
rect 19628 22964 19656 23190
rect 19904 23174 20024 23202
rect 19904 23118 19932 23174
rect 19892 23112 19944 23118
rect 20088 23100 20116 23258
rect 20180 23118 20208 24006
rect 20272 23594 20300 24210
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20364 23526 20392 24636
rect 20444 24618 20496 24624
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20456 23730 20484 24074
rect 20548 23730 20576 24754
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20640 23866 20668 24618
rect 20732 23866 20760 25162
rect 20824 24954 20852 25230
rect 20812 24948 20864 24954
rect 20812 24890 20864 24896
rect 21008 24886 21036 25230
rect 21376 24886 21404 26386
rect 21468 25702 21496 29106
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21928 28082 21956 28358
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21560 26081 21588 26318
rect 21546 26072 21602 26081
rect 21652 26042 21680 27270
rect 21744 26450 21772 27610
rect 22190 27432 22246 27441
rect 22190 27367 22192 27376
rect 22244 27367 22246 27376
rect 22192 27338 22244 27344
rect 22190 27160 22246 27169
rect 22296 27146 22324 29192
rect 22480 28082 22508 29446
rect 22572 29209 22600 29446
rect 22558 29200 22614 29209
rect 22664 29186 22692 29990
rect 22756 29850 22784 30534
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22756 29306 22784 29582
rect 22744 29300 22796 29306
rect 22744 29242 22796 29248
rect 22664 29170 22784 29186
rect 22664 29164 22796 29170
rect 22664 29158 22744 29164
rect 22558 29135 22614 29144
rect 22744 29106 22796 29112
rect 22652 28960 22704 28966
rect 22650 28928 22652 28937
rect 22704 28928 22706 28937
rect 22650 28863 22706 28872
rect 22664 28082 22692 28863
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22246 27118 22324 27146
rect 22190 27095 22246 27104
rect 22098 27024 22154 27033
rect 22098 26959 22100 26968
rect 22152 26959 22154 26968
rect 22284 26988 22336 26994
rect 22100 26930 22152 26936
rect 22284 26930 22336 26936
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 21546 26007 21602 26016
rect 21640 26036 21692 26042
rect 21640 25978 21692 25984
rect 21652 25838 21680 25978
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 22020 25498 22048 26318
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 22204 25294 22232 26726
rect 22296 26586 22324 26930
rect 22664 26761 22692 26930
rect 22650 26752 22706 26761
rect 22650 26687 22706 26696
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22466 26208 22522 26217
rect 22466 26143 22522 26152
rect 22480 25906 22508 26143
rect 22468 25900 22520 25906
rect 22468 25842 22520 25848
rect 22376 25764 22428 25770
rect 22376 25706 22428 25712
rect 22388 25294 22416 25706
rect 21640 25288 21692 25294
rect 22100 25288 22152 25294
rect 21692 25248 21772 25276
rect 21640 25230 21692 25236
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 21364 24880 21416 24886
rect 21364 24822 21416 24828
rect 21468 24818 21496 25162
rect 21546 24984 21602 24993
rect 21546 24919 21548 24928
rect 21600 24919 21602 24928
rect 21548 24890 21600 24896
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 20824 24206 20852 24754
rect 21364 24744 21416 24750
rect 20902 24712 20958 24721
rect 20902 24647 20904 24656
rect 20956 24647 20958 24656
rect 21270 24712 21326 24721
rect 21364 24686 21416 24692
rect 21270 24647 21326 24656
rect 20904 24618 20956 24624
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21100 24206 21128 24550
rect 21178 24440 21234 24449
rect 21178 24375 21234 24384
rect 21192 24206 21220 24375
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20996 24064 21048 24070
rect 21100 24041 21128 24142
rect 20996 24006 21048 24012
rect 21086 24032 21142 24041
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20456 23254 20484 23666
rect 20444 23248 20496 23254
rect 20444 23190 20496 23196
rect 19892 23054 19944 23060
rect 19996 23072 20116 23100
rect 20168 23112 20220 23118
rect 19435 22936 19472 22964
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19444 22642 19472 22936
rect 19511 22936 19656 22964
rect 19511 22778 19539 22936
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19511 22772 19576 22778
rect 19511 22732 19524 22772
rect 19996 22760 20024 23072
rect 20220 23072 20392 23100
rect 20168 23054 20220 23060
rect 20258 22944 20314 22953
rect 20258 22879 20314 22888
rect 19524 22714 19576 22720
rect 19904 22732 20024 22760
rect 20168 22772 20220 22778
rect 19616 22704 19668 22710
rect 19614 22672 19616 22681
rect 19668 22672 19670 22681
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19524 22636 19576 22642
rect 19614 22607 19670 22616
rect 19798 22672 19854 22681
rect 19904 22642 19932 22732
rect 20272 22760 20300 22879
rect 20220 22732 20300 22760
rect 20168 22714 20220 22720
rect 20364 22642 20392 23072
rect 20456 22642 20484 23190
rect 20548 23118 20576 23666
rect 20640 23118 20668 23802
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20732 23254 20760 23666
rect 20720 23248 20772 23254
rect 20720 23190 20772 23196
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 19798 22607 19854 22616
rect 19892 22636 19944 22642
rect 19524 22578 19576 22584
rect 19260 22545 19288 22578
rect 19246 22536 19302 22545
rect 19352 22522 19380 22578
rect 19352 22494 19472 22522
rect 19246 22471 19302 22480
rect 19444 22098 19472 22494
rect 19536 22234 19564 22578
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19156 21956 19208 21962
rect 19208 21916 19288 21944
rect 19156 21898 19208 21904
rect 19154 21856 19210 21865
rect 19154 21791 19210 21800
rect 19168 21554 19196 21791
rect 19260 21570 19288 21916
rect 19352 21690 19380 22034
rect 19340 21684 19392 21690
rect 19444 21672 19472 22034
rect 19628 21894 19656 22374
rect 19812 22098 19840 22607
rect 20352 22636 20404 22642
rect 19892 22578 19944 22584
rect 20272 22596 20352 22624
rect 19904 22114 19932 22578
rect 20272 22438 20300 22596
rect 20352 22578 20404 22584
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20548 22522 20576 22918
rect 20640 22817 20668 23054
rect 20626 22808 20682 22817
rect 20732 22778 20760 23190
rect 20916 23118 20944 24006
rect 21008 23662 21036 24006
rect 21086 23967 21142 23976
rect 21192 23905 21220 24142
rect 21178 23896 21234 23905
rect 21088 23860 21140 23866
rect 21284 23866 21312 24647
rect 21376 23866 21404 24686
rect 21468 24070 21496 24754
rect 21744 24410 21772 25248
rect 22100 25230 22152 25236
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22376 25288 22428 25294
rect 22468 25288 22520 25294
rect 22376 25230 22428 25236
rect 22466 25256 22468 25265
rect 22520 25256 22522 25265
rect 22112 25158 22140 25230
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22388 24886 22416 25230
rect 22466 25191 22522 25200
rect 21824 24880 21876 24886
rect 22376 24880 22428 24886
rect 21824 24822 21876 24828
rect 21914 24848 21970 24857
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21548 24200 21600 24206
rect 21546 24168 21548 24177
rect 21600 24168 21602 24177
rect 21546 24103 21602 24112
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21652 23866 21680 24346
rect 21178 23831 21234 23840
rect 21272 23860 21324 23866
rect 21088 23802 21140 23808
rect 21272 23802 21324 23808
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20626 22743 20682 22752
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20364 22494 20576 22522
rect 20260 22432 20312 22438
rect 20074 22400 20130 22409
rect 19996 22358 20074 22386
rect 19996 22234 20024 22358
rect 20260 22374 20312 22380
rect 20074 22335 20130 22344
rect 19984 22228 20036 22234
rect 20272 22216 20300 22374
rect 20364 22273 20392 22494
rect 20536 22432 20588 22438
rect 20534 22400 20536 22409
rect 20588 22400 20590 22409
rect 20534 22335 20590 22344
rect 19984 22170 20036 22176
rect 20088 22188 20300 22216
rect 20350 22264 20406 22273
rect 20640 22250 20668 22578
rect 20732 22522 20760 22714
rect 20732 22494 20852 22522
rect 20916 22506 20944 23054
rect 21100 22930 21128 23802
rect 21376 23594 21404 23802
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 23588 21416 23594
rect 21364 23530 21416 23536
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21008 22902 21128 22930
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20350 22199 20406 22208
rect 20456 22222 20668 22250
rect 19800 22092 19852 22098
rect 19904 22086 20024 22114
rect 19800 22034 19852 22040
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21672 20024 22086
rect 19444 21644 19656 21672
rect 19340 21626 19392 21632
rect 19156 21548 19208 21554
rect 19260 21542 19472 21570
rect 19628 21554 19656 21644
rect 19720 21644 20024 21672
rect 19156 21490 19208 21496
rect 18984 21406 19104 21434
rect 19156 21412 19208 21418
rect 18984 21026 19012 21406
rect 19156 21354 19208 21360
rect 18984 20998 19104 21026
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18984 20806 19012 20878
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18786 20496 18842 20505
rect 18786 20431 18842 20440
rect 18984 19990 19012 20742
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18970 19816 19026 19825
rect 18800 19514 18828 19790
rect 18970 19751 19026 19760
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18800 18766 18828 19314
rect 18892 19310 18920 19654
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18984 19174 19012 19751
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18786 18456 18842 18465
rect 18786 18391 18788 18400
rect 18840 18391 18842 18400
rect 18788 18362 18840 18368
rect 18616 18154 18736 18170
rect 18604 18148 18736 18154
rect 18656 18142 18736 18148
rect 18604 18090 18656 18096
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17882 18552 18022
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 17684 17672 17736 17678
rect 18432 17649 18460 17682
rect 18418 17640 18474 17649
rect 17684 17614 17736 17620
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 17338 17540 17478
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17512 16794 17540 17274
rect 17604 16794 17632 17546
rect 17696 17202 17724 17614
rect 18340 17598 18418 17626
rect 18340 17202 18368 17598
rect 18418 17575 18474 17584
rect 18524 17202 18552 17818
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 17696 16998 17724 17138
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 18340 16658 18368 17138
rect 18616 17134 18644 18090
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17814 18736 18022
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18892 17338 18920 18770
rect 19076 17882 19104 20998
rect 19168 20992 19196 21354
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19246 21176 19302 21185
rect 19246 21111 19302 21120
rect 19260 20992 19288 21111
rect 19168 20964 19288 20992
rect 19168 20058 19196 20964
rect 19352 20942 19380 21286
rect 19444 21010 19472 21542
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19628 21146 19656 21490
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19524 20800 19576 20806
rect 19720 20788 19748 21644
rect 20088 21570 20116 22188
rect 20456 22166 20484 22222
rect 20444 22160 20496 22166
rect 20166 22128 20222 22137
rect 20222 22086 20300 22114
rect 20444 22102 20496 22108
rect 20534 22128 20590 22137
rect 20166 22063 20222 22072
rect 20272 22030 20300 22086
rect 20732 22098 20760 22374
rect 20824 22166 20852 22494
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 21008 22386 21036 22902
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21100 22642 21128 22714
rect 21192 22642 21220 23054
rect 21284 22982 21312 23462
rect 21364 23316 21416 23322
rect 21468 23304 21496 23666
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21416 23276 21496 23304
rect 21364 23258 21416 23264
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21376 22710 21404 23258
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21560 22778 21588 23190
rect 21652 23118 21680 23530
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21364 22704 21416 22710
rect 21364 22646 21416 22652
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21364 22568 21416 22574
rect 21284 22528 21364 22556
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 20916 22358 21036 22386
rect 20812 22160 20864 22166
rect 20812 22102 20864 22108
rect 20534 22063 20590 22072
rect 20720 22092 20772 22098
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20442 21992 20498 22001
rect 20272 21729 20300 21966
rect 20442 21927 20498 21936
rect 20456 21894 20484 21927
rect 20444 21888 20496 21894
rect 20350 21856 20406 21865
rect 20444 21830 20496 21836
rect 20350 21791 20406 21800
rect 20258 21720 20314 21729
rect 20258 21655 20314 21664
rect 19904 21554 20116 21570
rect 19892 21548 20116 21554
rect 19944 21542 20116 21548
rect 19892 21490 19944 21496
rect 19800 21344 19852 21350
rect 19798 21312 19800 21321
rect 19892 21344 19944 21350
rect 19852 21312 19854 21321
rect 19892 21286 19944 21292
rect 19798 21247 19854 21256
rect 19904 21026 19932 21286
rect 19812 20998 19932 21026
rect 19982 21040 20038 21049
rect 19812 20806 19840 20998
rect 19982 20975 20038 20984
rect 19892 20936 19944 20942
rect 19890 20904 19892 20913
rect 19944 20904 19946 20913
rect 19890 20839 19946 20848
rect 19576 20760 19748 20788
rect 19800 20800 19852 20806
rect 19524 20742 19576 20748
rect 19800 20742 19852 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19430 20632 19486 20641
rect 19574 20635 19882 20644
rect 19486 20576 19932 20584
rect 19430 20567 19932 20576
rect 19444 20556 19932 20567
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19260 20233 19288 20402
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19246 20224 19302 20233
rect 19246 20159 19302 20168
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19340 19916 19392 19922
rect 19444 19904 19472 20334
rect 19392 19876 19472 19904
rect 19340 19858 19392 19864
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19168 19446 19196 19790
rect 19352 19514 19380 19858
rect 19524 19848 19576 19854
rect 19444 19808 19524 19836
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19156 19236 19208 19242
rect 19156 19178 19208 19184
rect 19168 18290 19196 19178
rect 19260 18834 19288 19450
rect 19352 19378 19380 19450
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19444 18358 19472 19808
rect 19524 19790 19576 19796
rect 19524 19712 19576 19718
rect 19511 19660 19524 19700
rect 19628 19700 19656 20402
rect 19720 19825 19748 20402
rect 19904 20398 19932 20556
rect 19996 20534 20024 20975
rect 20088 20806 20116 21542
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 20800 20128 20806
rect 20180 20777 20208 21422
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 21049 20300 21286
rect 20258 21040 20314 21049
rect 20258 20975 20314 20984
rect 20364 20942 20392 21791
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20076 20742 20128 20748
rect 20166 20768 20222 20777
rect 20166 20703 20222 20712
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19982 20360 20038 20369
rect 19812 20244 19840 20334
rect 20038 20318 20208 20346
rect 19982 20295 20038 20304
rect 19812 20216 20116 20244
rect 20088 19854 20116 20216
rect 20180 19990 20208 20318
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20076 19848 20128 19854
rect 19706 19816 19762 19825
rect 20076 19790 20128 19796
rect 19706 19751 19762 19760
rect 19576 19672 19656 19700
rect 19984 19712 20036 19718
rect 19511 19654 19576 19660
rect 19984 19654 20036 19660
rect 19511 19496 19539 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19511 19468 19564 19496
rect 19536 18698 19564 19468
rect 19892 19440 19944 19446
rect 19890 19408 19892 19417
rect 19944 19408 19946 19417
rect 19996 19378 20024 19654
rect 19890 19343 19946 19352
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19720 18873 19748 19178
rect 20088 19174 20116 19790
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19706 18864 19762 18873
rect 19706 18799 19762 18808
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19432 18352 19484 18358
rect 19352 18312 19432 18340
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16794 18644 17070
rect 18892 16794 18920 17274
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19168 16998 19196 17138
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18510 16552 18566 16561
rect 18510 16487 18566 16496
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15706 17172 15982
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 15016 15632 15068 15638
rect 15014 15600 15016 15609
rect 15568 15632 15620 15638
rect 15068 15600 15070 15609
rect 14740 15564 14792 15570
rect 15568 15574 15620 15580
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 15014 15535 15070 15544
rect 14740 15506 14792 15512
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14568 14278 14596 15302
rect 14752 15162 14780 15506
rect 15028 15162 15056 15535
rect 17420 15502 17448 15846
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17972 15434 18000 15846
rect 18524 15638 18552 16487
rect 19076 16114 19104 16594
rect 19168 16590 19196 16934
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 16114 19196 16526
rect 19260 16454 19288 17002
rect 19352 16454 19380 18312
rect 19432 18294 19484 18300
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19522 17912 19578 17921
rect 19522 17847 19578 17856
rect 19536 17678 19564 17847
rect 19720 17678 19748 18294
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19812 17678 19840 18022
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19260 15910 19288 16390
rect 19444 16250 19472 17546
rect 19904 17524 19932 18362
rect 19996 18290 20024 18906
rect 20088 18698 20116 19110
rect 20272 18970 20300 20810
rect 20350 20632 20406 20641
rect 20350 20567 20406 20576
rect 20364 20330 20392 20567
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20364 19281 20392 19722
rect 20350 19272 20406 19281
rect 20350 19207 20406 19216
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20364 18850 20392 19207
rect 20272 18834 20392 18850
rect 20260 18828 20392 18834
rect 20312 18822 20392 18828
rect 20260 18770 20312 18776
rect 20352 18760 20404 18766
rect 20456 18748 20484 21558
rect 20548 21554 20576 22063
rect 20720 22034 20772 22040
rect 20824 21622 20852 22102
rect 20916 22030 20944 22358
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 21008 21162 21036 22170
rect 21100 21962 21128 22442
rect 21178 22128 21234 22137
rect 21178 22063 21180 22072
rect 21232 22063 21234 22072
rect 21180 22034 21232 22040
rect 21284 22030 21312 22528
rect 21364 22510 21416 22516
rect 21364 22160 21416 22166
rect 21364 22102 21416 22108
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21100 21690 21128 21898
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 21086 21584 21142 21593
rect 21086 21519 21088 21528
rect 21140 21519 21142 21528
rect 21088 21490 21140 21496
rect 21008 21134 21128 21162
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20628 20936 20680 20942
rect 20680 20896 20760 20924
rect 20628 20878 20680 20884
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 19854 20576 20402
rect 20640 19922 20668 20742
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 19378 20576 19790
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20404 18720 20484 18748
rect 20352 18702 20404 18708
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 17678 20024 18226
rect 20088 17678 20116 18634
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 18154 20208 18566
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20166 17640 20222 17649
rect 20166 17575 20222 17584
rect 20180 17524 20208 17575
rect 19904 17496 20024 17524
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19890 17232 19946 17241
rect 19800 17196 19852 17202
rect 19890 17167 19892 17176
rect 19800 17138 19852 17144
rect 19944 17167 19946 17176
rect 19892 17138 19944 17144
rect 19812 16726 19840 17138
rect 19904 16794 19932 17138
rect 19996 16998 20024 17496
rect 20088 17496 20208 17524
rect 20088 17202 20116 17496
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 20272 16590 20300 16934
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20364 16250 20392 18702
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20456 18426 20484 18566
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20640 18290 20668 19382
rect 20732 19334 20760 20896
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20824 20641 20852 20742
rect 20810 20632 20866 20641
rect 20810 20567 20866 20576
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 19922 20852 20334
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19446 20852 19858
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20732 19306 20852 19334
rect 20824 19242 20852 19306
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20810 19000 20866 19009
rect 20810 18935 20866 18944
rect 20628 18284 20680 18290
rect 20824 18272 20852 18935
rect 20916 18426 20944 19790
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20904 18284 20956 18290
rect 20824 18244 20904 18272
rect 20628 18226 20680 18232
rect 20904 18226 20956 18232
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 17116 20484 18158
rect 20534 17912 20590 17921
rect 20534 17847 20590 17856
rect 20548 17218 20576 17847
rect 20640 17338 20668 18226
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 17610 20760 18090
rect 21008 17678 21036 21014
rect 21100 20534 21128 21134
rect 21192 21010 21220 21830
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21100 20262 21128 20334
rect 21088 20256 21140 20262
rect 21086 20224 21088 20233
rect 21140 20224 21142 20233
rect 21086 20159 21142 20168
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21100 19378 21128 19994
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21100 17785 21128 19314
rect 21192 18426 21220 20810
rect 21284 20602 21312 21966
rect 21376 21690 21404 22102
rect 21468 22012 21496 22714
rect 21560 22409 21588 22714
rect 21652 22681 21680 23054
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21638 22672 21694 22681
rect 21638 22607 21694 22616
rect 21640 22432 21692 22438
rect 21546 22400 21602 22409
rect 21640 22374 21692 22380
rect 21546 22335 21602 22344
rect 21652 22234 21680 22374
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21744 22098 21772 22918
rect 21836 22574 21864 24822
rect 22376 24822 22428 24828
rect 21914 24783 21916 24792
rect 21968 24783 21970 24792
rect 21916 24754 21968 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22006 24440 22062 24449
rect 22062 24398 22140 24426
rect 22006 24375 22062 24384
rect 22112 24206 22140 24398
rect 22388 24206 22416 24550
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 21914 23896 21970 23905
rect 21914 23831 21970 23840
rect 22008 23860 22060 23866
rect 21928 23361 21956 23831
rect 22008 23802 22060 23808
rect 22020 23769 22048 23802
rect 22100 23792 22152 23798
rect 22006 23760 22062 23769
rect 22100 23734 22152 23740
rect 22006 23695 22062 23704
rect 21914 23352 21970 23361
rect 21914 23287 21916 23296
rect 21968 23287 21970 23296
rect 21916 23258 21968 23264
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21928 22710 21956 23054
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21824 22568 21876 22574
rect 21824 22510 21876 22516
rect 21822 22400 21878 22409
rect 21822 22335 21878 22344
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21548 22024 21600 22030
rect 21468 21984 21548 22012
rect 21548 21966 21600 21972
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21560 21554 21588 21966
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21652 21729 21680 21830
rect 21638 21720 21694 21729
rect 21836 21706 21864 22335
rect 21638 21655 21694 21664
rect 21744 21678 21864 21706
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21192 17882 21220 18362
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 20996 17672 21048 17678
rect 20902 17640 20958 17649
rect 20720 17604 20772 17610
rect 20772 17564 20852 17592
rect 20996 17614 21048 17620
rect 20902 17575 20958 17584
rect 20720 17546 20772 17552
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20548 17190 20760 17218
rect 20456 17088 20668 17116
rect 20456 16726 20484 17088
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20640 16590 20668 17088
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20732 16454 20760 17190
rect 20824 16658 20852 17564
rect 20916 17338 20944 17575
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 21100 17270 21128 17711
rect 21180 17672 21232 17678
rect 21284 17660 21312 19654
rect 21376 19009 21404 21490
rect 21454 21312 21510 21321
rect 21454 21247 21510 21256
rect 21468 19938 21496 21247
rect 21560 20942 21588 21490
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21652 20602 21680 21655
rect 21744 21146 21772 21678
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21914 21584 21970 21593
rect 21836 21146 21864 21558
rect 21914 21519 21916 21528
rect 21968 21519 21970 21528
rect 21916 21490 21968 21496
rect 22020 21434 22048 22918
rect 22112 22642 22140 23734
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22204 22953 22232 23666
rect 22284 23588 22336 23594
rect 22284 23530 22336 23536
rect 22296 23361 22324 23530
rect 22282 23352 22338 23361
rect 22282 23287 22338 23296
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22190 22944 22246 22953
rect 22190 22879 22246 22888
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22296 22574 22324 23122
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22204 22098 22232 22442
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21928 21406 22048 21434
rect 21928 21321 21956 21406
rect 22008 21344 22060 21350
rect 21914 21312 21970 21321
rect 22008 21286 22060 21292
rect 21914 21247 21970 21256
rect 22020 21146 22048 21286
rect 22204 21146 22232 21490
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 22008 21140 22060 21146
rect 22192 21140 22244 21146
rect 22008 21082 22060 21088
rect 22112 21100 22192 21128
rect 21822 21040 21878 21049
rect 21822 20975 21878 20984
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21652 20058 21680 20538
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21468 19910 21588 19938
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21468 19689 21496 19790
rect 21454 19680 21510 19689
rect 21454 19615 21510 19624
rect 21560 19446 21588 19910
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 19145 21496 19178
rect 21454 19136 21510 19145
rect 21454 19071 21510 19080
rect 21362 19000 21418 19009
rect 21652 18986 21680 19994
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21744 19378 21772 19926
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21362 18935 21418 18944
rect 21468 18958 21680 18986
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21376 18737 21404 18838
rect 21468 18766 21496 18958
rect 21732 18896 21784 18902
rect 21730 18864 21732 18873
rect 21784 18864 21786 18873
rect 21730 18799 21786 18808
rect 21456 18760 21508 18766
rect 21362 18728 21418 18737
rect 21456 18702 21508 18708
rect 21362 18663 21418 18672
rect 21836 18612 21864 20975
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22020 20074 22048 20470
rect 21928 20046 22048 20074
rect 21928 19854 21956 20046
rect 22112 19922 22140 21100
rect 22192 21082 22244 21088
rect 22296 20942 22324 22374
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22204 20262 22232 20878
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19990 22232 20198
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21916 19848 21968 19854
rect 22296 19836 22324 20742
rect 21916 19790 21968 19796
rect 22204 19808 22324 19836
rect 21928 19514 21956 19790
rect 22100 19712 22152 19718
rect 22006 19680 22062 19689
rect 22100 19654 22152 19660
rect 22006 19615 22062 19624
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21914 19408 21970 19417
rect 21914 19343 21970 19352
rect 21928 19174 21956 19343
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21928 18766 21956 19110
rect 22020 18902 22048 19615
rect 22112 19310 22140 19654
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 22204 18834 22232 19808
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 19009 22324 19246
rect 22282 19000 22338 19009
rect 22282 18935 22338 18944
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 21916 18760 21968 18766
rect 22100 18760 22152 18766
rect 21916 18702 21968 18708
rect 22098 18728 22100 18737
rect 22152 18728 22154 18737
rect 22098 18663 22154 18672
rect 21652 18584 21864 18612
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21376 17746 21404 18362
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21560 17882 21588 18226
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21232 17632 21312 17660
rect 21456 17672 21508 17678
rect 21362 17640 21418 17649
rect 21180 17614 21232 17620
rect 21456 17614 21508 17620
rect 21362 17575 21364 17584
rect 21416 17575 21418 17584
rect 21364 17546 21416 17552
rect 21468 17513 21496 17614
rect 21454 17504 21510 17513
rect 21454 17439 21510 17448
rect 21088 17264 21140 17270
rect 21364 17264 21416 17270
rect 21088 17206 21140 17212
rect 21362 17232 21364 17241
rect 21416 17232 21418 17241
rect 21362 17167 21418 17176
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 21100 16590 21128 16934
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21376 16522 21404 17167
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21468 16590 21496 17070
rect 21560 16658 21588 17818
rect 21652 17241 21680 18584
rect 22112 18442 22140 18663
rect 22192 18624 22244 18630
rect 22190 18592 22192 18601
rect 22244 18592 22246 18601
rect 22190 18527 22246 18536
rect 22112 18414 22232 18442
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21732 18148 21784 18154
rect 21732 18090 21784 18096
rect 21638 17232 21694 17241
rect 21744 17202 21772 18090
rect 21836 17921 21864 18226
rect 21822 17912 21878 17921
rect 21822 17847 21878 17856
rect 21836 17660 21864 17847
rect 21928 17814 21956 18226
rect 22008 18080 22060 18086
rect 22006 18048 22008 18057
rect 22060 18048 22062 18057
rect 22006 17983 22062 17992
rect 22020 17814 22048 17983
rect 22204 17921 22232 18414
rect 22388 18068 22416 24142
rect 22558 24032 22614 24041
rect 22558 23967 22614 23976
rect 22572 23730 22600 23967
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22468 23588 22520 23594
rect 22468 23530 22520 23536
rect 22480 21622 22508 23530
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22572 22030 22600 22578
rect 22664 22522 22692 26318
rect 22756 25140 22784 29106
rect 22848 25362 22876 33884
rect 22928 33866 22980 33872
rect 23032 33590 23060 34342
rect 23020 33584 23072 33590
rect 23020 33526 23072 33532
rect 23124 33436 23152 36615
rect 23216 35834 23244 36722
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23492 35630 23520 37046
rect 23584 35766 23612 37062
rect 23664 36576 23716 36582
rect 23664 36518 23716 36524
rect 23572 35760 23624 35766
rect 23572 35702 23624 35708
rect 23480 35624 23532 35630
rect 23480 35566 23532 35572
rect 23492 35193 23520 35566
rect 23478 35184 23534 35193
rect 23478 35119 23480 35128
rect 23532 35119 23534 35128
rect 23480 35090 23532 35096
rect 23296 34536 23348 34542
rect 23296 34478 23348 34484
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 23216 33522 23244 34138
rect 23308 33561 23336 34478
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23294 33552 23350 33561
rect 23204 33516 23256 33522
rect 23294 33487 23350 33496
rect 23204 33458 23256 33464
rect 23032 33408 23152 33436
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22940 30938 22968 31282
rect 22928 30932 22980 30938
rect 22928 30874 22980 30880
rect 22926 30696 22982 30705
rect 22926 30631 22982 30640
rect 22940 30394 22968 30631
rect 22928 30388 22980 30394
rect 22928 30330 22980 30336
rect 22926 30152 22982 30161
rect 22926 30087 22982 30096
rect 22940 29646 22968 30087
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 23032 29170 23060 33408
rect 23216 32910 23244 33458
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23112 30592 23164 30598
rect 23216 30580 23244 32846
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23164 30552 23244 30580
rect 23112 30534 23164 30540
rect 23110 30424 23166 30433
rect 23110 30359 23166 30368
rect 23124 29714 23152 30359
rect 23216 29889 23244 30552
rect 23308 30258 23336 31758
rect 23296 30252 23348 30258
rect 23296 30194 23348 30200
rect 23296 30116 23348 30122
rect 23296 30058 23348 30064
rect 23202 29880 23258 29889
rect 23202 29815 23258 29824
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 23110 29608 23166 29617
rect 23166 29566 23244 29594
rect 23110 29543 23166 29552
rect 23112 29504 23164 29510
rect 23112 29446 23164 29452
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 22928 29096 22980 29102
rect 22926 29064 22928 29073
rect 22980 29064 22982 29073
rect 22926 28999 22982 29008
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 22940 27130 22968 27338
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22928 25900 22980 25906
rect 22928 25842 22980 25848
rect 22940 25498 22968 25842
rect 22928 25492 22980 25498
rect 22928 25434 22980 25440
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22836 25152 22888 25158
rect 22756 25112 22836 25140
rect 22836 25094 22888 25100
rect 22742 24984 22798 24993
rect 22742 24919 22744 24928
rect 22796 24919 22798 24928
rect 22744 24890 22796 24896
rect 22848 24818 22876 25094
rect 23032 24834 23060 25366
rect 23124 24886 23152 29446
rect 23216 29170 23244 29566
rect 23308 29238 23336 30058
rect 23296 29232 23348 29238
rect 23296 29174 23348 29180
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23216 28762 23244 29106
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23400 27606 23428 33798
rect 23676 33522 23704 36518
rect 23768 35834 23796 37606
rect 23952 37274 23980 38830
rect 24504 38350 24532 38966
rect 24584 38956 24636 38962
rect 24584 38898 24636 38904
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 24596 38554 24624 38898
rect 24584 38548 24636 38554
rect 24584 38490 24636 38496
rect 24124 38344 24176 38350
rect 24124 38286 24176 38292
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24032 38208 24084 38214
rect 24032 38150 24084 38156
rect 24044 38010 24072 38150
rect 24032 38004 24084 38010
rect 24032 37946 24084 37952
rect 23860 37246 23980 37274
rect 24136 37262 24164 38286
rect 24216 37732 24268 37738
rect 24216 37674 24268 37680
rect 24228 37398 24256 37674
rect 24780 37670 24808 38898
rect 24872 38010 24900 39306
rect 25412 39296 25464 39302
rect 25412 39238 25464 39244
rect 25424 38962 25452 39238
rect 25976 38962 26004 39442
rect 26240 39296 26292 39302
rect 26240 39238 26292 39244
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25964 38956 26016 38962
rect 25964 38898 26016 38904
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 25332 37874 25360 38694
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 25412 38276 25464 38282
rect 25412 38218 25464 38224
rect 25424 38185 25452 38218
rect 25780 38208 25832 38214
rect 25410 38176 25466 38185
rect 25780 38150 25832 38156
rect 25410 38111 25466 38120
rect 24860 37868 24912 37874
rect 24860 37810 24912 37816
rect 25044 37868 25096 37874
rect 25044 37810 25096 37816
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24216 37392 24268 37398
rect 24216 37334 24268 37340
rect 24768 37324 24820 37330
rect 24768 37266 24820 37272
rect 23860 37194 23888 37246
rect 23952 37244 23980 37246
rect 24032 37256 24084 37262
rect 23952 37216 24032 37244
rect 24032 37198 24084 37204
rect 24124 37256 24176 37262
rect 24400 37256 24452 37262
rect 24124 37198 24176 37204
rect 24214 37224 24270 37233
rect 23848 37188 23900 37194
rect 24400 37198 24452 37204
rect 24214 37159 24216 37168
rect 23848 37130 23900 37136
rect 24268 37159 24270 37168
rect 24216 37130 24268 37136
rect 24412 36718 24440 37198
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24596 36922 24624 37062
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 24400 36712 24452 36718
rect 24400 36654 24452 36660
rect 24308 36576 24360 36582
rect 24308 36518 24360 36524
rect 24320 36242 24348 36518
rect 24308 36236 24360 36242
rect 24308 36178 24360 36184
rect 23756 35828 23808 35834
rect 23756 35770 23808 35776
rect 24320 35698 24348 36178
rect 24412 35698 24440 36654
rect 24780 36174 24808 37266
rect 24872 36854 24900 37810
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 24860 36848 24912 36854
rect 24860 36790 24912 36796
rect 24768 36168 24820 36174
rect 24964 36156 24992 37198
rect 25056 37126 25084 37810
rect 25228 37664 25280 37670
rect 25228 37606 25280 37612
rect 25240 37398 25268 37606
rect 25228 37392 25280 37398
rect 25228 37334 25280 37340
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 25044 36168 25096 36174
rect 24964 36128 25044 36156
rect 24768 36110 24820 36116
rect 25044 36110 25096 36116
rect 24492 35760 24544 35766
rect 24492 35702 24544 35708
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24412 35222 24440 35634
rect 24504 35290 24532 35702
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24688 35290 24716 35566
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24492 35284 24544 35290
rect 24492 35226 24544 35232
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 24400 35216 24452 35222
rect 24688 35170 24716 35226
rect 24400 35158 24452 35164
rect 24596 35142 24716 35170
rect 24872 35154 24900 35430
rect 24860 35148 24912 35154
rect 23756 34672 23808 34678
rect 23756 34614 23808 34620
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23492 31482 23520 31622
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23492 30802 23520 31418
rect 23584 31090 23612 33254
rect 23676 33017 23704 33458
rect 23662 33008 23718 33017
rect 23662 32943 23718 32952
rect 23676 32008 23704 32943
rect 23768 32434 23796 34614
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24400 34468 24452 34474
rect 24400 34410 24452 34416
rect 23848 34400 23900 34406
rect 23848 34342 23900 34348
rect 23860 33998 23888 34342
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 24032 33924 24084 33930
rect 24308 33924 24360 33930
rect 24032 33866 24084 33872
rect 24136 33884 24308 33912
rect 24044 33697 24072 33866
rect 24030 33688 24086 33697
rect 24030 33623 24086 33632
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23676 31980 23796 32008
rect 23664 31748 23716 31754
rect 23664 31690 23716 31696
rect 23676 31482 23704 31690
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 23768 31142 23796 31980
rect 23860 31890 23888 32302
rect 23952 32230 23980 32846
rect 24136 32434 24164 33884
rect 24308 33866 24360 33872
rect 24412 33658 24440 34410
rect 24504 33946 24532 34546
rect 24596 34202 24624 35142
rect 24860 35090 24912 35096
rect 24952 35148 25004 35154
rect 24952 35090 25004 35096
rect 24964 34762 24992 35090
rect 24688 34734 24992 34762
rect 24688 34678 24716 34734
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24584 34196 24636 34202
rect 24584 34138 24636 34144
rect 24674 33960 24730 33969
rect 24504 33918 24674 33946
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24216 33584 24268 33590
rect 24216 33526 24268 33532
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24124 32292 24176 32298
rect 24124 32234 24176 32240
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 32065 23980 32166
rect 23938 32056 23994 32065
rect 23938 31991 23994 32000
rect 23848 31884 23900 31890
rect 23848 31826 23900 31832
rect 23860 31346 23888 31826
rect 24030 31648 24086 31657
rect 24030 31583 24086 31592
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23756 31136 23808 31142
rect 23662 31104 23718 31113
rect 23584 31062 23662 31090
rect 23756 31078 23808 31084
rect 23662 31039 23718 31048
rect 23768 30920 23796 31078
rect 23676 30892 23796 30920
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23572 30796 23624 30802
rect 23572 30738 23624 30744
rect 23480 30388 23532 30394
rect 23480 30330 23532 30336
rect 23492 30190 23520 30330
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 23584 30138 23612 30738
rect 23676 30598 23704 30892
rect 23940 30864 23992 30870
rect 23940 30806 23992 30812
rect 23848 30728 23900 30734
rect 23846 30696 23848 30705
rect 23900 30696 23902 30705
rect 23846 30631 23902 30640
rect 23664 30592 23716 30598
rect 23664 30534 23716 30540
rect 23676 30258 23704 30534
rect 23952 30394 23980 30806
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 24044 30258 24072 31583
rect 24136 30870 24164 32234
rect 24124 30864 24176 30870
rect 24124 30806 24176 30812
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 23848 30184 23900 30190
rect 23584 30132 23848 30138
rect 23584 30126 23900 30132
rect 23584 30110 23888 30126
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 23492 29646 23520 29990
rect 23584 29714 23612 30110
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23676 29850 23704 29990
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23570 29608 23626 29617
rect 23570 29543 23572 29552
rect 23624 29543 23626 29552
rect 23664 29572 23716 29578
rect 23572 29514 23624 29520
rect 23664 29514 23716 29520
rect 23676 29306 23704 29514
rect 23768 29306 23796 29990
rect 23860 29458 23888 29990
rect 23860 29430 23980 29458
rect 23846 29336 23902 29345
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23756 29300 23808 29306
rect 23846 29271 23848 29280
rect 23756 29242 23808 29248
rect 23900 29271 23902 29280
rect 23848 29242 23900 29248
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 23676 28762 23704 29106
rect 23952 28994 23980 29430
rect 23860 28966 23980 28994
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23664 27872 23716 27878
rect 23664 27814 23716 27820
rect 23388 27600 23440 27606
rect 23294 27568 23350 27577
rect 23388 27542 23440 27548
rect 23478 27568 23534 27577
rect 23294 27503 23350 27512
rect 23308 27169 23336 27503
rect 23294 27160 23350 27169
rect 23294 27095 23350 27104
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23202 26480 23258 26489
rect 23202 26415 23258 26424
rect 23216 25906 23244 26415
rect 23308 26382 23336 26862
rect 23296 26376 23348 26382
rect 23400 26353 23428 27542
rect 23478 27503 23534 27512
rect 23572 27532 23624 27538
rect 23492 26994 23520 27503
rect 23572 27474 23624 27480
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23492 26586 23520 26930
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23296 26318 23348 26324
rect 23386 26344 23442 26353
rect 23386 26279 23442 26288
rect 23480 26308 23532 26314
rect 23400 26042 23428 26279
rect 23480 26250 23532 26256
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 25702 23428 25842
rect 23492 25838 23520 26250
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23204 25288 23256 25294
rect 23400 25265 23428 25638
rect 23204 25230 23256 25236
rect 23386 25256 23442 25265
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22940 24806 23060 24834
rect 23112 24880 23164 24886
rect 23112 24822 23164 24828
rect 22848 24614 22876 24754
rect 22836 24608 22888 24614
rect 22834 24576 22836 24585
rect 22888 24576 22890 24585
rect 22834 24511 22890 24520
rect 22834 24032 22890 24041
rect 22834 23967 22890 23976
rect 22744 22636 22796 22642
rect 22848 22624 22876 23967
rect 22940 23322 22968 24806
rect 23216 24750 23244 25230
rect 23386 25191 23442 25200
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23032 23798 23060 24550
rect 23216 24410 23244 24686
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 23308 24274 23336 25094
rect 23492 24274 23520 25774
rect 23584 25242 23612 27474
rect 23676 25906 23704 27814
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 23768 26897 23796 27406
rect 23754 26888 23810 26897
rect 23754 26823 23810 26832
rect 23768 26586 23796 26823
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23756 26376 23808 26382
rect 23860 26364 23888 28966
rect 24044 27470 24072 30194
rect 24124 30184 24176 30190
rect 24124 30126 24176 30132
rect 24136 30025 24164 30126
rect 24122 30016 24178 30025
rect 24122 29951 24178 29960
rect 24124 29504 24176 29510
rect 24124 29446 24176 29452
rect 24136 28762 24164 29446
rect 24228 29238 24256 33526
rect 24596 33522 24624 33918
rect 24674 33895 24730 33904
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24596 33134 24624 33458
rect 24504 33106 24624 33134
rect 24688 33114 24716 33798
rect 24676 33108 24728 33114
rect 24504 32994 24532 33106
rect 24676 33050 24728 33056
rect 24504 32966 24716 32994
rect 24492 32904 24544 32910
rect 24492 32846 24544 32852
rect 24504 32570 24532 32846
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24596 32434 24624 32710
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24308 32360 24360 32366
rect 24308 32302 24360 32308
rect 24320 31385 24348 32302
rect 24688 32298 24716 32966
rect 24780 32960 24808 34614
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24872 34202 24900 34478
rect 24865 34196 24917 34202
rect 24865 34138 24917 34144
rect 24964 33862 24992 34734
rect 25056 34542 25084 36110
rect 25424 36106 25452 38111
rect 25792 38010 25820 38150
rect 26160 38010 26188 38286
rect 25780 38004 25832 38010
rect 25780 37946 25832 37952
rect 26148 38004 26200 38010
rect 26148 37946 26200 37952
rect 25780 37800 25832 37806
rect 26252 37788 26280 39238
rect 26344 38350 26372 39578
rect 27068 39568 27120 39574
rect 26896 39516 27068 39522
rect 26896 39510 27120 39516
rect 26896 39494 27108 39510
rect 26896 39438 26924 39494
rect 27172 39438 27200 40326
rect 27252 40180 27304 40186
rect 27252 40122 27304 40128
rect 27264 39438 27292 40122
rect 27632 40118 27660 40326
rect 27620 40112 27672 40118
rect 27620 40054 27672 40060
rect 27436 40044 27488 40050
rect 27436 39986 27488 39992
rect 27448 39846 27476 39986
rect 27724 39930 27752 40938
rect 27540 39914 27752 39930
rect 27528 39908 27752 39914
rect 27580 39902 27752 39908
rect 27528 39850 27580 39856
rect 27436 39840 27488 39846
rect 27436 39782 27488 39788
rect 27620 39840 27672 39846
rect 27620 39782 27672 39788
rect 26884 39432 26936 39438
rect 26884 39374 26936 39380
rect 27068 39432 27120 39438
rect 27068 39374 27120 39380
rect 27160 39432 27212 39438
rect 27160 39374 27212 39380
rect 27252 39432 27304 39438
rect 27252 39374 27304 39380
rect 26896 39030 26924 39374
rect 26884 39024 26936 39030
rect 26884 38966 26936 38972
rect 27080 38962 27108 39374
rect 27252 39296 27304 39302
rect 27252 39238 27304 39244
rect 27344 39296 27396 39302
rect 27344 39238 27396 39244
rect 27264 39098 27292 39238
rect 27252 39092 27304 39098
rect 27252 39034 27304 39040
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 27252 38956 27304 38962
rect 27252 38898 27304 38904
rect 26332 38344 26384 38350
rect 26332 38286 26384 38292
rect 26516 38344 26568 38350
rect 26516 38286 26568 38292
rect 26332 37800 26384 37806
rect 25832 37760 25912 37788
rect 25780 37742 25832 37748
rect 25884 36582 25912 37760
rect 26252 37760 26332 37788
rect 26252 37670 26280 37760
rect 26332 37742 26384 37748
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 26252 36786 26280 37334
rect 26528 37126 26556 38286
rect 26700 37664 26752 37670
rect 26700 37606 26752 37612
rect 26712 37262 26740 37606
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 26516 37120 26568 37126
rect 26516 37062 26568 37068
rect 26608 37120 26660 37126
rect 26608 37062 26660 37068
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26424 36780 26476 36786
rect 26476 36740 26556 36768
rect 26424 36722 26476 36728
rect 26332 36644 26384 36650
rect 26332 36586 26384 36592
rect 25872 36576 25924 36582
rect 25872 36518 25924 36524
rect 25884 36378 25912 36518
rect 25872 36372 25924 36378
rect 25872 36314 25924 36320
rect 25596 36304 25648 36310
rect 25596 36246 25648 36252
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 25148 35562 25176 35634
rect 25332 35630 25360 36042
rect 25424 36009 25452 36042
rect 25504 36032 25556 36038
rect 25410 36000 25466 36009
rect 25504 35974 25556 35980
rect 25410 35935 25466 35944
rect 25412 35828 25464 35834
rect 25412 35770 25464 35776
rect 25320 35624 25372 35630
rect 25320 35566 25372 35572
rect 25136 35556 25188 35562
rect 25136 35498 25188 35504
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25240 35290 25268 35430
rect 25228 35284 25280 35290
rect 25228 35226 25280 35232
rect 25240 35086 25268 35226
rect 25228 35080 25280 35086
rect 25228 35022 25280 35028
rect 25424 34610 25452 35770
rect 25516 35086 25544 35974
rect 25608 35698 25636 36246
rect 25884 36122 25912 36314
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 25792 36094 25912 36122
rect 25792 35834 25820 36094
rect 25976 35873 26004 36178
rect 26344 36106 26372 36586
rect 26422 36408 26478 36417
rect 26422 36343 26478 36352
rect 26332 36100 26384 36106
rect 26332 36042 26384 36048
rect 26436 36038 26464 36343
rect 26056 36032 26108 36038
rect 26056 35974 26108 35980
rect 26424 36032 26476 36038
rect 26424 35974 26476 35980
rect 25962 35864 26018 35873
rect 25780 35828 25832 35834
rect 26068 35834 26096 35974
rect 25962 35799 26018 35808
rect 26056 35828 26108 35834
rect 25780 35770 25832 35776
rect 26056 35770 26108 35776
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 26148 35556 26200 35562
rect 26148 35498 26200 35504
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25872 35216 25924 35222
rect 25872 35158 25924 35164
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25780 35012 25832 35018
rect 25780 34954 25832 34960
rect 25688 34672 25740 34678
rect 25688 34614 25740 34620
rect 25412 34604 25464 34610
rect 25412 34546 25464 34552
rect 25044 34536 25096 34542
rect 25044 34478 25096 34484
rect 25056 34241 25084 34478
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25042 34232 25098 34241
rect 25042 34167 25098 34176
rect 25044 34128 25096 34134
rect 25148 34116 25176 34342
rect 25096 34088 25176 34116
rect 25044 34070 25096 34076
rect 24952 33856 25004 33862
rect 24858 33824 24914 33833
rect 24952 33798 25004 33804
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24858 33759 24914 33768
rect 24872 33590 24900 33759
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 24950 33416 25006 33425
rect 24872 33300 24900 33390
rect 25056 33402 25084 33798
rect 25424 33522 25452 34546
rect 25596 34400 25648 34406
rect 25596 34342 25648 34348
rect 25608 34241 25636 34342
rect 25594 34232 25650 34241
rect 25594 34167 25650 34176
rect 25700 34105 25728 34614
rect 25686 34096 25742 34105
rect 25686 34031 25742 34040
rect 25504 33992 25556 33998
rect 25504 33934 25556 33940
rect 25516 33697 25544 33934
rect 25688 33924 25740 33930
rect 25688 33866 25740 33872
rect 25502 33688 25558 33697
rect 25502 33623 25558 33632
rect 25228 33516 25280 33522
rect 25228 33458 25280 33464
rect 25412 33516 25464 33522
rect 25596 33516 25648 33522
rect 25464 33476 25544 33504
rect 25412 33458 25464 33464
rect 25006 33374 25084 33402
rect 24950 33351 25006 33360
rect 24872 33272 25176 33300
rect 24780 32932 24992 32960
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 24872 32570 24900 32778
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24872 32434 24900 32506
rect 24964 32434 24992 32932
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 25056 32570 25084 32710
rect 25044 32564 25096 32570
rect 25044 32506 25096 32512
rect 25148 32450 25176 33272
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 25056 32422 25176 32450
rect 24676 32292 24728 32298
rect 24728 32252 24808 32280
rect 24676 32234 24728 32240
rect 24674 32192 24730 32201
rect 24596 32150 24674 32178
rect 24400 31816 24452 31822
rect 24400 31758 24452 31764
rect 24412 31482 24440 31758
rect 24596 31482 24624 32150
rect 24674 32127 24730 32136
rect 24676 32020 24728 32026
rect 24676 31962 24728 31968
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24306 31376 24362 31385
rect 24306 31311 24362 31320
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 24412 30938 24440 31214
rect 24504 30938 24532 31418
rect 24582 31104 24638 31113
rect 24582 31039 24638 31048
rect 24596 30938 24624 31039
rect 24308 30932 24360 30938
rect 24308 30874 24360 30880
rect 24400 30932 24452 30938
rect 24400 30874 24452 30880
rect 24492 30932 24544 30938
rect 24492 30874 24544 30880
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24320 30841 24348 30874
rect 24306 30832 24362 30841
rect 24596 30802 24624 30874
rect 24688 30802 24716 31962
rect 24780 31822 24808 32252
rect 24964 31940 24992 32370
rect 24872 31912 24992 31940
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24780 31414 24808 31758
rect 24872 31414 24900 31912
rect 24950 31512 25006 31521
rect 25056 31498 25084 32422
rect 25136 32360 25188 32366
rect 25136 32302 25188 32308
rect 25148 31958 25176 32302
rect 25240 32230 25268 33458
rect 25516 32910 25544 33476
rect 25596 33458 25648 33464
rect 25504 32904 25556 32910
rect 25332 32864 25504 32892
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25226 32056 25282 32065
rect 25226 31991 25282 32000
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 25006 31470 25084 31498
rect 24950 31447 25006 31456
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24860 31408 24912 31414
rect 24860 31350 24912 31356
rect 24766 31104 24822 31113
rect 24766 31039 24822 31048
rect 24780 30802 24808 31039
rect 24306 30767 24362 30776
rect 24584 30796 24636 30802
rect 24320 30054 24348 30767
rect 24584 30738 24636 30744
rect 24676 30796 24728 30802
rect 24676 30738 24728 30744
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24412 29306 24440 30534
rect 24400 29300 24452 29306
rect 24400 29242 24452 29248
rect 24216 29232 24268 29238
rect 24216 29174 24268 29180
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24124 28756 24176 28762
rect 24124 28698 24176 28704
rect 24320 28506 24348 29106
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24412 28762 24440 28902
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24320 28478 24440 28506
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 24320 28218 24348 28358
rect 24412 28218 24440 28478
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24400 28212 24452 28218
rect 24400 28154 24452 28160
rect 24504 27606 24532 30602
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24584 30320 24636 30326
rect 24584 30262 24636 30268
rect 24674 30288 24730 30297
rect 24596 29646 24624 30262
rect 24780 30258 24808 30534
rect 24674 30223 24730 30232
rect 24768 30252 24820 30258
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24596 29170 24624 29582
rect 24688 29170 24716 30223
rect 24768 30194 24820 30200
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24688 29073 24716 29106
rect 24780 29102 24808 29582
rect 24872 29510 24900 31350
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24964 30977 24992 31282
rect 24950 30968 25006 30977
rect 25006 30926 25084 30954
rect 24950 30903 25006 30912
rect 24952 30796 25004 30802
rect 24952 30738 25004 30744
rect 24964 29782 24992 30738
rect 25056 30666 25084 30926
rect 25044 30660 25096 30666
rect 25044 30602 25096 30608
rect 25148 30394 25176 31894
rect 25240 31822 25268 31991
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25332 31414 25360 32864
rect 25504 32846 25556 32852
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25504 32428 25556 32434
rect 25504 32370 25556 32376
rect 25320 31408 25372 31414
rect 25240 31368 25320 31396
rect 25240 30580 25268 31368
rect 25320 31350 25372 31356
rect 25424 31226 25452 32370
rect 25516 31498 25544 32370
rect 25608 32230 25636 33458
rect 25700 33454 25728 33866
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25596 32224 25648 32230
rect 25594 32192 25596 32201
rect 25648 32192 25650 32201
rect 25594 32127 25650 32136
rect 25700 32042 25728 33254
rect 25792 32910 25820 34954
rect 25884 34610 25912 35158
rect 25976 35086 26004 35430
rect 25964 35080 26016 35086
rect 25964 35022 26016 35028
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 26068 34610 26096 34886
rect 25872 34604 25924 34610
rect 25872 34546 25924 34552
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 25884 33998 25912 34546
rect 25872 33992 25924 33998
rect 26068 33980 26096 34546
rect 26160 34542 26188 35498
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26148 34536 26200 34542
rect 26148 34478 26200 34484
rect 26252 34134 26280 35430
rect 26436 34678 26464 35974
rect 26528 35834 26556 36740
rect 26620 36378 26648 37062
rect 26804 36786 26832 37198
rect 26988 36854 27016 37198
rect 27080 37126 27108 38898
rect 27160 38208 27212 38214
rect 27264 38196 27292 38898
rect 27356 38350 27384 39238
rect 27448 38944 27476 39782
rect 27632 39574 27660 39782
rect 27620 39568 27672 39574
rect 27620 39510 27672 39516
rect 27816 39386 27844 41006
rect 27908 40594 27936 41958
rect 28724 41540 28776 41546
rect 28724 41482 28776 41488
rect 28356 41132 28408 41138
rect 28356 41074 28408 41080
rect 28368 40934 28396 41074
rect 28736 41070 28764 41482
rect 28816 41268 28868 41274
rect 28816 41210 28868 41216
rect 28828 41070 28856 41210
rect 28724 41064 28776 41070
rect 28724 41006 28776 41012
rect 28816 41064 28868 41070
rect 28816 41006 28868 41012
rect 29104 41018 29132 41958
rect 29184 41472 29236 41478
rect 29184 41414 29236 41420
rect 29196 41386 29408 41414
rect 29276 41064 29328 41070
rect 29104 40990 29224 41018
rect 29276 41006 29328 41012
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 27896 40588 27948 40594
rect 27896 40530 27948 40536
rect 29196 40526 29224 40990
rect 29184 40520 29236 40526
rect 29184 40462 29236 40468
rect 27896 40384 27948 40390
rect 27896 40326 27948 40332
rect 28816 40384 28868 40390
rect 28816 40326 28868 40332
rect 29000 40384 29052 40390
rect 29000 40326 29052 40332
rect 27908 39506 27936 40326
rect 27988 40112 28040 40118
rect 27988 40054 28040 40060
rect 27896 39500 27948 39506
rect 27896 39442 27948 39448
rect 27632 39358 27844 39386
rect 27528 38956 27580 38962
rect 27448 38916 27528 38944
rect 27528 38898 27580 38904
rect 27540 38350 27568 38898
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27528 38344 27580 38350
rect 27528 38286 27580 38292
rect 27264 38168 27476 38196
rect 27160 38150 27212 38156
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 26976 36848 27028 36854
rect 26976 36790 27028 36796
rect 26792 36780 26844 36786
rect 26792 36722 26844 36728
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26700 36236 26752 36242
rect 26700 36178 26752 36184
rect 26712 35834 26740 36178
rect 26988 36106 27016 36790
rect 27172 36786 27200 38150
rect 27448 37874 27476 38168
rect 27436 37868 27488 37874
rect 27436 37810 27488 37816
rect 27528 37868 27580 37874
rect 27632 37856 27660 39358
rect 28000 38282 28028 40054
rect 28724 39500 28776 39506
rect 28724 39442 28776 39448
rect 28264 39296 28316 39302
rect 28264 39238 28316 39244
rect 28078 38448 28134 38457
rect 28276 38418 28304 39238
rect 28736 38486 28764 39442
rect 28828 38894 28856 40326
rect 28908 39976 28960 39982
rect 28908 39918 28960 39924
rect 28920 39438 28948 39918
rect 28908 39432 28960 39438
rect 28908 39374 28960 39380
rect 28816 38888 28868 38894
rect 28816 38830 28868 38836
rect 28724 38480 28776 38486
rect 28724 38422 28776 38428
rect 28920 38418 28948 39374
rect 28078 38383 28134 38392
rect 28264 38412 28316 38418
rect 28092 38350 28120 38383
rect 28264 38354 28316 38360
rect 28908 38412 28960 38418
rect 28908 38354 28960 38360
rect 28080 38344 28132 38350
rect 28080 38286 28132 38292
rect 27988 38276 28040 38282
rect 27988 38218 28040 38224
rect 27580 37828 27660 37856
rect 27528 37810 27580 37816
rect 27448 37330 27476 37810
rect 27436 37324 27488 37330
rect 27436 37266 27488 37272
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 27540 36292 27568 37810
rect 27712 37664 27764 37670
rect 27712 37606 27764 37612
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 27632 36786 27660 37062
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27632 36394 27660 36722
rect 27724 36718 27752 37606
rect 27712 36712 27764 36718
rect 27712 36654 27764 36660
rect 28000 36417 28028 38218
rect 28814 38040 28870 38049
rect 28814 37975 28816 37984
rect 28868 37975 28870 37984
rect 28816 37946 28868 37952
rect 28448 37936 28500 37942
rect 28448 37878 28500 37884
rect 28354 36816 28410 36825
rect 28080 36780 28132 36786
rect 28354 36751 28356 36760
rect 28080 36722 28132 36728
rect 28408 36751 28410 36760
rect 28356 36722 28408 36728
rect 27986 36408 28042 36417
rect 27632 36366 27752 36394
rect 27540 36264 27660 36292
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 26700 35828 26752 35834
rect 26700 35770 26752 35776
rect 26712 35290 26740 35770
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 26700 35284 26752 35290
rect 26700 35226 26752 35232
rect 26700 34944 26752 34950
rect 26700 34886 26752 34892
rect 26712 34746 26740 34886
rect 26700 34740 26752 34746
rect 26700 34682 26752 34688
rect 26424 34672 26476 34678
rect 26424 34614 26476 34620
rect 26424 34468 26476 34474
rect 26424 34410 26476 34416
rect 26516 34468 26568 34474
rect 26516 34410 26568 34416
rect 26436 34202 26464 34410
rect 26528 34202 26556 34410
rect 26424 34196 26476 34202
rect 26424 34138 26476 34144
rect 26516 34196 26568 34202
rect 26516 34138 26568 34144
rect 26240 34128 26292 34134
rect 26240 34070 26292 34076
rect 26516 34060 26568 34066
rect 26568 34020 26648 34048
rect 26516 34002 26568 34008
rect 26148 33992 26200 33998
rect 26068 33952 26148 33980
rect 25872 33934 25924 33940
rect 26148 33934 26200 33940
rect 25964 33856 26016 33862
rect 25964 33798 26016 33804
rect 26056 33856 26108 33862
rect 26056 33798 26108 33804
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25608 32014 25728 32042
rect 25608 31686 25636 32014
rect 25792 31822 25820 32846
rect 25884 32434 25912 33390
rect 25976 33114 26004 33798
rect 25964 33108 26016 33114
rect 25964 33050 26016 33056
rect 26068 32586 26096 33798
rect 26160 33114 26188 33934
rect 26238 33552 26294 33561
rect 26238 33487 26240 33496
rect 26292 33487 26294 33496
rect 26240 33458 26292 33464
rect 26516 33448 26568 33454
rect 26516 33390 26568 33396
rect 26240 33380 26292 33386
rect 26240 33322 26292 33328
rect 26332 33380 26384 33386
rect 26332 33322 26384 33328
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 26252 32910 26280 33322
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 25976 32558 26096 32586
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25976 32178 26004 32558
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26240 32428 26292 32434
rect 26240 32370 26292 32376
rect 25884 32150 26004 32178
rect 25884 31822 25912 32150
rect 26068 32008 26096 32370
rect 26252 32026 26280 32370
rect 26344 32348 26372 33322
rect 26424 33108 26476 33114
rect 26424 33050 26476 33056
rect 26436 32910 26464 33050
rect 26424 32904 26476 32910
rect 26424 32846 26476 32852
rect 26424 32768 26476 32774
rect 26424 32710 26476 32716
rect 26436 32502 26464 32710
rect 26424 32496 26476 32502
rect 26528 32473 26556 33390
rect 26424 32438 26476 32444
rect 26514 32464 26570 32473
rect 26514 32399 26570 32408
rect 26344 32320 26464 32348
rect 26332 32224 26384 32230
rect 26330 32192 26332 32201
rect 26384 32192 26386 32201
rect 26330 32127 26386 32136
rect 25976 31980 26096 32008
rect 26240 32020 26292 32026
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25516 31470 25728 31498
rect 25884 31482 25912 31758
rect 25976 31482 26004 31980
rect 26240 31962 26292 31968
rect 26332 31952 26384 31958
rect 26332 31894 26384 31900
rect 26240 31884 26292 31890
rect 26240 31826 26292 31832
rect 26148 31816 26200 31822
rect 26068 31776 26148 31804
rect 26068 31521 26096 31776
rect 26148 31758 26200 31764
rect 26054 31512 26110 31521
rect 25608 31346 25636 31470
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25424 31198 25636 31226
rect 25320 31136 25372 31142
rect 25320 31078 25372 31084
rect 25332 30734 25360 31078
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25424 30580 25452 30670
rect 25504 30660 25556 30666
rect 25504 30602 25556 30608
rect 25240 30552 25452 30580
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25318 30288 25374 30297
rect 25424 30258 25452 30552
rect 25516 30258 25544 30602
rect 25608 30258 25636 31198
rect 25318 30223 25320 30232
rect 25372 30223 25374 30232
rect 25412 30252 25464 30258
rect 25320 30194 25372 30200
rect 25412 30194 25464 30200
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25410 30152 25466 30161
rect 25410 30087 25412 30096
rect 25464 30087 25466 30096
rect 25412 30058 25464 30064
rect 25516 30002 25544 30194
rect 25148 29974 25544 30002
rect 25608 30002 25636 30194
rect 25700 30190 25728 31470
rect 25872 31476 25924 31482
rect 25792 31436 25872 31464
rect 25792 30870 25820 31436
rect 25872 31418 25924 31424
rect 25964 31476 26016 31482
rect 26054 31447 26110 31456
rect 25964 31418 26016 31424
rect 26252 31414 26280 31826
rect 26240 31408 26292 31414
rect 25962 31376 26018 31385
rect 26240 31350 26292 31356
rect 26344 31346 26372 31894
rect 25962 31311 26018 31320
rect 26332 31340 26384 31346
rect 25976 31210 26004 31311
rect 26332 31282 26384 31288
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25872 31136 25924 31142
rect 26056 31136 26108 31142
rect 25872 31078 25924 31084
rect 25962 31104 26018 31113
rect 25884 30977 25912 31078
rect 26056 31078 26108 31084
rect 25962 31039 26018 31048
rect 25870 30968 25926 30977
rect 25870 30903 25926 30912
rect 25780 30864 25832 30870
rect 25780 30806 25832 30812
rect 25778 30560 25834 30569
rect 25884 30546 25912 30903
rect 25976 30648 26004 31039
rect 26068 30818 26096 31078
rect 26160 30938 26188 31214
rect 26436 31142 26464 32320
rect 26516 32292 26568 32298
rect 26516 32234 26568 32240
rect 26528 31346 26556 32234
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26424 31136 26476 31142
rect 26424 31078 26476 31084
rect 26330 30968 26386 30977
rect 26148 30932 26200 30938
rect 26330 30903 26386 30912
rect 26148 30874 26200 30880
rect 26344 30870 26372 30903
rect 26332 30864 26384 30870
rect 26068 30790 26188 30818
rect 26516 30864 26568 30870
rect 26384 30824 26464 30852
rect 26332 30806 26384 30812
rect 26056 30660 26108 30666
rect 25976 30620 26056 30648
rect 26056 30602 26108 30608
rect 25834 30518 25912 30546
rect 25778 30495 25834 30504
rect 25792 30258 25820 30495
rect 25870 30288 25926 30297
rect 25780 30252 25832 30258
rect 25870 30223 25926 30232
rect 25780 30194 25832 30200
rect 25688 30184 25740 30190
rect 25688 30126 25740 30132
rect 25778 30152 25834 30161
rect 25778 30087 25780 30096
rect 25832 30087 25834 30096
rect 25780 30058 25832 30064
rect 25608 29974 25820 30002
rect 25148 29850 25176 29974
rect 25226 29880 25282 29889
rect 25136 29844 25188 29850
rect 25792 29850 25820 29974
rect 25226 29815 25228 29824
rect 25136 29786 25188 29792
rect 25280 29815 25282 29824
rect 25780 29844 25832 29850
rect 25228 29786 25280 29792
rect 25780 29786 25832 29792
rect 24952 29776 25004 29782
rect 24952 29718 25004 29724
rect 25148 29578 25176 29786
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 24950 29472 25006 29481
rect 24950 29407 25006 29416
rect 24964 29322 24992 29407
rect 24964 29294 25176 29322
rect 25240 29306 25268 29582
rect 25688 29504 25740 29510
rect 25688 29446 25740 29452
rect 24964 29238 24992 29294
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 25042 29200 25098 29209
rect 25042 29135 25044 29144
rect 25096 29135 25098 29144
rect 25148 29152 25176 29294
rect 25228 29300 25280 29306
rect 25228 29242 25280 29248
rect 25504 29300 25556 29306
rect 25504 29242 25556 29248
rect 25412 29164 25464 29170
rect 25148 29124 25412 29152
rect 25044 29106 25096 29112
rect 25412 29106 25464 29112
rect 24768 29096 24820 29102
rect 24674 29064 24730 29073
rect 24768 29038 24820 29044
rect 24674 28999 24730 29008
rect 24674 28792 24730 28801
rect 24674 28727 24730 28736
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24400 27328 24452 27334
rect 24306 27296 24362 27305
rect 24400 27270 24452 27276
rect 24306 27231 24362 27240
rect 23808 26336 23888 26364
rect 23756 26318 23808 26324
rect 24320 26314 24348 27231
rect 24412 26926 24440 27270
rect 24504 26926 24532 27542
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24400 26920 24452 26926
rect 24400 26862 24452 26868
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24596 26586 24624 27406
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 23940 26308 23992 26314
rect 23940 26250 23992 26256
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23676 25673 23704 25842
rect 23662 25664 23718 25673
rect 23662 25599 23718 25608
rect 23952 25294 23980 26250
rect 24400 25968 24452 25974
rect 24688 25956 24716 28727
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 25056 28082 25084 28358
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 25318 27976 25374 27985
rect 25318 27911 25374 27920
rect 25332 27538 25360 27911
rect 25320 27532 25372 27538
rect 25372 27492 25452 27520
rect 25320 27474 25372 27480
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 24452 25928 24716 25956
rect 24400 25910 24452 25916
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24124 25832 24176 25838
rect 24228 25809 24256 25842
rect 24308 25832 24360 25838
rect 24124 25774 24176 25780
rect 24214 25800 24270 25809
rect 23940 25288 23992 25294
rect 23584 25214 23704 25242
rect 23940 25230 23992 25236
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24818 23612 25094
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23572 24608 23624 24614
rect 23570 24576 23572 24585
rect 23624 24576 23626 24585
rect 23570 24511 23626 24520
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23480 24268 23532 24274
rect 23532 24228 23612 24256
rect 23480 24210 23532 24216
rect 23388 24132 23440 24138
rect 23216 24092 23388 24120
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 23112 22976 23164 22982
rect 23112 22918 23164 22924
rect 23018 22808 23074 22817
rect 23018 22743 23074 22752
rect 22796 22596 22876 22624
rect 22928 22636 22980 22642
rect 22744 22578 22796 22584
rect 22928 22578 22980 22584
rect 22664 22494 22876 22522
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22560 21888 22612 21894
rect 22558 21856 22560 21865
rect 22612 21856 22614 21865
rect 22558 21791 22614 21800
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22480 20942 22508 21422
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22480 20534 22508 20878
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22466 20088 22522 20097
rect 22572 20074 22600 21791
rect 22664 21622 22692 22374
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 22756 21486 22784 21966
rect 22848 21706 22876 22494
rect 22940 21865 22968 22578
rect 22926 21856 22982 21865
rect 22926 21791 22982 21800
rect 22848 21678 22968 21706
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22744 21480 22796 21486
rect 22650 21448 22706 21457
rect 22744 21422 22796 21428
rect 22650 21383 22706 21392
rect 22522 20046 22600 20074
rect 22466 20023 22522 20032
rect 22468 19984 22520 19990
rect 22468 19926 22520 19932
rect 22480 18902 22508 19926
rect 22664 19666 22692 21383
rect 22848 21321 22876 21490
rect 22940 21434 22968 21678
rect 23032 21536 23060 22743
rect 23124 22030 23152 22918
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21865 23152 21966
rect 23110 21856 23166 21865
rect 23110 21791 23166 21800
rect 23112 21548 23164 21554
rect 23032 21508 23112 21536
rect 23112 21490 23164 21496
rect 22940 21406 23152 21434
rect 22928 21344 22980 21350
rect 22834 21312 22890 21321
rect 22928 21286 22980 21292
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22834 21247 22890 21256
rect 22742 21176 22798 21185
rect 22742 21111 22798 21120
rect 22756 21010 22784 21111
rect 22848 21078 22876 21247
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22756 20777 22784 20946
rect 22834 20904 22890 20913
rect 22834 20839 22890 20848
rect 22742 20768 22798 20777
rect 22742 20703 22798 20712
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22756 19786 22784 19994
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22572 19638 22692 19666
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22480 18222 22508 18566
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22388 18040 22508 18068
rect 22190 17912 22246 17921
rect 22190 17847 22246 17856
rect 21916 17808 21968 17814
rect 22008 17808 22060 17814
rect 21968 17768 22008 17796
rect 21916 17750 21968 17756
rect 22008 17750 22060 17756
rect 21916 17672 21968 17678
rect 21836 17632 21916 17660
rect 21916 17614 21968 17620
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22388 17252 22416 17614
rect 22480 17338 22508 18040
rect 22572 17882 22600 19638
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22664 19334 22692 19450
rect 22664 19306 22784 19334
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22664 18358 22692 19178
rect 22756 18834 22784 19306
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22848 18578 22876 20839
rect 22940 20466 22968 21286
rect 23032 20505 23060 21286
rect 23124 20942 23152 21406
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23018 20496 23074 20505
rect 22928 20460 22980 20466
rect 23018 20431 23074 20440
rect 22928 20402 22980 20408
rect 23124 20380 23152 20878
rect 23032 20352 23152 20380
rect 22926 19680 22982 19689
rect 22926 19615 22982 19624
rect 22940 18970 22968 19615
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 22756 18550 22876 18578
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22296 17224 22416 17252
rect 21638 17167 21694 17176
rect 21732 17196 21784 17202
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 20272 15706 20300 15982
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 13372 9654 13400 14214
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 11624 6798 11652 9590
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 18524 5574 18552 15574
rect 21376 15570 21404 16118
rect 21652 15978 21680 17167
rect 21732 17138 21784 17144
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16454 21956 16934
rect 22020 16574 22048 17002
rect 22100 16584 22152 16590
rect 22020 16546 22100 16574
rect 22100 16526 22152 16532
rect 22296 16454 22324 17224
rect 22480 16674 22508 17274
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22388 16658 22508 16674
rect 22376 16652 22508 16658
rect 22428 16646 22508 16652
rect 22376 16594 22428 16600
rect 22468 16584 22520 16590
rect 22560 16584 22612 16590
rect 22468 16526 22520 16532
rect 22558 16552 22560 16561
rect 22612 16552 22614 16561
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22480 16250 22508 16526
rect 22664 16522 22692 17206
rect 22558 16487 22614 16496
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 22480 15706 22508 16186
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 22756 15434 22784 18550
rect 23032 18222 23060 20352
rect 23110 19816 23166 19825
rect 23110 19751 23166 19760
rect 23124 19514 23152 19751
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 22928 18216 22980 18222
rect 22834 18184 22890 18193
rect 22928 18158 22980 18164
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22834 18119 22890 18128
rect 22848 17338 22876 18119
rect 22940 17610 22968 18158
rect 23124 17678 23152 18566
rect 23216 17882 23244 24092
rect 23388 24074 23440 24080
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23308 23322 23336 23734
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 22574 23336 22918
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23400 22137 23428 23734
rect 23492 23730 23520 24006
rect 23584 23730 23612 24228
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23492 23118 23520 23666
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23492 22778 23520 23054
rect 23572 22976 23624 22982
rect 23676 22964 23704 25214
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23768 24342 23796 24754
rect 24044 24410 24072 25230
rect 24136 24886 24164 25774
rect 24308 25774 24360 25780
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24964 25786 24992 26930
rect 25056 26586 25084 26930
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25240 25838 25268 26998
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25332 26382 25360 26862
rect 25424 26450 25452 27492
rect 25516 26450 25544 29242
rect 25700 29170 25728 29446
rect 25688 29164 25740 29170
rect 25688 29106 25740 29112
rect 25700 28490 25728 29106
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25884 28082 25912 30223
rect 26068 30054 26096 30602
rect 25964 30048 26016 30054
rect 25964 29990 26016 29996
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 25608 27334 25636 27406
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25504 26444 25556 26450
rect 25504 26386 25556 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25228 25832 25280 25838
rect 25226 25800 25228 25809
rect 25280 25800 25282 25809
rect 24214 25735 24270 25744
rect 24320 25129 24348 25774
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24492 25424 24544 25430
rect 24492 25366 24544 25372
rect 24400 25220 24452 25226
rect 24400 25162 24452 25168
rect 24306 25120 24362 25129
rect 24306 25055 24362 25064
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 23756 24336 23808 24342
rect 24136 24290 24164 24822
rect 24320 24698 24348 25055
rect 24412 24818 24440 25162
rect 24504 24954 24532 25366
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24596 24993 24624 25230
rect 24582 24984 24638 24993
rect 24492 24948 24544 24954
rect 24582 24919 24584 24928
rect 24492 24890 24544 24896
rect 24636 24919 24638 24928
rect 24584 24890 24636 24896
rect 24400 24812 24452 24818
rect 24504 24800 24532 24890
rect 24688 24886 24716 25434
rect 24872 25362 24900 25774
rect 24964 25758 25176 25786
rect 25148 25498 25176 25758
rect 25226 25735 25282 25744
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25424 25430 25452 26386
rect 25608 25906 25636 27270
rect 25700 26994 25728 27814
rect 25884 27713 25912 28018
rect 25870 27704 25926 27713
rect 25870 27639 25926 27648
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25596 25900 25648 25906
rect 25596 25842 25648 25848
rect 25412 25424 25464 25430
rect 25412 25366 25464 25372
rect 24860 25356 24912 25362
rect 24780 25316 24860 25344
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24584 24812 24636 24818
rect 24504 24772 24584 24800
rect 24400 24754 24452 24760
rect 24584 24754 24636 24760
rect 24412 24721 24440 24754
rect 23756 24278 23808 24284
rect 23952 24262 24164 24290
rect 24228 24670 24348 24698
rect 24398 24712 24454 24721
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23768 23526 23796 23802
rect 23952 23730 23980 24262
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23952 23322 23980 23666
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 23676 22936 23980 22964
rect 23572 22918 23624 22924
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23584 22624 23612 22918
rect 23756 22636 23808 22642
rect 23584 22596 23704 22624
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23386 22128 23442 22137
rect 23386 22063 23442 22072
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23308 21321 23336 21830
rect 23294 21312 23350 21321
rect 23294 21247 23350 21256
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23308 20466 23336 21082
rect 23400 20942 23428 21898
rect 23492 21146 23520 22510
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23584 21622 23612 22442
rect 23676 22030 23704 22596
rect 23756 22578 23808 22584
rect 23768 22098 23796 22578
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23308 20097 23336 20198
rect 23294 20088 23350 20097
rect 23294 20023 23350 20032
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19378 23336 19858
rect 23492 19802 23520 20402
rect 23584 19825 23612 21422
rect 23676 21049 23704 21830
rect 23860 21622 23888 21966
rect 23848 21616 23900 21622
rect 23952 21593 23980 22936
rect 24044 22001 24072 24142
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 23730 24164 24006
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24124 23044 24176 23050
rect 24124 22986 24176 22992
rect 24030 21992 24086 22001
rect 24030 21927 24032 21936
rect 24084 21927 24086 21936
rect 24032 21898 24084 21904
rect 23848 21558 23900 21564
rect 23938 21584 23994 21593
rect 24136 21554 24164 22986
rect 24228 22234 24256 24670
rect 24596 24682 24624 24754
rect 24398 24647 24454 24656
rect 24492 24676 24544 24682
rect 24492 24618 24544 24624
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24504 24562 24532 24618
rect 24320 24138 24348 24550
rect 24504 24534 24716 24562
rect 24308 24132 24360 24138
rect 24308 24074 24360 24080
rect 24584 24132 24636 24138
rect 24584 24074 24636 24080
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24306 23488 24362 23497
rect 24306 23423 24362 23432
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24124 21548 24176 21554
rect 23994 21528 24072 21536
rect 23938 21519 24072 21528
rect 23952 21508 24072 21519
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23848 21480 23900 21486
rect 23900 21440 23980 21468
rect 23848 21422 23900 21428
rect 23662 21040 23718 21049
rect 23662 20975 23718 20984
rect 23662 20904 23718 20913
rect 23662 20839 23718 20848
rect 23676 20806 23704 20839
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20262 23704 20742
rect 23768 20262 23796 21422
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23860 20874 23888 21286
rect 23952 20942 23980 21440
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24044 20874 24072 21508
rect 24176 21508 24256 21536
rect 24124 21490 24176 21496
rect 24228 20890 24256 21508
rect 24320 21128 24348 23423
rect 24412 22778 24440 24006
rect 24596 23225 24624 24074
rect 24582 23216 24638 23225
rect 24582 23151 24638 23160
rect 24596 22778 24624 23151
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24398 22672 24454 22681
rect 24398 22607 24400 22616
rect 24452 22607 24454 22616
rect 24492 22636 24544 22642
rect 24400 22578 24452 22584
rect 24492 22578 24544 22584
rect 24412 22234 24440 22578
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24504 21894 24532 22578
rect 24688 22166 24716 24534
rect 24780 24410 24808 25316
rect 24860 25298 24912 25304
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 25332 24886 25360 25162
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25320 24880 25372 24886
rect 25320 24822 25372 24828
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24780 24206 24808 24346
rect 24872 24206 24900 24618
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24872 23848 24900 24142
rect 24780 23820 24900 23848
rect 24780 23730 24808 23820
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24872 23225 24900 23666
rect 24858 23216 24914 23225
rect 24858 23151 24914 23160
rect 24964 23050 24992 24550
rect 25056 24410 25084 24822
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25044 23792 25096 23798
rect 25148 23780 25176 24686
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25096 23752 25176 23780
rect 25044 23734 25096 23740
rect 25044 23588 25096 23594
rect 25044 23530 25096 23536
rect 25056 23186 25084 23530
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25148 23322 25176 23462
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24780 22642 24808 22986
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24872 22522 24900 22986
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25148 22710 25176 22918
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 24872 22494 25084 22522
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24584 22160 24636 22166
rect 24584 22102 24636 22108
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24766 22128 24822 22137
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21486 24532 21830
rect 24596 21622 24624 22102
rect 24766 22063 24822 22072
rect 24780 22030 24808 22063
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24688 21865 24716 21898
rect 24768 21888 24820 21894
rect 24674 21856 24730 21865
rect 24768 21830 24820 21836
rect 24674 21791 24730 21800
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24492 21480 24544 21486
rect 24544 21440 24624 21468
rect 24492 21422 24544 21428
rect 24400 21140 24452 21146
rect 24320 21100 24400 21128
rect 24400 21082 24452 21088
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 24032 20868 24084 20874
rect 24228 20862 24348 20890
rect 24032 20810 24084 20816
rect 23940 20800 23992 20806
rect 23846 20768 23902 20777
rect 24216 20800 24268 20806
rect 24030 20768 24086 20777
rect 23992 20748 24030 20754
rect 23940 20742 24030 20748
rect 23952 20726 24030 20742
rect 23846 20703 23902 20712
rect 24216 20742 24268 20748
rect 24030 20703 24086 20712
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23860 20074 23888 20703
rect 23938 20632 23994 20641
rect 23938 20567 23994 20576
rect 23676 20046 23888 20074
rect 23400 19774 23520 19802
rect 23570 19816 23626 19825
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23294 19272 23350 19281
rect 23294 19207 23350 19216
rect 23308 18601 23336 19207
rect 23400 18970 23428 19774
rect 23570 19751 23626 19760
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23492 19242 23520 19654
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23480 18896 23532 18902
rect 23584 18884 23612 19382
rect 23532 18856 23612 18884
rect 23480 18838 23532 18844
rect 23676 18766 23704 20046
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19378 23796 19654
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23860 18986 23888 19858
rect 23952 19378 23980 20567
rect 24030 20496 24086 20505
rect 24086 20466 24164 20482
rect 24228 20466 24256 20742
rect 24086 20460 24176 20466
rect 24086 20454 24124 20460
rect 24030 20431 24086 20440
rect 24124 20402 24176 20408
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24214 20360 24270 20369
rect 24044 19990 24072 20334
rect 24214 20295 24270 20304
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 24136 19446 24164 19994
rect 24228 19990 24256 20295
rect 24320 20262 24348 20862
rect 24412 20398 24440 21082
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24504 20602 24532 20742
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24596 20534 24624 21440
rect 24688 20874 24716 21791
rect 24780 21690 24808 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24780 20924 24808 21626
rect 24872 21486 24900 22374
rect 24964 21486 24992 22374
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 24860 20936 24912 20942
rect 24780 20896 24860 20924
rect 24860 20878 24912 20884
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24584 20528 24636 20534
rect 24964 20482 24992 21422
rect 25056 21049 25084 22494
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25240 21978 25268 24006
rect 25332 23866 25360 24550
rect 25424 24410 25452 25366
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25516 24274 25544 24754
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25516 23866 25544 24210
rect 25608 24206 25636 24822
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 22692 25360 23462
rect 25412 23248 25464 23254
rect 25412 23190 25464 23196
rect 25424 23089 25452 23190
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25332 22664 25452 22692
rect 25148 21876 25176 21966
rect 25240 21950 25360 21978
rect 25148 21848 25268 21876
rect 25042 21040 25098 21049
rect 25042 20975 25098 20984
rect 25240 20942 25268 21848
rect 25332 21593 25360 21950
rect 25318 21584 25374 21593
rect 25318 21519 25374 21528
rect 25320 21140 25372 21146
rect 25424 21128 25452 22664
rect 25608 22658 25636 24142
rect 25700 24070 25728 26726
rect 25884 26586 25912 26930
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25780 26376 25832 26382
rect 25884 26353 25912 26522
rect 25976 26450 26004 29990
rect 26068 29510 26096 29990
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 26160 28994 26188 30790
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 26252 29102 26280 30058
rect 26332 29572 26384 29578
rect 26332 29514 26384 29520
rect 26436 29560 26464 30824
rect 26516 30806 26568 30812
rect 26528 30716 26556 30806
rect 26620 30784 26648 34020
rect 26700 33992 26752 33998
rect 26698 33960 26700 33969
rect 26752 33960 26754 33969
rect 26698 33895 26754 33904
rect 26712 33697 26740 33895
rect 26698 33688 26754 33697
rect 26698 33623 26754 33632
rect 26804 33590 26832 35566
rect 26884 35080 26936 35086
rect 26884 35022 26936 35028
rect 26896 34921 26924 35022
rect 26882 34912 26938 34921
rect 26882 34847 26938 34856
rect 26988 34610 27016 36042
rect 27344 35692 27396 35698
rect 27540 35680 27568 36264
rect 27396 35652 27568 35680
rect 27344 35634 27396 35640
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 26976 34604 27028 34610
rect 26976 34546 27028 34552
rect 26884 34536 26936 34542
rect 26884 34478 26936 34484
rect 26792 33584 26844 33590
rect 26792 33526 26844 33532
rect 26896 33318 26924 34478
rect 27172 34406 27200 35566
rect 27632 35290 27660 36264
rect 27620 35284 27672 35290
rect 27620 35226 27672 35232
rect 27724 34746 27752 36366
rect 28092 36378 28120 36722
rect 27986 36343 28042 36352
rect 28080 36372 28132 36378
rect 28000 36145 28028 36343
rect 28080 36314 28132 36320
rect 28172 36372 28224 36378
rect 28172 36314 28224 36320
rect 27986 36136 28042 36145
rect 27986 36071 28042 36080
rect 27896 36032 27948 36038
rect 27896 35974 27948 35980
rect 27988 36032 28040 36038
rect 27988 35974 28040 35980
rect 27908 35601 27936 35974
rect 27894 35592 27950 35601
rect 27894 35527 27950 35536
rect 27896 35216 27948 35222
rect 27896 35158 27948 35164
rect 27712 34740 27764 34746
rect 27712 34682 27764 34688
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 27160 34400 27212 34406
rect 27160 34342 27212 34348
rect 27344 34400 27396 34406
rect 27344 34342 27396 34348
rect 27158 34232 27214 34241
rect 27068 34196 27120 34202
rect 27158 34167 27214 34176
rect 27068 34138 27120 34144
rect 27080 33998 27108 34138
rect 27172 33998 27200 34167
rect 27068 33992 27120 33998
rect 27068 33934 27120 33940
rect 27160 33992 27212 33998
rect 27212 33952 27292 33980
rect 27160 33934 27212 33940
rect 26884 33312 26936 33318
rect 26884 33254 26936 33260
rect 26792 33108 26844 33114
rect 26792 33050 26844 33056
rect 26700 32768 26752 32774
rect 26700 32710 26752 32716
rect 26712 31346 26740 32710
rect 26804 32026 26832 33050
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 26884 32768 26936 32774
rect 26884 32710 26936 32716
rect 26896 32570 26924 32710
rect 26884 32564 26936 32570
rect 26884 32506 26936 32512
rect 26884 32428 26936 32434
rect 26884 32370 26936 32376
rect 26896 32201 26924 32370
rect 26988 32366 27016 32846
rect 26976 32360 27028 32366
rect 26976 32302 27028 32308
rect 26976 32224 27028 32230
rect 26882 32192 26938 32201
rect 26976 32166 27028 32172
rect 26882 32127 26938 32136
rect 26988 32065 27016 32166
rect 26974 32056 27030 32065
rect 26792 32020 26844 32026
rect 26974 31991 27030 32000
rect 26792 31962 26844 31968
rect 27080 31906 27108 33934
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 26884 31884 26936 31890
rect 26988 31878 27108 31906
rect 26988 31872 27016 31878
rect 26936 31844 27016 31872
rect 26884 31826 26936 31832
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 27068 31816 27120 31822
rect 27172 31804 27200 33798
rect 27264 33590 27292 33952
rect 27252 33584 27304 33590
rect 27252 33526 27304 33532
rect 27356 33386 27384 34342
rect 27540 34082 27568 34546
rect 27802 34368 27858 34377
rect 27724 34326 27802 34354
rect 27724 34134 27752 34326
rect 27802 34303 27858 34312
rect 27620 34128 27672 34134
rect 27448 34054 27568 34082
rect 27618 34096 27620 34105
rect 27712 34128 27764 34134
rect 27672 34096 27674 34105
rect 27448 33930 27476 34054
rect 27712 34070 27764 34076
rect 27618 34031 27674 34040
rect 27908 33998 27936 35158
rect 28000 34388 28028 35974
rect 28184 35630 28212 36314
rect 28354 36272 28410 36281
rect 28460 36242 28488 37878
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28724 37392 28776 37398
rect 28644 37340 28724 37346
rect 28644 37334 28776 37340
rect 28644 37318 28764 37334
rect 28644 36786 28672 37318
rect 28920 37233 28948 37742
rect 28906 37224 28962 37233
rect 28906 37159 28962 37168
rect 28722 36952 28778 36961
rect 28722 36887 28778 36896
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28540 36712 28592 36718
rect 28540 36654 28592 36660
rect 28552 36242 28580 36654
rect 28644 36553 28672 36722
rect 28630 36544 28686 36553
rect 28630 36479 28686 36488
rect 28736 36378 28764 36887
rect 29012 36786 29040 40326
rect 29184 40044 29236 40050
rect 29104 40004 29184 40032
rect 29104 39846 29132 40004
rect 29184 39986 29236 39992
rect 29092 39840 29144 39846
rect 29092 39782 29144 39788
rect 29184 39296 29236 39302
rect 29184 39238 29236 39244
rect 29092 38752 29144 38758
rect 29092 38694 29144 38700
rect 29104 37874 29132 38694
rect 29196 38350 29224 39238
rect 29288 39098 29316 41006
rect 29380 40730 29408 41386
rect 29644 41268 29696 41274
rect 29644 41210 29696 41216
rect 29460 40928 29512 40934
rect 29460 40870 29512 40876
rect 29552 40928 29604 40934
rect 29552 40870 29604 40876
rect 29368 40724 29420 40730
rect 29368 40666 29420 40672
rect 29368 40384 29420 40390
rect 29368 40326 29420 40332
rect 29380 39370 29408 40326
rect 29368 39364 29420 39370
rect 29368 39306 29420 39312
rect 29276 39092 29328 39098
rect 29276 39034 29328 39040
rect 29368 39092 29420 39098
rect 29368 39034 29420 39040
rect 29380 38962 29408 39034
rect 29368 38956 29420 38962
rect 29368 38898 29420 38904
rect 29276 38548 29328 38554
rect 29276 38490 29328 38496
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29092 37868 29144 37874
rect 29092 37810 29144 37816
rect 29288 37330 29316 38490
rect 29368 38412 29420 38418
rect 29368 38354 29420 38360
rect 29380 37618 29408 38354
rect 29472 37874 29500 40870
rect 29564 39098 29592 40870
rect 29656 40186 29684 41210
rect 29748 40730 29960 40746
rect 29736 40724 29960 40730
rect 29788 40718 29960 40724
rect 29736 40666 29788 40672
rect 29828 40588 29880 40594
rect 29828 40530 29880 40536
rect 29736 40384 29788 40390
rect 29736 40326 29788 40332
rect 29644 40180 29696 40186
rect 29644 40122 29696 40128
rect 29656 39098 29684 40122
rect 29552 39092 29604 39098
rect 29552 39034 29604 39040
rect 29644 39092 29696 39098
rect 29644 39034 29696 39040
rect 29644 38956 29696 38962
rect 29644 38898 29696 38904
rect 29656 38010 29684 38898
rect 29644 38004 29696 38010
rect 29644 37946 29696 37952
rect 29460 37868 29512 37874
rect 29460 37810 29512 37816
rect 29552 37664 29604 37670
rect 29380 37590 29500 37618
rect 29552 37606 29604 37612
rect 29276 37324 29328 37330
rect 29276 37266 29328 37272
rect 29276 37120 29328 37126
rect 29276 37062 29328 37068
rect 29184 36848 29236 36854
rect 29184 36790 29236 36796
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28814 36408 28870 36417
rect 28724 36372 28776 36378
rect 28814 36343 28870 36352
rect 28724 36314 28776 36320
rect 28828 36310 28856 36343
rect 28816 36304 28868 36310
rect 28816 36246 28868 36252
rect 28920 36242 28948 36586
rect 29000 36576 29052 36582
rect 29092 36576 29144 36582
rect 29000 36518 29052 36524
rect 29090 36544 29092 36553
rect 29144 36544 29146 36553
rect 28354 36207 28410 36216
rect 28448 36236 28500 36242
rect 28368 36038 28396 36207
rect 28448 36178 28500 36184
rect 28540 36236 28592 36242
rect 28540 36178 28592 36184
rect 28632 36236 28684 36242
rect 28632 36178 28684 36184
rect 28908 36236 28960 36242
rect 28908 36178 28960 36184
rect 28552 36038 28580 36178
rect 28356 36032 28408 36038
rect 28356 35974 28408 35980
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28552 35873 28580 35974
rect 28538 35864 28594 35873
rect 28538 35799 28594 35808
rect 28264 35692 28316 35698
rect 28264 35634 28316 35640
rect 28172 35624 28224 35630
rect 28172 35566 28224 35572
rect 28172 35488 28224 35494
rect 28172 35430 28224 35436
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 28092 34542 28120 35022
rect 28184 34746 28212 35430
rect 28276 35222 28304 35634
rect 28644 35290 28672 36178
rect 28724 36032 28776 36038
rect 28724 35974 28776 35980
rect 28632 35284 28684 35290
rect 28632 35226 28684 35232
rect 28264 35216 28316 35222
rect 28264 35158 28316 35164
rect 28356 35148 28408 35154
rect 28356 35090 28408 35096
rect 28368 34746 28396 35090
rect 28448 34944 28500 34950
rect 28448 34886 28500 34892
rect 28540 34944 28592 34950
rect 28540 34886 28592 34892
rect 28460 34746 28488 34886
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 28356 34740 28408 34746
rect 28356 34682 28408 34688
rect 28448 34740 28500 34746
rect 28448 34682 28500 34688
rect 28080 34536 28132 34542
rect 28080 34478 28132 34484
rect 28552 34406 28580 34886
rect 28540 34400 28592 34406
rect 28000 34360 28120 34388
rect 27986 34096 28042 34105
rect 27986 34031 27988 34040
rect 28040 34031 28042 34040
rect 27988 34002 28040 34008
rect 28092 33998 28120 34360
rect 28262 34368 28318 34377
rect 28540 34342 28592 34348
rect 28262 34303 28318 34312
rect 28276 33998 28304 34303
rect 28356 34060 28408 34066
rect 28356 34002 28408 34008
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27896 33992 27948 33998
rect 27896 33934 27948 33940
rect 28080 33992 28132 33998
rect 28264 33992 28316 33998
rect 28132 33952 28212 33980
rect 28080 33934 28132 33940
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27344 33380 27396 33386
rect 27344 33322 27396 33328
rect 27344 32972 27396 32978
rect 27344 32914 27396 32920
rect 27252 32768 27304 32774
rect 27252 32710 27304 32716
rect 27264 32434 27292 32710
rect 27356 32570 27384 32914
rect 27540 32910 27568 33934
rect 27620 33856 27672 33862
rect 27618 33824 27620 33833
rect 27712 33856 27764 33862
rect 27672 33824 27674 33833
rect 28080 33856 28132 33862
rect 27764 33816 28028 33844
rect 27712 33798 27764 33804
rect 27618 33759 27674 33768
rect 27632 32978 27660 33759
rect 27724 33658 27752 33798
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 27712 33312 27764 33318
rect 27712 33254 27764 33260
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 27528 32904 27580 32910
rect 27448 32864 27528 32892
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27252 32428 27304 32434
rect 27252 32370 27304 32376
rect 27344 32360 27396 32366
rect 27344 32302 27396 32308
rect 27356 31890 27384 32302
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 27120 31776 27200 31804
rect 27068 31758 27120 31764
rect 26804 31362 26832 31758
rect 26976 31680 27028 31686
rect 26976 31622 27028 31628
rect 27068 31680 27120 31686
rect 27068 31622 27120 31628
rect 26700 31340 26752 31346
rect 26804 31334 26924 31362
rect 26700 31282 26752 31288
rect 26620 30756 26832 30784
rect 26528 30688 26648 30716
rect 26514 30288 26570 30297
rect 26514 30223 26516 30232
rect 26568 30223 26570 30232
rect 26516 30194 26568 30200
rect 26516 29572 26568 29578
rect 26436 29532 26516 29560
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26068 28966 26188 28994
rect 26068 27470 26096 28966
rect 26252 28626 26280 29038
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 26344 28490 26372 29514
rect 26436 29170 26464 29532
rect 26516 29514 26568 29520
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26422 28792 26478 28801
rect 26422 28727 26424 28736
rect 26476 28727 26478 28736
rect 26424 28698 26476 28704
rect 26620 28694 26648 30688
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26712 30054 26740 30534
rect 26804 30258 26832 30756
rect 26792 30252 26844 30258
rect 26792 30194 26844 30200
rect 26700 30048 26752 30054
rect 26700 29990 26752 29996
rect 26804 29850 26832 30194
rect 26896 30122 26924 31334
rect 26988 30870 27016 31622
rect 27080 31521 27108 31622
rect 27066 31512 27122 31521
rect 27066 31447 27122 31456
rect 26976 30864 27028 30870
rect 26976 30806 27028 30812
rect 26974 30424 27030 30433
rect 26974 30359 27030 30368
rect 26884 30116 26936 30122
rect 26884 30058 26936 30064
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26700 29776 26752 29782
rect 26700 29718 26752 29724
rect 26608 28688 26660 28694
rect 26528 28648 26608 28676
rect 26240 28484 26292 28490
rect 26240 28426 26292 28432
rect 26332 28484 26384 28490
rect 26332 28426 26384 28432
rect 26148 28416 26200 28422
rect 26148 28358 26200 28364
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 26068 26897 26096 27270
rect 26160 26994 26188 28358
rect 26252 28218 26280 28426
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 26054 26888 26110 26897
rect 26054 26823 26110 26832
rect 26068 26586 26096 26823
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25780 26318 25832 26324
rect 25870 26344 25926 26353
rect 25792 25974 25820 26318
rect 25870 26279 25926 26288
rect 25976 25974 26004 26386
rect 26160 26382 26188 26930
rect 26252 26586 26280 27882
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 26344 27606 26372 27814
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 26436 27538 26464 28358
rect 26528 27577 26556 28648
rect 26608 28630 26660 28636
rect 26712 28558 26740 29718
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26608 28416 26660 28422
rect 26608 28358 26660 28364
rect 26514 27568 26570 27577
rect 26424 27532 26476 27538
rect 26514 27503 26570 27512
rect 26424 27474 26476 27480
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26436 27112 26464 27338
rect 26528 27305 26556 27406
rect 26514 27296 26570 27305
rect 26514 27231 26570 27240
rect 26516 27124 26568 27130
rect 26436 27084 26516 27112
rect 26516 27066 26568 27072
rect 26332 27056 26384 27062
rect 26332 26998 26384 27004
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 25780 25968 25832 25974
rect 25780 25910 25832 25916
rect 25964 25968 26016 25974
rect 25964 25910 26016 25916
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26056 25832 26108 25838
rect 26146 25800 26202 25809
rect 26108 25780 26146 25786
rect 26056 25774 26146 25780
rect 26068 25758 26146 25774
rect 26146 25735 26202 25744
rect 26252 25673 26280 25842
rect 26238 25664 26294 25673
rect 26238 25599 26294 25608
rect 26344 24818 26372 26998
rect 26516 26852 26568 26858
rect 26516 26794 26568 26800
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26436 26246 26464 26318
rect 26424 26240 26476 26246
rect 26424 26182 26476 26188
rect 26436 25106 26464 26182
rect 26528 25362 26556 26794
rect 26516 25356 26568 25362
rect 26516 25298 26568 25304
rect 26514 25120 26570 25129
rect 26436 25078 26514 25106
rect 26514 25055 26570 25064
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26620 24614 26648 28358
rect 26804 28082 26832 29786
rect 26896 29578 26924 30058
rect 26884 29572 26936 29578
rect 26884 29514 26936 29520
rect 26896 28762 26924 29514
rect 26988 29306 27016 30359
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27080 29889 27108 29990
rect 27066 29880 27122 29889
rect 27066 29815 27122 29824
rect 26976 29300 27028 29306
rect 26976 29242 27028 29248
rect 27080 29238 27108 29815
rect 27172 29628 27200 31776
rect 27252 31748 27304 31754
rect 27304 31708 27384 31736
rect 27252 31690 27304 31696
rect 27356 31346 27384 31708
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 27252 31136 27304 31142
rect 27356 31113 27384 31282
rect 27252 31078 27304 31084
rect 27342 31104 27398 31113
rect 27264 29764 27292 31078
rect 27342 31039 27398 31048
rect 27448 30258 27476 32864
rect 27528 32846 27580 32852
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 27540 30802 27568 32302
rect 27632 31822 27660 32914
rect 27724 32910 27752 33254
rect 27816 33153 27844 33458
rect 27894 33280 27950 33289
rect 27894 33215 27950 33224
rect 27802 33144 27858 33153
rect 27908 33114 27936 33215
rect 27802 33079 27858 33088
rect 27896 33108 27948 33114
rect 27896 33050 27948 33056
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27724 31754 27752 32846
rect 27816 32434 27844 32846
rect 27804 32428 27856 32434
rect 28000 32416 28028 33816
rect 28080 33798 28132 33804
rect 28092 33697 28120 33798
rect 28078 33688 28134 33697
rect 28078 33623 28080 33632
rect 28132 33623 28134 33632
rect 28080 33594 28132 33600
rect 27804 32370 27856 32376
rect 27908 32388 28028 32416
rect 27816 31958 27844 32370
rect 27804 31952 27856 31958
rect 27804 31894 27856 31900
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27908 31464 27936 32388
rect 27988 32292 28040 32298
rect 27988 32234 28040 32240
rect 28000 31958 28028 32234
rect 27988 31952 28040 31958
rect 27988 31894 28040 31900
rect 28092 31906 28120 33594
rect 28184 33522 28212 33952
rect 28264 33934 28316 33940
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28276 33318 28304 33934
rect 28368 33833 28396 34002
rect 28644 33946 28672 35226
rect 28736 35086 28764 35974
rect 29012 35698 29040 36518
rect 29090 36479 29146 36488
rect 29092 36168 29144 36174
rect 29090 36136 29092 36145
rect 29144 36136 29146 36145
rect 29090 36071 29146 36080
rect 29196 35834 29224 36790
rect 29288 35834 29316 37062
rect 29472 36825 29500 37590
rect 29564 37466 29592 37606
rect 29552 37460 29604 37466
rect 29552 37402 29604 37408
rect 29748 37346 29776 40326
rect 29552 37324 29604 37330
rect 29552 37266 29604 37272
rect 29656 37318 29776 37346
rect 29458 36816 29514 36825
rect 29368 36780 29420 36786
rect 29564 36802 29592 37266
rect 29656 37262 29684 37318
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 29748 36922 29776 37198
rect 29840 37097 29868 40530
rect 29932 38894 29960 40718
rect 30104 40588 30156 40594
rect 30104 40530 30156 40536
rect 29920 38888 29972 38894
rect 29920 38830 29972 38836
rect 29826 37088 29882 37097
rect 29826 37023 29882 37032
rect 29736 36916 29788 36922
rect 29736 36858 29788 36864
rect 29564 36774 29684 36802
rect 29458 36751 29460 36760
rect 29368 36722 29420 36728
rect 29512 36751 29514 36760
rect 29460 36722 29512 36728
rect 29380 36224 29408 36722
rect 29458 36680 29514 36689
rect 29458 36615 29514 36624
rect 29472 36378 29500 36615
rect 29460 36372 29512 36378
rect 29460 36314 29512 36320
rect 29380 36196 29592 36224
rect 29564 36088 29592 36196
rect 29472 36060 29592 36088
rect 29184 35828 29236 35834
rect 29184 35770 29236 35776
rect 29276 35828 29328 35834
rect 29276 35770 29328 35776
rect 29092 35760 29144 35766
rect 29090 35728 29092 35737
rect 29144 35728 29146 35737
rect 29000 35692 29052 35698
rect 29090 35663 29146 35672
rect 29000 35634 29052 35640
rect 29274 35592 29330 35601
rect 28908 35556 28960 35562
rect 29274 35527 29330 35536
rect 28908 35498 28960 35504
rect 28816 35488 28868 35494
rect 28816 35430 28868 35436
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28828 34066 28856 35430
rect 28920 35154 28948 35498
rect 29092 35488 29144 35494
rect 29092 35430 29144 35436
rect 28908 35148 28960 35154
rect 28908 35090 28960 35096
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 28816 34060 28868 34066
rect 28816 34002 28868 34008
rect 28920 33998 28948 34478
rect 28908 33992 28960 33998
rect 28644 33918 28856 33946
rect 28908 33934 28960 33940
rect 28354 33824 28410 33833
rect 28354 33759 28410 33768
rect 28540 33448 28592 33454
rect 28540 33390 28592 33396
rect 28264 33312 28316 33318
rect 28264 33254 28316 33260
rect 28552 33114 28580 33390
rect 28632 33380 28684 33386
rect 28632 33322 28684 33328
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 28448 32904 28500 32910
rect 28448 32846 28500 32852
rect 28172 32768 28224 32774
rect 28172 32710 28224 32716
rect 28184 32434 28212 32710
rect 28264 32564 28316 32570
rect 28264 32506 28316 32512
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 27632 31436 27936 31464
rect 27632 31346 27660 31436
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27804 31340 27856 31346
rect 27804 31282 27856 31288
rect 27620 31136 27672 31142
rect 27620 31078 27672 31084
rect 27632 30870 27660 31078
rect 27620 30864 27672 30870
rect 27620 30806 27672 30812
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27264 29736 27384 29764
rect 27252 29640 27304 29646
rect 27172 29600 27252 29628
rect 27252 29582 27304 29588
rect 27068 29232 27120 29238
rect 27068 29174 27120 29180
rect 27264 28994 27292 29582
rect 27356 29481 27384 29736
rect 27448 29714 27476 29786
rect 27436 29708 27488 29714
rect 27436 29650 27488 29656
rect 27448 29578 27476 29650
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27342 29472 27398 29481
rect 27342 29407 27398 29416
rect 27448 29238 27476 29514
rect 27540 29306 27568 30738
rect 27724 30569 27752 31282
rect 27710 30560 27766 30569
rect 27710 30495 27766 30504
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27436 29232 27488 29238
rect 27342 29200 27398 29209
rect 27436 29174 27488 29180
rect 27342 29135 27344 29144
rect 27396 29135 27398 29144
rect 27344 29106 27396 29112
rect 27264 28966 27384 28994
rect 26884 28756 26936 28762
rect 26884 28698 26936 28704
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 26884 28620 26936 28626
rect 26884 28562 26936 28568
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 26700 27872 26752 27878
rect 26700 27814 26752 27820
rect 26790 27840 26846 27849
rect 26712 26217 26740 27814
rect 26790 27775 26846 27784
rect 26804 27470 26832 27775
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26804 26246 26832 26726
rect 26896 26586 26924 28562
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 27172 27826 27200 28698
rect 27356 28694 27384 28966
rect 27344 28688 27396 28694
rect 27344 28630 27396 28636
rect 27448 28626 27476 29174
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27540 28762 27568 29106
rect 27528 28756 27580 28762
rect 27528 28698 27580 28704
rect 27436 28620 27488 28626
rect 27436 28562 27488 28568
rect 27540 28506 27568 28698
rect 27448 28478 27568 28506
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27264 28082 27292 28358
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27264 27928 27292 28018
rect 27344 27940 27396 27946
rect 27264 27900 27344 27928
rect 27344 27882 27396 27888
rect 27448 27826 27476 28478
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 28082 27568 28358
rect 27632 28082 27660 29990
rect 27724 29850 27752 30330
rect 27816 29850 27844 31282
rect 27908 31142 27936 31436
rect 27896 31136 27948 31142
rect 27896 31078 27948 31084
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27724 28937 27752 29242
rect 27710 28928 27766 28937
rect 27710 28863 27766 28872
rect 27816 28801 27844 29786
rect 27896 29232 27948 29238
rect 28000 29220 28028 31894
rect 28092 31878 28212 31906
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 28092 31346 28120 31758
rect 28184 31686 28212 31878
rect 28172 31680 28224 31686
rect 28172 31622 28224 31628
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 28170 30968 28226 30977
rect 28170 30903 28172 30912
rect 28224 30903 28226 30912
rect 28172 30874 28224 30880
rect 28172 30388 28224 30394
rect 28172 30330 28224 30336
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 27948 29192 28028 29220
rect 27896 29174 27948 29180
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27802 28792 27858 28801
rect 27802 28727 27858 28736
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27724 28393 27752 28494
rect 27710 28384 27766 28393
rect 27710 28319 27766 28328
rect 27724 28218 27752 28319
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27528 27940 27580 27946
rect 27724 27928 27752 28018
rect 27580 27900 27752 27928
rect 27528 27882 27580 27888
rect 26884 26580 26936 26586
rect 27080 26568 27108 27814
rect 27172 27798 27384 27826
rect 27448 27798 27752 27826
rect 27250 27704 27306 27713
rect 27356 27674 27384 27798
rect 27250 27639 27306 27648
rect 27344 27668 27396 27674
rect 27264 27402 27292 27639
rect 27344 27610 27396 27616
rect 27526 27568 27582 27577
rect 27526 27503 27582 27512
rect 27540 27470 27568 27503
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27252 27396 27304 27402
rect 27252 27338 27304 27344
rect 27160 27328 27212 27334
rect 27160 27270 27212 27276
rect 27250 27296 27306 27305
rect 27172 27130 27200 27270
rect 27356 27282 27384 27406
rect 27306 27254 27384 27282
rect 27250 27231 27306 27240
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27080 26540 27109 26568
rect 26884 26522 26936 26528
rect 27081 26432 27109 26540
rect 27080 26404 27109 26432
rect 26792 26240 26844 26246
rect 26698 26208 26754 26217
rect 26792 26182 26844 26188
rect 26698 26143 26754 26152
rect 26712 25294 26740 26143
rect 26792 25696 26844 25702
rect 26792 25638 26844 25644
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 25884 24274 25912 24550
rect 26349 24410 26556 24426
rect 26332 24404 26556 24410
rect 26384 24398 26556 24404
rect 26332 24346 26384 24352
rect 26528 24290 26556 24398
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 26436 24262 26556 24290
rect 26148 24200 26200 24206
rect 25778 24168 25834 24177
rect 26148 24142 26200 24148
rect 25778 24103 25834 24112
rect 25872 24132 25924 24138
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25700 23730 25728 24006
rect 25792 23905 25820 24103
rect 25872 24074 25924 24080
rect 25778 23896 25834 23905
rect 25884 23866 25912 24074
rect 26160 24070 26188 24142
rect 26148 24064 26200 24070
rect 25962 24032 26018 24041
rect 26148 24006 26200 24012
rect 26286 24064 26338 24070
rect 26338 24012 26377 24018
rect 26286 24006 26377 24012
rect 26298 23990 26377 24006
rect 25962 23967 26018 23976
rect 25778 23831 25834 23840
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25976 23798 26004 23967
rect 26146 23896 26202 23905
rect 26349 23882 26377 23990
rect 26146 23831 26202 23840
rect 26344 23854 26377 23882
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 26056 23724 26108 23730
rect 26160 23712 26188 23831
rect 26108 23684 26188 23712
rect 26056 23666 26108 23672
rect 25964 23588 26016 23594
rect 25964 23530 26016 23536
rect 26056 23588 26108 23594
rect 26056 23530 26108 23536
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25372 21100 25452 21128
rect 25516 22630 25636 22658
rect 25320 21082 25372 21088
rect 25516 21060 25544 22630
rect 25596 22160 25648 22166
rect 25594 22128 25596 22137
rect 25648 22128 25650 22137
rect 25594 22063 25650 22072
rect 25596 22024 25648 22030
rect 25594 21992 25596 22001
rect 25648 21992 25650 22001
rect 25594 21927 25650 21936
rect 25608 21690 25636 21927
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25424 21032 25544 21060
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 24584 20470 24636 20476
rect 24780 20466 24992 20482
rect 24768 20460 24992 20466
rect 24820 20454 24992 20460
rect 24768 20402 24820 20408
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 24768 20324 24820 20330
rect 24768 20266 24820 20272
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24780 20058 24808 20266
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 25134 20224 25190 20233
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24216 19984 24268 19990
rect 24216 19926 24268 19932
rect 24582 19952 24638 19961
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23768 18958 23888 18986
rect 23768 18766 23796 18958
rect 24136 18834 24164 19382
rect 24228 18970 24256 19926
rect 24582 19887 24638 19896
rect 24596 19854 24624 19887
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 23294 18592 23350 18601
rect 23294 18527 23350 18536
rect 23308 18358 23336 18527
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 22928 17604 22980 17610
rect 22928 17546 22980 17552
rect 22940 17338 22968 17546
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 23124 17202 23152 17614
rect 23308 17338 23336 17750
rect 23492 17678 23520 18702
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 18057 23888 18634
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23952 18290 23980 18566
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24044 18086 24072 18702
rect 24136 18426 24164 18770
rect 24320 18766 24348 19722
rect 24412 19514 24440 19790
rect 24400 19508 24452 19514
rect 24400 19450 24452 19456
rect 24688 19378 24716 19790
rect 24780 19786 24808 19994
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24872 19394 24900 19926
rect 24964 19854 24992 20198
rect 25134 20159 25190 20168
rect 25148 19990 25176 20159
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24872 19378 24992 19394
rect 24676 19372 24728 19378
rect 24872 19372 25004 19378
rect 24872 19366 24952 19372
rect 24676 19314 24728 19320
rect 24952 19314 25004 19320
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24398 19000 24454 19009
rect 24596 18970 24624 19110
rect 24398 18935 24454 18944
rect 24492 18964 24544 18970
rect 24412 18766 24440 18935
rect 24492 18906 24544 18912
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24124 18420 24176 18426
rect 24412 18408 24440 18702
rect 24124 18362 24176 18368
rect 24320 18380 24440 18408
rect 24122 18320 24178 18329
rect 24122 18255 24124 18264
rect 24176 18255 24178 18264
rect 24124 18226 24176 18232
rect 24032 18080 24084 18086
rect 23846 18048 23902 18057
rect 24032 18022 24084 18028
rect 23846 17983 23902 17992
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23662 17640 23718 17649
rect 23492 17542 23520 17614
rect 23662 17575 23664 17584
rect 23716 17575 23718 17584
rect 23664 17546 23716 17552
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23124 17066 23152 17138
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 23308 16998 23336 17274
rect 23400 17252 23428 17478
rect 24320 17270 24348 18380
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 23480 17264 23532 17270
rect 23400 17224 23480 17252
rect 24308 17264 24360 17270
rect 23480 17206 23532 17212
rect 23570 17232 23626 17241
rect 24308 17206 24360 17212
rect 23570 17167 23572 17176
rect 23624 17167 23626 17176
rect 23572 17138 23624 17144
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 24412 16726 24440 18226
rect 24504 18154 24532 18906
rect 24688 18902 24716 19314
rect 24952 19236 25004 19242
rect 24952 19178 25004 19184
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24688 18290 24716 18838
rect 24964 18698 24992 19178
rect 25056 18970 25084 19654
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 25148 18873 25176 19790
rect 25134 18864 25190 18873
rect 25134 18799 25190 18808
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 24766 18320 24822 18329
rect 24676 18284 24728 18290
rect 24766 18255 24822 18264
rect 24676 18226 24728 18232
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24492 18148 24544 18154
rect 24492 18090 24544 18096
rect 24504 17610 24532 18090
rect 24596 17678 24624 18158
rect 24688 17882 24716 18226
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24780 17746 24808 18255
rect 25056 18086 25084 18566
rect 25240 18426 25268 20878
rect 25424 20602 25452 21032
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25516 20806 25544 20878
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 20398 25544 20742
rect 25608 20602 25636 20742
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25700 20262 25728 23054
rect 25792 22438 25820 23462
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25884 22545 25912 23054
rect 25870 22536 25926 22545
rect 25870 22471 25872 22480
rect 25924 22471 25926 22480
rect 25872 22442 25924 22448
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25792 22030 25820 22374
rect 25976 22273 26004 23530
rect 26068 23497 26096 23530
rect 26054 23488 26110 23497
rect 26054 23423 26110 23432
rect 26056 23180 26108 23186
rect 26160 23168 26188 23684
rect 26344 23225 26372 23854
rect 26108 23140 26188 23168
rect 26330 23216 26386 23225
rect 26330 23151 26386 23160
rect 26056 23122 26108 23128
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22642 26280 22918
rect 26344 22794 26372 23151
rect 26436 23118 26464 24262
rect 26620 23118 26648 24550
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26712 23118 26740 24278
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26424 22976 26476 22982
rect 26476 22936 26556 22964
rect 26424 22918 26476 22924
rect 26344 22766 26464 22794
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26148 22432 26200 22438
rect 26148 22374 26200 22380
rect 25962 22264 26018 22273
rect 25962 22199 26018 22208
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25778 21584 25834 21593
rect 25884 21554 25912 21830
rect 25778 21519 25780 21528
rect 25832 21519 25834 21528
rect 25872 21548 25924 21554
rect 25780 21490 25832 21496
rect 25872 21490 25924 21496
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25884 21078 25912 21286
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25332 19514 25360 20198
rect 25424 20058 25452 20198
rect 25792 20058 25820 20402
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25780 20052 25832 20058
rect 25780 19994 25832 20000
rect 25884 19938 25912 21014
rect 25976 20534 26004 22199
rect 26056 22160 26108 22166
rect 26056 22102 26108 22108
rect 26068 21622 26096 22102
rect 26160 22098 26188 22374
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 26332 22024 26384 22030
rect 26252 22001 26332 22012
rect 26238 21992 26332 22001
rect 26148 21956 26200 21962
rect 26294 21984 26332 21992
rect 26332 21966 26384 21972
rect 26238 21927 26294 21936
rect 26148 21898 26200 21904
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 26160 20942 26188 21898
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 25964 20528 26016 20534
rect 25964 20470 26016 20476
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25608 19910 25912 19938
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25148 17882 25176 18226
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 25332 17678 25360 19314
rect 25424 18426 25452 19858
rect 25608 19514 25636 19910
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25700 18970 25728 19450
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25502 18728 25558 18737
rect 25502 18663 25558 18672
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25516 18306 25544 18663
rect 25424 18290 25544 18306
rect 25412 18284 25544 18290
rect 25464 18278 25544 18284
rect 25596 18284 25648 18290
rect 25412 18226 25464 18232
rect 25596 18226 25648 18232
rect 25424 17882 25452 18226
rect 25608 17882 25636 18226
rect 25688 18216 25740 18222
rect 25688 18158 25740 18164
rect 25700 17921 25728 18158
rect 25686 17912 25742 17921
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25596 17876 25648 17882
rect 25686 17847 25742 17856
rect 25596 17818 25648 17824
rect 25792 17678 25820 19790
rect 25976 19689 26004 20470
rect 25962 19680 26018 19689
rect 25962 19615 26018 19624
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25976 19009 26004 19246
rect 25962 19000 26018 19009
rect 25962 18935 26018 18944
rect 26068 18714 26096 20878
rect 26160 19922 26188 20878
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20466 26280 20742
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26238 20360 26294 20369
rect 26238 20295 26240 20304
rect 26292 20295 26294 20304
rect 26240 20266 26292 20272
rect 26344 19922 26372 21558
rect 26436 21350 26464 22766
rect 26528 21876 26556 22936
rect 26608 22568 26660 22574
rect 26608 22510 26660 22516
rect 26620 22030 26648 22510
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26528 21848 26648 21876
rect 26620 21554 26648 21848
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26424 21344 26476 21350
rect 26424 21286 26476 21292
rect 26422 21040 26478 21049
rect 26620 21010 26648 21490
rect 26712 21418 26740 22170
rect 26804 22030 26832 25638
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 26896 24177 26924 24210
rect 26882 24168 26938 24177
rect 26882 24103 26938 24112
rect 26976 24132 27028 24138
rect 26976 24074 27028 24080
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26896 22710 26924 24006
rect 26988 23730 27016 24074
rect 27080 23798 27108 26404
rect 27264 26382 27292 26930
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27252 26376 27304 26382
rect 27356 26353 27384 26862
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27252 26318 27304 26324
rect 27342 26344 27398 26353
rect 27342 26279 27398 26288
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27264 25809 27292 26182
rect 27356 25974 27384 26279
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27250 25800 27306 25809
rect 27250 25735 27306 25744
rect 27356 25294 27384 25910
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 27252 25152 27304 25158
rect 27252 25094 27304 25100
rect 27160 24880 27212 24886
rect 27160 24822 27212 24828
rect 27172 24410 27200 24822
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 27068 23792 27120 23798
rect 27068 23734 27120 23740
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26988 23118 27016 23666
rect 27172 23497 27200 24006
rect 27158 23488 27214 23497
rect 27158 23423 27214 23432
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26976 22024 27028 22030
rect 26976 21966 27028 21972
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 26422 20975 26478 20984
rect 26608 21004 26660 21010
rect 26436 20942 26464 20975
rect 26608 20946 26660 20952
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26514 20904 26570 20913
rect 26514 20839 26570 20848
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26436 20058 26464 20334
rect 26424 20052 26476 20058
rect 26424 19994 26476 20000
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26160 19242 26188 19858
rect 26528 19854 26556 20839
rect 26606 20632 26662 20641
rect 26606 20567 26662 20576
rect 26620 19854 26648 20567
rect 26804 20262 26832 21422
rect 26896 21078 26924 21830
rect 26988 21690 27016 21966
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 27080 21690 27108 21830
rect 26976 21684 27028 21690
rect 26976 21626 27028 21632
rect 27068 21684 27120 21690
rect 27068 21626 27120 21632
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26884 21072 26936 21078
rect 26884 21014 26936 21020
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26896 20777 26924 20878
rect 26882 20768 26938 20777
rect 26882 20703 26938 20712
rect 26988 20602 27016 21490
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 27080 20466 27108 21626
rect 27172 21350 27200 22918
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27172 20505 27200 21286
rect 27264 21146 27292 25094
rect 27356 24818 27384 25230
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27448 23798 27476 26726
rect 27540 24954 27568 27406
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27632 26994 27660 27066
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27632 26586 27660 26930
rect 27724 26790 27752 27798
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27620 26580 27672 26586
rect 27620 26522 27672 26528
rect 27632 26450 27660 26522
rect 27620 26444 27672 26450
rect 27816 26432 27844 28086
rect 27908 27402 27936 28970
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 26994 27936 27338
rect 28000 27130 28028 29192
rect 28092 29034 28120 30262
rect 28080 29028 28132 29034
rect 28080 28970 28132 28976
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 28092 27674 28120 28018
rect 28184 27849 28212 30330
rect 28276 29850 28304 32506
rect 28356 32428 28408 32434
rect 28356 32370 28408 32376
rect 28368 31482 28396 32370
rect 28356 31476 28408 31482
rect 28356 31418 28408 31424
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28368 30190 28396 31282
rect 28460 30938 28488 32846
rect 28644 32230 28672 33322
rect 28828 32774 28856 33918
rect 28920 33590 28948 33934
rect 28908 33584 28960 33590
rect 28908 33526 28960 33532
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 28908 32972 28960 32978
rect 28908 32914 28960 32920
rect 28724 32768 28776 32774
rect 28816 32768 28868 32774
rect 28724 32710 28776 32716
rect 28814 32736 28816 32745
rect 28868 32736 28870 32745
rect 28736 32570 28764 32710
rect 28814 32671 28870 32680
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28920 32450 28948 32914
rect 29012 32842 29040 33458
rect 29104 32910 29132 35430
rect 29184 34196 29236 34202
rect 29184 34138 29236 34144
rect 29092 32904 29144 32910
rect 29092 32846 29144 32852
rect 29000 32836 29052 32842
rect 29000 32778 29052 32784
rect 29104 32450 29132 32846
rect 28736 32434 28948 32450
rect 29012 32434 29132 32450
rect 28724 32428 28948 32434
rect 28776 32422 28948 32428
rect 29000 32428 29132 32434
rect 28724 32370 28776 32376
rect 29052 32422 29132 32428
rect 29000 32370 29052 32376
rect 28816 32360 28868 32366
rect 29012 32314 29040 32370
rect 28816 32302 28868 32308
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 31890 28672 32166
rect 28632 31884 28684 31890
rect 28552 31844 28632 31872
rect 28448 30932 28500 30938
rect 28448 30874 28500 30880
rect 28448 30660 28500 30666
rect 28448 30602 28500 30608
rect 28356 30184 28408 30190
rect 28356 30126 28408 30132
rect 28460 30054 28488 30602
rect 28552 30326 28580 31844
rect 28632 31826 28684 31832
rect 28828 31822 28856 32302
rect 28920 32286 29040 32314
rect 28920 31822 28948 32286
rect 29092 31884 29144 31890
rect 29092 31826 29144 31832
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28908 31816 28960 31822
rect 28908 31758 28960 31764
rect 28724 30864 28776 30870
rect 28722 30832 28724 30841
rect 28776 30832 28778 30841
rect 28632 30796 28684 30802
rect 28828 30802 28856 31758
rect 28920 31278 28948 31758
rect 29104 31686 29132 31826
rect 29092 31680 29144 31686
rect 29092 31622 29144 31628
rect 28908 31272 28960 31278
rect 28908 31214 28960 31220
rect 28908 31136 28960 31142
rect 28908 31078 28960 31084
rect 28722 30767 28778 30776
rect 28816 30796 28868 30802
rect 28632 30738 28684 30744
rect 28816 30738 28868 30744
rect 28540 30320 28592 30326
rect 28540 30262 28592 30268
rect 28644 30054 28672 30738
rect 28920 30734 28948 31078
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28828 30394 28856 30534
rect 28816 30388 28868 30394
rect 28816 30330 28868 30336
rect 28920 30258 28948 30670
rect 29196 30376 29224 34138
rect 29288 33114 29316 35527
rect 29368 34536 29420 34542
rect 29368 34478 29420 34484
rect 29276 33108 29328 33114
rect 29276 33050 29328 33056
rect 29274 33008 29330 33017
rect 29380 32978 29408 34478
rect 29472 33998 29500 36060
rect 29552 34740 29604 34746
rect 29656 34728 29684 36774
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 29748 36417 29776 36586
rect 29734 36408 29790 36417
rect 29734 36343 29736 36352
rect 29788 36343 29790 36352
rect 29736 36314 29788 36320
rect 29748 35834 29776 36314
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29604 34700 29684 34728
rect 29552 34682 29604 34688
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 29748 33590 29776 35566
rect 29840 35154 29868 37023
rect 29932 36281 29960 38830
rect 30012 38276 30064 38282
rect 30012 38218 30064 38224
rect 30024 37670 30052 38218
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 30024 37194 30052 37606
rect 30012 37188 30064 37194
rect 30012 37130 30064 37136
rect 30024 36786 30052 37130
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 29918 36272 29974 36281
rect 29918 36207 29974 36216
rect 30116 36174 30144 40530
rect 31036 40526 31064 41958
rect 31208 40928 31260 40934
rect 31208 40870 31260 40876
rect 30748 40520 30800 40526
rect 30748 40462 30800 40468
rect 31024 40520 31076 40526
rect 31024 40462 31076 40468
rect 30380 40452 30432 40458
rect 30380 40394 30432 40400
rect 30392 40050 30420 40394
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30576 40186 30604 40326
rect 30564 40180 30616 40186
rect 30564 40122 30616 40128
rect 30380 40044 30432 40050
rect 30380 39986 30432 39992
rect 30564 39908 30616 39914
rect 30564 39850 30616 39856
rect 30288 38412 30340 38418
rect 30288 38354 30340 38360
rect 30300 37874 30328 38354
rect 30576 37890 30604 39850
rect 30760 38350 30788 40462
rect 30932 39296 30984 39302
rect 30932 39238 30984 39244
rect 30944 39098 30972 39238
rect 30932 39092 30984 39098
rect 30932 39034 30984 39040
rect 31220 38962 31248 40870
rect 31496 40526 31524 41958
rect 31484 40520 31536 40526
rect 31484 40462 31536 40468
rect 31300 40384 31352 40390
rect 31300 40326 31352 40332
rect 31668 40384 31720 40390
rect 31668 40326 31720 40332
rect 31208 38956 31260 38962
rect 31208 38898 31260 38904
rect 30840 38752 30892 38758
rect 30840 38694 30892 38700
rect 30852 38350 30880 38694
rect 31116 38548 31168 38554
rect 31116 38490 31168 38496
rect 30932 38480 30984 38486
rect 30932 38422 30984 38428
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30840 38344 30892 38350
rect 30840 38286 30892 38292
rect 30484 37874 30604 37890
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30472 37868 30604 37874
rect 30524 37862 30604 37868
rect 30472 37810 30524 37816
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30196 36916 30248 36922
rect 30196 36858 30248 36864
rect 30104 36168 30156 36174
rect 30104 36110 30156 36116
rect 30102 35728 30158 35737
rect 30102 35663 30158 35672
rect 30116 35494 30144 35663
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 30012 35216 30064 35222
rect 30012 35158 30064 35164
rect 29828 35148 29880 35154
rect 29828 35090 29880 35096
rect 29840 33810 29868 35090
rect 30024 35018 30052 35158
rect 30208 35086 30236 36858
rect 30392 36582 30420 37062
rect 30380 36576 30432 36582
rect 30286 36544 30342 36553
rect 30380 36518 30432 36524
rect 30286 36479 30342 36488
rect 30300 36174 30328 36479
rect 30288 36168 30340 36174
rect 30288 36110 30340 36116
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30392 35698 30420 35974
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 30012 35012 30064 35018
rect 30012 34954 30064 34960
rect 29920 34944 29972 34950
rect 29920 34886 29972 34892
rect 29932 34746 29960 34886
rect 30300 34746 30328 35566
rect 30852 35086 30880 38286
rect 30944 37262 30972 38422
rect 31128 38350 31156 38490
rect 31024 38344 31076 38350
rect 31024 38286 31076 38292
rect 31116 38344 31168 38350
rect 31116 38286 31168 38292
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 31036 35850 31064 38286
rect 31208 37800 31260 37806
rect 31208 37742 31260 37748
rect 31220 37330 31248 37742
rect 31312 37738 31340 40326
rect 31680 39438 31708 40326
rect 31668 39432 31720 39438
rect 31668 39374 31720 39380
rect 31944 39296 31996 39302
rect 31944 39238 31996 39244
rect 32036 39296 32088 39302
rect 32036 39238 32088 39244
rect 31956 38962 31984 39238
rect 31944 38956 31996 38962
rect 31944 38898 31996 38904
rect 31392 38820 31444 38826
rect 31392 38762 31444 38768
rect 31576 38820 31628 38826
rect 31576 38762 31628 38768
rect 31300 37732 31352 37738
rect 31300 37674 31352 37680
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31116 37256 31168 37262
rect 31116 37198 31168 37204
rect 31128 37126 31156 37198
rect 31116 37120 31168 37126
rect 31116 37062 31168 37068
rect 31128 36145 31156 37062
rect 31312 36854 31340 37674
rect 31404 37262 31432 38762
rect 31588 38554 31616 38762
rect 31576 38548 31628 38554
rect 31576 38490 31628 38496
rect 31956 38282 31984 38898
rect 31944 38276 31996 38282
rect 31944 38218 31996 38224
rect 31760 38208 31812 38214
rect 31760 38150 31812 38156
rect 31852 38208 31904 38214
rect 31852 38150 31904 38156
rect 31392 37256 31444 37262
rect 31392 37198 31444 37204
rect 31300 36848 31352 36854
rect 31300 36790 31352 36796
rect 31114 36136 31170 36145
rect 31114 36071 31170 36080
rect 30944 35822 31064 35850
rect 30944 35290 30972 35822
rect 31024 35760 31076 35766
rect 31024 35702 31076 35708
rect 30932 35284 30984 35290
rect 30932 35226 30984 35232
rect 31036 35154 31064 35702
rect 31024 35148 31076 35154
rect 31024 35090 31076 35096
rect 30840 35080 30892 35086
rect 30840 35022 30892 35028
rect 30656 35012 30708 35018
rect 30656 34954 30708 34960
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 30288 34740 30340 34746
rect 30288 34682 30340 34688
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30576 34066 30604 34342
rect 30668 34066 30696 34954
rect 31404 34950 31432 37198
rect 31772 36718 31800 38150
rect 31864 37670 31892 38150
rect 31852 37664 31904 37670
rect 31852 37606 31904 37612
rect 31760 36712 31812 36718
rect 31760 36654 31812 36660
rect 31760 35488 31812 35494
rect 31760 35430 31812 35436
rect 31772 35154 31800 35430
rect 31760 35148 31812 35154
rect 31760 35090 31812 35096
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31404 34202 31432 34886
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 30564 34060 30616 34066
rect 30564 34002 30616 34008
rect 30656 34060 30708 34066
rect 30656 34002 30708 34008
rect 29840 33782 30052 33810
rect 29736 33584 29788 33590
rect 29736 33526 29788 33532
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29274 32943 29276 32952
rect 29328 32943 29330 32952
rect 29368 32972 29420 32978
rect 29276 32914 29328 32920
rect 29368 32914 29420 32920
rect 29276 32836 29328 32842
rect 29276 32778 29328 32784
rect 29368 32836 29420 32842
rect 29368 32778 29420 32784
rect 29288 30802 29316 32778
rect 29380 32230 29408 32778
rect 29472 32570 29500 33254
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 29460 32564 29512 32570
rect 29460 32506 29512 32512
rect 29368 32224 29420 32230
rect 29368 32166 29420 32172
rect 29380 31754 29408 32166
rect 29564 31822 29592 33050
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29644 32836 29696 32842
rect 29644 32778 29696 32784
rect 29656 32570 29684 32778
rect 29644 32564 29696 32570
rect 29644 32506 29696 32512
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29380 31726 29500 31754
rect 29368 31680 29420 31686
rect 29368 31622 29420 31628
rect 29276 30796 29328 30802
rect 29276 30738 29328 30744
rect 29288 30394 29316 30738
rect 29012 30348 29224 30376
rect 29276 30388 29328 30394
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28722 30152 28778 30161
rect 28722 30087 28778 30096
rect 28736 30054 28764 30087
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28276 28694 28304 29786
rect 28644 29646 28672 29990
rect 28828 29850 28856 30194
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28920 29730 28948 30194
rect 28736 29702 28948 29730
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28632 29640 28684 29646
rect 28632 29582 28684 29588
rect 28264 28688 28316 28694
rect 28264 28630 28316 28636
rect 28264 28484 28316 28490
rect 28460 28472 28488 29582
rect 28538 29336 28594 29345
rect 28736 29306 28764 29702
rect 28814 29472 28870 29481
rect 28814 29407 28870 29416
rect 28538 29271 28594 29280
rect 28724 29300 28776 29306
rect 28552 29238 28580 29271
rect 28724 29242 28776 29248
rect 28540 29232 28592 29238
rect 28540 29174 28592 29180
rect 28540 29028 28592 29034
rect 28540 28970 28592 28976
rect 28632 29028 28684 29034
rect 28632 28970 28684 28976
rect 28552 28626 28580 28970
rect 28644 28937 28672 28970
rect 28630 28928 28686 28937
rect 28630 28863 28686 28872
rect 28736 28762 28764 29242
rect 28828 28762 28856 29407
rect 29012 29152 29040 30348
rect 29276 30330 29328 30336
rect 29184 30252 29236 30258
rect 29184 30194 29236 30200
rect 29090 30016 29146 30025
rect 29090 29951 29146 29960
rect 29104 29850 29132 29951
rect 29092 29844 29144 29850
rect 29092 29786 29144 29792
rect 29092 29572 29144 29578
rect 29196 29560 29224 30194
rect 29144 29532 29224 29560
rect 29092 29514 29144 29520
rect 29104 29306 29132 29514
rect 29288 29458 29316 30330
rect 29380 29889 29408 31622
rect 29472 30258 29500 31726
rect 29564 31346 29592 31758
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 29552 31136 29604 31142
rect 29552 31078 29604 31084
rect 29564 30938 29592 31078
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29366 29880 29422 29889
rect 29366 29815 29422 29824
rect 29196 29430 29316 29458
rect 29196 29306 29224 29430
rect 29274 29336 29330 29345
rect 29092 29300 29144 29306
rect 29092 29242 29144 29248
rect 29184 29300 29236 29306
rect 29274 29271 29330 29280
rect 29184 29242 29236 29248
rect 29092 29164 29144 29170
rect 29012 29124 29092 29152
rect 29092 29106 29144 29112
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28724 28756 28776 28762
rect 28724 28698 28776 28704
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28540 28620 28592 28626
rect 28540 28562 28592 28568
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28316 28444 28488 28472
rect 28264 28426 28316 28432
rect 28356 27940 28408 27946
rect 28356 27882 28408 27888
rect 28170 27840 28226 27849
rect 28170 27775 28226 27784
rect 28080 27668 28132 27674
rect 28080 27610 28132 27616
rect 28092 27470 28120 27610
rect 28184 27470 28212 27775
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27620 26386 27672 26392
rect 27724 26404 27844 26432
rect 27724 25974 27752 26404
rect 27804 26370 27856 26376
rect 28000 26364 28028 26930
rect 28092 26897 28120 27066
rect 28078 26888 28134 26897
rect 28078 26823 28134 26832
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 27856 26336 28028 26364
rect 27804 26312 27856 26318
rect 27988 26240 28040 26246
rect 27988 26182 28040 26188
rect 28000 26042 28028 26182
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 27988 26036 28040 26042
rect 27988 25978 28040 25984
rect 27712 25968 27764 25974
rect 27712 25910 27764 25916
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27540 24410 27568 24754
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27632 24154 27660 25638
rect 27724 24410 27752 25706
rect 27804 24608 27856 24614
rect 27804 24550 27856 24556
rect 27712 24404 27764 24410
rect 27712 24346 27764 24352
rect 27816 24342 27844 24550
rect 27804 24336 27856 24342
rect 27804 24278 27856 24284
rect 27540 24138 27660 24154
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27528 24132 27660 24138
rect 27580 24126 27660 24132
rect 27528 24074 27580 24080
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27632 23730 27660 24126
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27344 23316 27396 23322
rect 27344 23258 27396 23264
rect 27356 21962 27384 23258
rect 27436 23112 27488 23118
rect 27436 23054 27488 23060
rect 27448 22778 27476 23054
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27436 22432 27488 22438
rect 27436 22374 27488 22380
rect 27448 22098 27476 22374
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27356 21146 27384 21626
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27158 20496 27214 20505
rect 27068 20460 27120 20466
rect 27158 20431 27214 20440
rect 27068 20402 27120 20408
rect 27264 20312 27292 20946
rect 27448 20806 27476 21490
rect 27344 20800 27396 20806
rect 27344 20742 27396 20748
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27356 20466 27384 20742
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27344 20324 27396 20330
rect 27264 20284 27344 20312
rect 27344 20266 27396 20272
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 26792 20256 26844 20262
rect 27448 20210 27476 20266
rect 26792 20198 26844 20204
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26148 19236 26200 19242
rect 26148 19178 26200 19184
rect 26160 18902 26188 19178
rect 26238 19136 26294 19145
rect 26238 19071 26294 19080
rect 26148 18896 26200 18902
rect 26148 18838 26200 18844
rect 26252 18766 26280 19071
rect 25884 18686 26096 18714
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26148 18692 26200 18698
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25884 17610 25912 18686
rect 26148 18634 26200 18640
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 25976 17610 26004 18566
rect 26068 18426 26096 18566
rect 26056 18420 26108 18426
rect 26056 18362 26108 18368
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 25504 17604 25556 17610
rect 25504 17546 25556 17552
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 24504 17066 24532 17546
rect 24688 17134 24716 17546
rect 24780 17338 24808 17546
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 25516 16794 25544 17546
rect 25608 17513 25636 17546
rect 25594 17504 25650 17513
rect 25594 17439 25650 17448
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 24400 16720 24452 16726
rect 24400 16662 24452 16668
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23032 16250 23060 16526
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 26068 15502 26096 18022
rect 26160 17882 26188 18634
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26344 17746 26372 19722
rect 26608 19372 26660 19378
rect 26436 19320 26608 19334
rect 26436 19314 26660 19320
rect 26436 19306 26648 19314
rect 26436 18426 26464 19306
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 26712 18154 26740 18566
rect 26700 18148 26752 18154
rect 26700 18090 26752 18096
rect 26712 17785 26740 18090
rect 26804 17882 26832 20198
rect 27264 20182 27476 20210
rect 27264 19990 27292 20182
rect 27342 20088 27398 20097
rect 27540 20058 27568 23462
rect 27632 22642 27660 23666
rect 27816 23662 27844 24142
rect 27908 24138 27936 25978
rect 27986 25392 28042 25401
rect 27986 25327 27988 25336
rect 28040 25327 28042 25336
rect 27988 25298 28040 25304
rect 27896 24132 27948 24138
rect 27896 24074 27948 24080
rect 27908 23866 27936 24074
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27816 23118 27844 23598
rect 27908 23361 27936 23666
rect 27894 23352 27950 23361
rect 27894 23287 27950 23296
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27724 22710 27752 22918
rect 27894 22808 27950 22817
rect 27894 22743 27950 22752
rect 27908 22710 27936 22743
rect 27712 22704 27764 22710
rect 27896 22704 27948 22710
rect 27764 22664 27844 22692
rect 27712 22646 27764 22652
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 22012 27660 22374
rect 27712 22024 27764 22030
rect 27632 21984 27712 22012
rect 27712 21966 27764 21972
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27342 20023 27398 20032
rect 27528 20052 27580 20058
rect 27252 19984 27304 19990
rect 27252 19926 27304 19932
rect 27356 19904 27384 20023
rect 27528 19994 27580 20000
rect 27436 19916 27488 19922
rect 27356 19876 27436 19904
rect 27436 19858 27488 19864
rect 27342 19816 27398 19825
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26976 19780 27028 19786
rect 27342 19751 27398 19760
rect 27436 19780 27488 19786
rect 26976 19722 27028 19728
rect 26896 18970 26924 19722
rect 26988 19334 27016 19722
rect 27356 19446 27384 19751
rect 27436 19722 27488 19728
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 26988 19310 27292 19334
rect 26988 19306 27304 19310
rect 27252 19304 27304 19306
rect 27252 19246 27304 19252
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26976 18896 27028 18902
rect 26976 18838 27028 18844
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26698 17776 26754 17785
rect 26332 17740 26384 17746
rect 26698 17711 26754 17720
rect 26332 17682 26384 17688
rect 26896 16182 26924 18158
rect 26988 17746 27016 18838
rect 27264 18766 27292 19110
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 27264 17678 27292 18566
rect 27448 17678 27476 19722
rect 27632 19446 27660 21830
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27724 21078 27752 21286
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27816 20398 27844 22664
rect 27896 22646 27948 22652
rect 28000 22506 28028 24006
rect 28092 23322 28120 26726
rect 28184 25906 28212 27270
rect 28368 26994 28396 27882
rect 28356 26988 28408 26994
rect 28356 26930 28408 26936
rect 28356 26852 28408 26858
rect 28356 26794 28408 26800
rect 28262 26752 28318 26761
rect 28262 26687 28318 26696
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28184 24818 28212 25842
rect 28276 25770 28304 26687
rect 28264 25764 28316 25770
rect 28264 25706 28316 25712
rect 28264 24948 28316 24954
rect 28264 24890 28316 24896
rect 28276 24818 28304 24890
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28172 24676 28224 24682
rect 28172 24618 28224 24624
rect 28184 24585 28212 24618
rect 28264 24608 28316 24614
rect 28170 24576 28226 24585
rect 28368 24596 28396 26794
rect 28460 26586 28488 28444
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28552 27946 28580 28426
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28644 28082 28672 28358
rect 28632 28076 28684 28082
rect 28632 28018 28684 28024
rect 28540 27940 28592 27946
rect 28540 27882 28592 27888
rect 28736 27674 28764 28494
rect 28724 27668 28776 27674
rect 28724 27610 28776 27616
rect 28724 27532 28776 27538
rect 28724 27474 28776 27480
rect 28632 26784 28684 26790
rect 28632 26726 28684 26732
rect 28448 26580 28500 26586
rect 28448 26522 28500 26528
rect 28644 26353 28672 26726
rect 28736 26518 28764 27474
rect 28816 26988 28868 26994
rect 28816 26930 28868 26936
rect 28724 26512 28776 26518
rect 28724 26454 28776 26460
rect 28630 26344 28686 26353
rect 28448 26308 28500 26314
rect 28630 26279 28686 26288
rect 28448 26250 28500 26256
rect 28460 25838 28488 26250
rect 28540 26240 28592 26246
rect 28724 26240 28776 26246
rect 28540 26182 28592 26188
rect 28644 26200 28724 26228
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28448 24744 28500 24750
rect 28448 24686 28500 24692
rect 28316 24568 28396 24596
rect 28264 24550 28316 24556
rect 28170 24511 28226 24520
rect 28460 23769 28488 24686
rect 28446 23760 28502 23769
rect 28446 23695 28502 23704
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 28080 23316 28132 23322
rect 28080 23258 28132 23264
rect 28080 22704 28132 22710
rect 28080 22646 28132 22652
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27908 22234 27936 22374
rect 28092 22234 28120 22646
rect 27896 22228 27948 22234
rect 27896 22170 27948 22176
rect 28080 22228 28132 22234
rect 28080 22170 28132 22176
rect 28080 22094 28132 22098
rect 28184 22094 28212 23462
rect 28552 23186 28580 26182
rect 28644 25809 28672 26200
rect 28724 26182 28776 26188
rect 28828 26042 28856 26930
rect 28920 26790 28948 28902
rect 29000 28688 29052 28694
rect 29000 28630 29052 28636
rect 29012 27470 29040 28630
rect 29104 28558 29132 29106
rect 29288 29102 29316 29271
rect 29380 29170 29408 29815
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29458 29200 29514 29209
rect 29368 29164 29420 29170
rect 29564 29170 29592 29582
rect 29458 29135 29460 29144
rect 29368 29106 29420 29112
rect 29512 29135 29514 29144
rect 29552 29164 29604 29170
rect 29460 29106 29512 29112
rect 29552 29106 29604 29112
rect 29276 29096 29328 29102
rect 29276 29038 29328 29044
rect 29184 28620 29236 28626
rect 29184 28562 29236 28568
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 28908 26784 28960 26790
rect 28908 26726 28960 26732
rect 28920 26586 28948 26726
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 28908 26444 28960 26450
rect 28908 26386 28960 26392
rect 28920 26217 28948 26386
rect 29196 26364 29224 28562
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29288 26489 29316 28086
rect 29380 27402 29408 29106
rect 29550 29064 29606 29073
rect 29550 28999 29606 29008
rect 29644 29028 29696 29034
rect 29368 27396 29420 27402
rect 29368 27338 29420 27344
rect 29460 27124 29512 27130
rect 29460 27066 29512 27072
rect 29472 26790 29500 27066
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29274 26480 29330 26489
rect 29564 26450 29592 28999
rect 29644 28970 29696 28976
rect 29656 27588 29684 28970
rect 29748 28626 29776 32846
rect 29932 32774 29960 33254
rect 29920 32768 29972 32774
rect 29920 32710 29972 32716
rect 29932 31657 29960 32710
rect 30024 32570 30052 33782
rect 30472 33312 30524 33318
rect 30472 33254 30524 33260
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30012 32564 30064 32570
rect 30012 32506 30064 32512
rect 30392 32434 30420 32846
rect 30012 32428 30064 32434
rect 30380 32428 30432 32434
rect 30012 32370 30064 32376
rect 30300 32388 30380 32416
rect 30024 32042 30052 32370
rect 30024 32014 30236 32042
rect 30104 31952 30156 31958
rect 30104 31894 30156 31900
rect 29918 31648 29974 31657
rect 29918 31583 29974 31592
rect 30116 30734 30144 31894
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 30012 30592 30064 30598
rect 30012 30534 30064 30540
rect 30024 29578 30052 30534
rect 30208 30410 30236 32014
rect 30300 31142 30328 32388
rect 30380 32370 30432 32376
rect 30484 32298 30512 33254
rect 30748 32564 30800 32570
rect 30748 32506 30800 32512
rect 30472 32292 30524 32298
rect 30472 32234 30524 32240
rect 30380 31680 30432 31686
rect 30380 31622 30432 31628
rect 30288 31136 30340 31142
rect 30288 31078 30340 31084
rect 30116 30382 30236 30410
rect 30288 30388 30340 30394
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 29736 28620 29788 28626
rect 29736 28562 29788 28568
rect 29828 27600 29880 27606
rect 29656 27560 29828 27588
rect 29828 27542 29880 27548
rect 29840 27402 29868 27542
rect 29828 27396 29880 27402
rect 29828 27338 29880 27344
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 29748 26858 29776 27270
rect 30024 27130 30052 29514
rect 30116 29102 30144 30382
rect 30288 30330 30340 30336
rect 30196 30320 30248 30326
rect 30196 30262 30248 30268
rect 30208 29753 30236 30262
rect 30194 29744 30250 29753
rect 30194 29679 30250 29688
rect 30300 29646 30328 30330
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30288 29504 30340 29510
rect 30288 29446 30340 29452
rect 30300 29170 30328 29446
rect 30392 29306 30420 31622
rect 30760 31226 30788 32506
rect 31392 32428 31444 32434
rect 31392 32370 31444 32376
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30852 31890 30880 32166
rect 31404 32026 31432 32370
rect 31392 32020 31444 32026
rect 31392 31962 31444 31968
rect 30840 31884 30892 31890
rect 30840 31826 30892 31832
rect 31024 31884 31076 31890
rect 31024 31826 31076 31832
rect 30760 31198 30880 31226
rect 30748 31136 30800 31142
rect 30748 31078 30800 31084
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 30484 30326 30512 30670
rect 30656 30660 30708 30666
rect 30656 30602 30708 30608
rect 30472 30320 30524 30326
rect 30472 30262 30524 30268
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30484 30054 30512 30126
rect 30668 30054 30696 30602
rect 30760 30394 30788 31078
rect 30748 30388 30800 30394
rect 30748 30330 30800 30336
rect 30472 30048 30524 30054
rect 30472 29990 30524 29996
rect 30564 30048 30616 30054
rect 30564 29990 30616 29996
rect 30656 30048 30708 30054
rect 30656 29990 30708 29996
rect 30484 29646 30512 29990
rect 30576 29850 30604 29990
rect 30852 29866 30880 31198
rect 30932 31204 30984 31210
rect 30932 31146 30984 31152
rect 30944 30734 30972 31146
rect 31036 31142 31064 31826
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 31668 31136 31720 31142
rect 31668 31078 31720 31084
rect 31760 31136 31812 31142
rect 31760 31078 31812 31084
rect 30932 30728 30984 30734
rect 31680 30705 31708 31078
rect 30932 30670 30984 30676
rect 31666 30696 31722 30705
rect 30944 30190 30972 30670
rect 31772 30666 31800 31078
rect 31666 30631 31722 30640
rect 31760 30660 31812 30666
rect 31392 30592 31444 30598
rect 31392 30534 31444 30540
rect 31024 30320 31076 30326
rect 31024 30262 31076 30268
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 30564 29844 30616 29850
rect 30564 29786 30616 29792
rect 30668 29838 30880 29866
rect 30562 29744 30618 29753
rect 30668 29714 30696 29838
rect 31036 29730 31064 30262
rect 31404 30258 31432 30534
rect 31680 30274 31708 30631
rect 31760 30602 31812 30608
rect 31680 30258 31800 30274
rect 31392 30252 31444 30258
rect 31576 30252 31628 30258
rect 31392 30194 31444 30200
rect 31496 30212 31576 30240
rect 30562 29679 30618 29688
rect 30656 29708 30708 29714
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30576 29578 30604 29679
rect 30656 29650 30708 29656
rect 31036 29702 31432 29730
rect 30564 29572 30616 29578
rect 30564 29514 30616 29520
rect 30380 29300 30432 29306
rect 30380 29242 30432 29248
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30104 29096 30156 29102
rect 30102 29064 30104 29073
rect 30156 29064 30158 29073
rect 30102 28999 30158 29008
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 30104 27872 30156 27878
rect 30104 27814 30156 27820
rect 30196 27872 30248 27878
rect 30196 27814 30248 27820
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 29736 26852 29788 26858
rect 29736 26794 29788 26800
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 29274 26415 29330 26424
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29840 26382 29868 26726
rect 30116 26625 30144 27814
rect 30208 27674 30236 27814
rect 30196 27668 30248 27674
rect 30196 27610 30248 27616
rect 30300 27470 30328 28494
rect 30392 28490 30420 29242
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30576 28966 30604 29106
rect 30668 29034 30696 29650
rect 30840 29572 30892 29578
rect 30840 29514 30892 29520
rect 30852 29238 30880 29514
rect 30840 29232 30892 29238
rect 30840 29174 30892 29180
rect 31036 29170 31064 29702
rect 31404 29646 31432 29702
rect 31116 29640 31168 29646
rect 31116 29582 31168 29588
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31128 29170 31156 29582
rect 31300 29572 31352 29578
rect 31300 29514 31352 29520
rect 31312 29322 31340 29514
rect 31496 29510 31524 30212
rect 31680 30252 31812 30258
rect 31680 30246 31760 30252
rect 31576 30194 31628 30200
rect 31760 30194 31812 30200
rect 31484 29504 31536 29510
rect 31484 29446 31536 29452
rect 31576 29504 31628 29510
rect 31576 29446 31628 29452
rect 31312 29294 31524 29322
rect 31588 29306 31616 29446
rect 31496 29186 31524 29294
rect 31576 29300 31628 29306
rect 31576 29242 31628 29248
rect 31668 29232 31720 29238
rect 31496 29180 31668 29186
rect 31496 29174 31720 29180
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 31116 29164 31168 29170
rect 31116 29106 31168 29112
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31496 29158 31708 29174
rect 30656 29028 30708 29034
rect 30656 28970 30708 28976
rect 30564 28960 30616 28966
rect 30564 28902 30616 28908
rect 30380 28484 30432 28490
rect 30380 28426 30432 28432
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30288 27464 30340 27470
rect 30288 27406 30340 27412
rect 30392 27033 30420 27950
rect 30576 27606 30604 28902
rect 30668 28082 30696 28970
rect 31036 28558 31064 29106
rect 31128 28762 31156 29106
rect 31116 28756 31168 28762
rect 31116 28698 31168 28704
rect 31404 28558 31432 29106
rect 31496 28665 31524 29158
rect 31772 28994 31800 30194
rect 31864 29850 31892 37606
rect 32048 37126 32076 39238
rect 32312 38344 32364 38350
rect 32312 38286 32364 38292
rect 32404 38344 32456 38350
rect 32404 38286 32456 38292
rect 32128 38276 32180 38282
rect 32128 38218 32180 38224
rect 32036 37120 32088 37126
rect 32036 37062 32088 37068
rect 32140 36961 32168 38218
rect 32324 38049 32352 38286
rect 32310 38040 32366 38049
rect 32416 38010 32444 38286
rect 32310 37975 32366 37984
rect 32404 38004 32456 38010
rect 32404 37946 32456 37952
rect 32692 37806 32720 41958
rect 32784 41818 32812 41958
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 32772 41812 32824 41818
rect 32772 41754 32824 41760
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 33232 39908 33284 39914
rect 33232 39850 33284 39856
rect 33244 38826 33272 39850
rect 33508 39840 33560 39846
rect 33508 39782 33560 39788
rect 33232 38820 33284 38826
rect 33232 38762 33284 38768
rect 32956 38208 33008 38214
rect 32956 38150 33008 38156
rect 32968 38010 32996 38150
rect 32956 38004 33008 38010
rect 32956 37946 33008 37952
rect 33140 37868 33192 37874
rect 33140 37810 33192 37816
rect 32680 37800 32732 37806
rect 32680 37742 32732 37748
rect 32220 37664 32272 37670
rect 32220 37606 32272 37612
rect 32232 37097 32260 37606
rect 33152 37466 33180 37810
rect 33244 37670 33272 38762
rect 33520 38010 33548 39782
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 33600 38752 33652 38758
rect 33600 38694 33652 38700
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 33232 37664 33284 37670
rect 33232 37606 33284 37612
rect 33140 37460 33192 37466
rect 33140 37402 33192 37408
rect 32218 37088 32274 37097
rect 32218 37023 32274 37032
rect 32126 36952 32182 36961
rect 32126 36887 32182 36896
rect 32140 36242 32168 36887
rect 32128 36236 32180 36242
rect 32128 36178 32180 36184
rect 31944 36032 31996 36038
rect 31942 36000 31944 36009
rect 31996 36000 31998 36009
rect 31942 35935 31998 35944
rect 32232 35816 32260 37023
rect 33152 36922 33180 37402
rect 33244 36922 33272 37606
rect 33612 37466 33640 38694
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 33968 37664 34020 37670
rect 33968 37606 34020 37612
rect 33600 37460 33652 37466
rect 33600 37402 33652 37408
rect 33980 37262 34008 37606
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 33968 37256 34020 37262
rect 33322 37224 33378 37233
rect 33968 37198 34020 37204
rect 33322 37159 33378 37168
rect 33336 37126 33364 37159
rect 33324 37120 33376 37126
rect 33324 37062 33376 37068
rect 33140 36916 33192 36922
rect 33140 36858 33192 36864
rect 33232 36916 33284 36922
rect 33232 36858 33284 36864
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 32310 36136 32366 36145
rect 32310 36071 32312 36080
rect 32364 36071 32366 36080
rect 32312 36042 32364 36048
rect 32680 36032 32732 36038
rect 32680 35974 32732 35980
rect 32140 35788 32260 35816
rect 32140 35018 32168 35788
rect 32220 35692 32272 35698
rect 32220 35634 32272 35640
rect 32232 35290 32260 35634
rect 32220 35284 32272 35290
rect 32220 35226 32272 35232
rect 32692 35222 32720 35974
rect 33060 35834 33088 36178
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 32680 35216 32732 35222
rect 32680 35158 32732 35164
rect 32312 35080 32364 35086
rect 32312 35022 32364 35028
rect 32128 35012 32180 35018
rect 32128 34954 32180 34960
rect 32324 34746 32352 35022
rect 32312 34740 32364 34746
rect 32312 34682 32364 34688
rect 32220 32564 32272 32570
rect 32220 32506 32272 32512
rect 32128 32224 32180 32230
rect 32128 32166 32180 32172
rect 32140 31929 32168 32166
rect 32126 31920 32182 31929
rect 32232 31890 32260 32506
rect 33048 32496 33100 32502
rect 33048 32438 33100 32444
rect 32772 32224 32824 32230
rect 32772 32166 32824 32172
rect 32126 31855 32182 31864
rect 32220 31884 32272 31890
rect 32220 31826 32272 31832
rect 32404 31816 32456 31822
rect 32404 31758 32456 31764
rect 32128 31680 32180 31686
rect 32128 31622 32180 31628
rect 32220 31680 32272 31686
rect 32220 31622 32272 31628
rect 32140 31346 32168 31622
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32232 30734 32260 31622
rect 32416 30938 32444 31758
rect 32404 30932 32456 30938
rect 32404 30874 32456 30880
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 31944 30592 31996 30598
rect 31944 30534 31996 30540
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 31956 30326 31984 30534
rect 31944 30320 31996 30326
rect 31944 30262 31996 30268
rect 32220 30252 32272 30258
rect 32220 30194 32272 30200
rect 32036 30184 32088 30190
rect 32036 30126 32088 30132
rect 31944 30048 31996 30054
rect 31944 29990 31996 29996
rect 31852 29844 31904 29850
rect 31852 29786 31904 29792
rect 31956 29617 31984 29990
rect 31942 29608 31998 29617
rect 32048 29578 32076 30126
rect 32232 29782 32260 30194
rect 32324 30054 32352 30534
rect 32312 30048 32364 30054
rect 32312 29990 32364 29996
rect 32220 29776 32272 29782
rect 32220 29718 32272 29724
rect 31942 29543 31998 29552
rect 32036 29572 32088 29578
rect 32036 29514 32088 29520
rect 31680 28966 31800 28994
rect 31482 28656 31538 28665
rect 31482 28591 31538 28600
rect 31024 28552 31076 28558
rect 31392 28552 31444 28558
rect 31024 28494 31076 28500
rect 31390 28520 31392 28529
rect 31444 28520 31446 28529
rect 30748 28484 30800 28490
rect 30748 28426 30800 28432
rect 30760 28218 30788 28426
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30656 28076 30708 28082
rect 30656 28018 30708 28024
rect 31036 27674 31064 28494
rect 31390 28455 31446 28464
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 31208 27668 31260 27674
rect 31208 27610 31260 27616
rect 30564 27600 30616 27606
rect 30616 27560 30788 27588
rect 30564 27542 30616 27548
rect 30760 27470 30788 27560
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30932 27464 30984 27470
rect 30984 27424 31156 27452
rect 30932 27406 30984 27412
rect 30668 27282 30696 27406
rect 31024 27328 31076 27334
rect 30746 27296 30802 27305
rect 30668 27254 30746 27282
rect 31024 27270 31076 27276
rect 30746 27231 30802 27240
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 30378 27024 30434 27033
rect 30944 26994 30972 27066
rect 31036 26994 31064 27270
rect 31128 27130 31156 27424
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 30378 26959 30434 26968
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 30196 26920 30248 26926
rect 30196 26862 30248 26868
rect 30102 26616 30158 26625
rect 30102 26551 30158 26560
rect 30208 26382 30236 26862
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30392 26450 30420 26726
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 29828 26376 29880 26382
rect 29196 26336 29408 26364
rect 29000 26240 29052 26246
rect 28906 26208 28962 26217
rect 29000 26182 29052 26188
rect 29092 26240 29144 26246
rect 29092 26182 29144 26188
rect 28906 26143 28962 26152
rect 28816 26036 28868 26042
rect 28816 25978 28868 25984
rect 28630 25800 28686 25809
rect 28630 25735 28686 25744
rect 28724 25764 28776 25770
rect 28724 25706 28776 25712
rect 28736 24886 28764 25706
rect 28828 24954 28856 25978
rect 28908 25832 28960 25838
rect 28908 25774 28960 25780
rect 28920 25362 28948 25774
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 29012 25242 29040 26182
rect 29104 25770 29132 26182
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 29184 25764 29236 25770
rect 29184 25706 29236 25712
rect 29196 25276 29224 25706
rect 29104 25272 29224 25276
rect 28920 25214 29040 25242
rect 29092 25266 29224 25272
rect 29144 25248 29224 25266
rect 29276 25288 29328 25294
rect 29380 25276 29408 26336
rect 29828 26318 29880 26324
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 30196 26376 30248 26382
rect 30196 26318 30248 26324
rect 29552 26240 29604 26246
rect 29932 26234 29960 26318
rect 29552 26182 29604 26188
rect 29656 26206 29960 26234
rect 29564 26042 29592 26182
rect 29552 26036 29604 26042
rect 29552 25978 29604 25984
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 29472 25430 29500 25910
rect 29552 25764 29604 25770
rect 29656 25752 29684 26206
rect 30104 25900 30156 25906
rect 30104 25842 30156 25848
rect 29604 25724 29684 25752
rect 29552 25706 29604 25712
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 29460 25424 29512 25430
rect 29460 25366 29512 25372
rect 29552 25424 29604 25430
rect 29552 25366 29604 25372
rect 29328 25248 29408 25276
rect 29276 25230 29328 25236
rect 28816 24948 28868 24954
rect 28816 24890 28868 24896
rect 28724 24880 28776 24886
rect 28724 24822 28776 24828
rect 28920 24818 28948 25214
rect 29092 25208 29144 25214
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24936 29132 25094
rect 29012 24908 29132 24936
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 29012 24682 29040 24908
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 28632 24676 28684 24682
rect 28632 24618 28684 24624
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 28540 23180 28592 23186
rect 28540 23122 28592 23128
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28538 23080 28594 23089
rect 28276 22953 28304 23054
rect 28538 23015 28594 23024
rect 28356 22976 28408 22982
rect 28262 22944 28318 22953
rect 28356 22918 28408 22924
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 28262 22879 28318 22888
rect 28276 22642 28304 22879
rect 28368 22642 28396 22918
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28368 22545 28396 22578
rect 28354 22536 28410 22545
rect 28354 22471 28410 22480
rect 28460 22438 28488 22918
rect 28552 22778 28580 23015
rect 28540 22772 28592 22778
rect 28540 22714 28592 22720
rect 28448 22432 28500 22438
rect 28552 22409 28580 22714
rect 28644 22642 28672 24618
rect 28724 24608 28776 24614
rect 28776 24568 28856 24596
rect 28724 24550 28776 24556
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28632 22432 28684 22438
rect 28448 22374 28500 22380
rect 28538 22400 28594 22409
rect 28460 22094 28488 22374
rect 28632 22374 28684 22380
rect 28538 22335 28594 22344
rect 28080 22092 28212 22094
rect 28132 22066 28212 22092
rect 28368 22066 28488 22094
rect 28080 22034 28132 22040
rect 28368 22030 28396 22066
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 27988 21888 28040 21894
rect 28264 21888 28316 21894
rect 27988 21830 28040 21836
rect 28092 21848 28264 21876
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27620 19440 27672 19446
rect 27620 19382 27672 19388
rect 27724 19174 27752 19654
rect 27816 19310 27844 20198
rect 27908 20058 27936 20470
rect 27896 20052 27948 20058
rect 27896 19994 27948 20000
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 28000 18766 28028 21830
rect 28092 21146 28120 21848
rect 28264 21830 28316 21836
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28184 21146 28212 21286
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28276 20602 28304 21490
rect 28356 21412 28408 21418
rect 28356 21354 28408 21360
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 28262 20496 28318 20505
rect 28262 20431 28264 20440
rect 28316 20431 28318 20440
rect 28264 20402 28316 20408
rect 28172 20392 28224 20398
rect 28224 20340 28304 20346
rect 28172 20334 28304 20340
rect 28184 20318 28304 20334
rect 28080 20256 28132 20262
rect 28078 20224 28080 20233
rect 28172 20256 28224 20262
rect 28132 20224 28134 20233
rect 28172 20198 28224 20204
rect 28078 20159 28134 20168
rect 28092 19854 28120 20159
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28184 19334 28212 20198
rect 28276 19854 28304 20318
rect 28368 20058 28396 21354
rect 28460 20466 28488 21830
rect 28552 21593 28580 21898
rect 28538 21584 28594 21593
rect 28644 21554 28672 22374
rect 28736 21554 28764 24278
rect 28828 22030 28856 24568
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 29012 23866 29040 24346
rect 29104 24138 29132 24686
rect 29092 24132 29144 24138
rect 29092 24074 29144 24080
rect 29460 24132 29512 24138
rect 29460 24074 29512 24080
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29472 23662 29500 24074
rect 29564 23798 29592 25366
rect 29552 23792 29604 23798
rect 29552 23734 29604 23740
rect 29460 23656 29512 23662
rect 29460 23598 29512 23604
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28538 21519 28594 21528
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28552 20466 28580 21422
rect 28644 20942 28672 21490
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28092 19306 28212 19334
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27988 18760 28040 18766
rect 27988 18702 28040 18708
rect 27632 18290 27660 18702
rect 28092 18426 28120 19306
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28080 18420 28132 18426
rect 28080 18362 28132 18368
rect 28184 18358 28212 19110
rect 28172 18352 28224 18358
rect 28172 18294 28224 18300
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 28368 16182 28396 19654
rect 28460 19514 28488 20198
rect 28644 19514 28672 20742
rect 28736 19786 28764 21490
rect 28828 20942 28856 21966
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28816 19712 28868 19718
rect 28816 19654 28868 19660
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 28356 16176 28408 16182
rect 28356 16118 28408 16124
rect 28828 15910 28856 19654
rect 28920 18698 28948 20878
rect 29104 20466 29132 21830
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29104 19854 29132 20402
rect 29196 19922 29224 21286
rect 29472 20942 29500 23598
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29184 19916 29236 19922
rect 29184 19858 29236 19864
rect 29092 19848 29144 19854
rect 29656 19825 29684 25434
rect 29736 25288 29788 25294
rect 30012 25288 30064 25294
rect 29736 25230 29788 25236
rect 30010 25256 30012 25265
rect 30064 25256 30066 25265
rect 29748 25129 29776 25230
rect 30010 25191 30066 25200
rect 29734 25120 29790 25129
rect 29734 25055 29790 25064
rect 30024 23866 30052 25191
rect 30116 24954 30144 25842
rect 30208 25226 30236 26318
rect 30288 26308 30340 26314
rect 30288 26250 30340 26256
rect 30196 25220 30248 25226
rect 30196 25162 30248 25168
rect 30104 24948 30156 24954
rect 30104 24890 30156 24896
rect 30208 24410 30236 25162
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 30012 23860 30064 23866
rect 30012 23802 30064 23808
rect 30300 22094 30328 26250
rect 30576 25226 30604 26726
rect 30668 26382 30696 26726
rect 30760 26586 30788 26930
rect 30748 26580 30800 26586
rect 30748 26522 30800 26528
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30852 25702 30880 26930
rect 31128 26586 31156 27066
rect 31220 26994 31248 27610
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 31220 26382 31248 26930
rect 31312 26586 31340 26930
rect 31496 26790 31524 27406
rect 31484 26784 31536 26790
rect 31484 26726 31536 26732
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 30932 26376 30984 26382
rect 30932 26318 30984 26324
rect 31208 26376 31260 26382
rect 31208 26318 31260 26324
rect 30944 25945 30972 26318
rect 31680 26234 31708 28966
rect 32048 28626 32076 29514
rect 32036 28620 32088 28626
rect 32036 28562 32088 28568
rect 32128 28484 32180 28490
rect 32128 28426 32180 28432
rect 32140 28218 32168 28426
rect 32128 28212 32180 28218
rect 32128 28154 32180 28160
rect 32128 28076 32180 28082
rect 32128 28018 32180 28024
rect 31760 27600 31812 27606
rect 31758 27568 31760 27577
rect 31812 27568 31814 27577
rect 31758 27503 31814 27512
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 31758 27160 31814 27169
rect 31814 27118 31892 27146
rect 31758 27095 31814 27104
rect 31864 27062 31892 27118
rect 31852 27056 31904 27062
rect 31852 26998 31904 27004
rect 31956 26994 31984 27406
rect 32140 26994 32168 28018
rect 32680 27464 32732 27470
rect 32680 27406 32732 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32220 27328 32272 27334
rect 32220 27270 32272 27276
rect 32232 26994 32260 27270
rect 31944 26988 31996 26994
rect 31944 26930 31996 26936
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 31852 26852 31904 26858
rect 31852 26794 31904 26800
rect 31588 26206 31708 26234
rect 30930 25936 30986 25945
rect 30930 25871 30986 25880
rect 30944 25770 30972 25871
rect 31116 25832 31168 25838
rect 31116 25774 31168 25780
rect 30932 25764 30984 25770
rect 30932 25706 30984 25712
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 31128 25498 31156 25774
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 31588 25294 31616 26206
rect 31864 25974 31892 26794
rect 32036 26784 32088 26790
rect 32036 26726 32088 26732
rect 32048 26314 32076 26726
rect 32140 26314 32168 26930
rect 32036 26308 32088 26314
rect 32036 26250 32088 26256
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 31852 25968 31904 25974
rect 31852 25910 31904 25916
rect 32140 25906 32168 26250
rect 32600 26042 32628 27338
rect 32692 27305 32720 27406
rect 32678 27296 32734 27305
rect 32678 27231 32734 27240
rect 32784 26518 32812 32166
rect 33060 32026 33088 32438
rect 33048 32020 33100 32026
rect 33048 31962 33100 31968
rect 33244 29306 33272 36858
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 33520 30394 33548 30670
rect 33508 30388 33560 30394
rect 33508 30330 33560 30336
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 32956 28756 33008 28762
rect 32956 28698 33008 28704
rect 32968 27402 32996 28698
rect 33060 28626 33088 29038
rect 33428 28762 33456 29106
rect 33692 29028 33744 29034
rect 33692 28970 33744 28976
rect 34060 29028 34112 29034
rect 34060 28970 34112 28976
rect 33508 28960 33560 28966
rect 33508 28902 33560 28908
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 33520 28558 33548 28902
rect 33508 28552 33560 28558
rect 33560 28512 33640 28540
rect 33508 28494 33560 28500
rect 33232 28416 33284 28422
rect 33232 28358 33284 28364
rect 33508 28416 33560 28422
rect 33508 28358 33560 28364
rect 33048 27600 33100 27606
rect 33046 27568 33048 27577
rect 33100 27568 33102 27577
rect 33244 27538 33272 28358
rect 33520 28082 33548 28358
rect 33612 28082 33640 28512
rect 33704 28082 33732 28970
rect 33968 28484 34020 28490
rect 33968 28426 34020 28432
rect 33980 28218 34008 28426
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 33508 28076 33560 28082
rect 33508 28018 33560 28024
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33692 28076 33744 28082
rect 33692 28018 33744 28024
rect 34072 27674 34100 28970
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 36280 28490 36308 29514
rect 36268 28484 36320 28490
rect 36268 28426 36320 28432
rect 36280 28082 36308 28426
rect 36268 28076 36320 28082
rect 36268 28018 36320 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34060 27668 34112 27674
rect 34060 27610 34112 27616
rect 33046 27503 33102 27512
rect 33232 27532 33284 27538
rect 33232 27474 33284 27480
rect 34072 27402 34100 27610
rect 32956 27396 33008 27402
rect 32956 27338 33008 27344
rect 34060 27396 34112 27402
rect 34060 27338 34112 27344
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33796 27130 33824 27270
rect 34072 27130 34100 27338
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 34060 27124 34112 27130
rect 34060 27066 34112 27072
rect 33876 26920 33928 26926
rect 33876 26862 33928 26868
rect 33888 26586 33916 26862
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 32772 26512 32824 26518
rect 32772 26454 32824 26460
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32494 25936 32550 25945
rect 32128 25900 32180 25906
rect 32494 25871 32550 25880
rect 32128 25842 32180 25848
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 30564 25220 30616 25226
rect 30564 25162 30616 25168
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31668 23792 31720 23798
rect 31496 23752 31668 23780
rect 31496 23633 31524 23752
rect 31772 23780 31800 25094
rect 31944 24608 31996 24614
rect 31944 24550 31996 24556
rect 31956 24410 31984 24550
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 32140 24274 32168 25842
rect 32508 25498 32536 25871
rect 32954 25528 33010 25537
rect 32496 25492 32548 25498
rect 32954 25463 32956 25472
rect 32496 25434 32548 25440
rect 33008 25463 33010 25472
rect 32956 25434 33008 25440
rect 32680 25356 32732 25362
rect 32680 25298 32732 25304
rect 32220 25152 32272 25158
rect 32220 25094 32272 25100
rect 32232 24818 32260 25094
rect 32692 24954 32720 25298
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 32968 24818 32996 25434
rect 33888 24954 33916 26522
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 36464 24818 36492 41958
rect 37660 38418 37688 41958
rect 43812 39364 43864 39370
rect 43812 39306 43864 39312
rect 43536 39296 43588 39302
rect 43824 39273 43852 39306
rect 43536 39238 43588 39244
rect 43810 39264 43866 39273
rect 37648 38412 37700 38418
rect 37648 38354 37700 38360
rect 42154 31240 42210 31249
rect 42154 31175 42210 31184
rect 42168 28694 42196 31175
rect 43548 28762 43576 39238
rect 43810 39199 43866 39208
rect 43536 28756 43588 28762
rect 43536 28698 43588 28704
rect 42156 28688 42208 28694
rect 42156 28630 42208 28636
rect 41880 28552 41932 28558
rect 41880 28494 41932 28500
rect 42340 28552 42392 28558
rect 42340 28494 42392 28500
rect 42800 28552 42852 28558
rect 42800 28494 42852 28500
rect 41892 28422 41920 28494
rect 41880 28416 41932 28422
rect 41880 28358 41932 28364
rect 41892 28218 41920 28358
rect 42352 28218 42380 28494
rect 41880 28212 41932 28218
rect 41880 28154 41932 28160
rect 42340 28212 42392 28218
rect 42340 28154 42392 28160
rect 42812 28150 42840 28494
rect 42984 28484 43036 28490
rect 42984 28426 43036 28432
rect 42996 28150 43024 28426
rect 43260 28416 43312 28422
rect 43260 28358 43312 28364
rect 42800 28144 42852 28150
rect 42800 28086 42852 28092
rect 42984 28144 43036 28150
rect 42984 28086 43036 28092
rect 43272 27878 43300 28358
rect 43810 28112 43866 28121
rect 43810 28047 43812 28056
rect 43864 28047 43866 28056
rect 43812 28018 43864 28024
rect 43260 27872 43312 27878
rect 43260 27814 43312 27820
rect 40682 27432 40738 27441
rect 40682 27367 40738 27376
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 33600 24812 33652 24818
rect 33600 24754 33652 24760
rect 36452 24812 36504 24818
rect 36452 24754 36504 24760
rect 32404 24744 32456 24750
rect 32404 24686 32456 24692
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 31720 23752 31800 23780
rect 31668 23734 31720 23740
rect 32324 23730 32352 24006
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 31482 23624 31538 23633
rect 31482 23559 31538 23568
rect 32324 23186 32352 23666
rect 32416 23322 32444 24686
rect 33140 23520 33192 23526
rect 33140 23462 33192 23468
rect 33152 23322 33180 23462
rect 33612 23322 33640 24754
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33796 24410 33824 24550
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33784 24064 33836 24070
rect 33784 24006 33836 24012
rect 33796 23866 33824 24006
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 32404 23316 32456 23322
rect 32404 23258 32456 23264
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 33600 23316 33652 23322
rect 33600 23258 33652 23264
rect 32312 23180 32364 23186
rect 32312 23122 32364 23128
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 30208 22066 30328 22094
rect 30208 21729 30236 22066
rect 30194 21720 30250 21729
rect 30194 21655 30250 21664
rect 30208 21146 30236 21655
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 29092 19790 29144 19796
rect 29642 19816 29698 19825
rect 29642 19751 29698 19760
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 29090 19000 29146 19009
rect 34934 19003 35242 19012
rect 29090 18935 29092 18944
rect 29144 18935 29146 18944
rect 29092 18906 29144 18912
rect 28908 18692 28960 18698
rect 28908 18634 28960 18640
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 40696 5817 40724 27367
rect 43260 25492 43312 25498
rect 43260 25434 43312 25440
rect 43272 17338 43300 25434
rect 43260 17332 43312 17338
rect 43260 17274 43312 17280
rect 43168 17196 43220 17202
rect 43168 17138 43220 17144
rect 43180 16969 43208 17138
rect 43166 16960 43222 16969
rect 43166 16895 43222 16904
rect 40682 5808 40738 5817
rect 40682 5743 40738 5752
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1228 4457 1256 4626
rect 1214 4448 1270 4457
rect 1214 4383 1270 4392
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 3146 4040 3202 4049
rect 3146 3975 3202 3984
rect 3160 3738 3188 3975
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 1216 3596 1268 3602
rect 1216 3538 1268 3544
rect 1228 3369 1256 3538
rect 1214 3360 1270 3369
rect 1214 3295 1270 3304
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 24674 2680 24730 2689
rect 34934 2683 35242 2692
rect 24674 2615 24676 2624
rect 24728 2615 24730 2624
rect 24676 2586 24728 2592
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 22480 800 22508 2450
rect 22466 0 22522 800
<< via2 >>
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 938 41384 994 41440
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 938 40296 994 40352
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 1214 39208 1270 39264
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 1214 38120 1270 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1214 37068 1216 37088
rect 1216 37068 1268 37088
rect 1268 37068 1270 37088
rect 1214 37032 1270 37068
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 938 35944 994 36000
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 938 34856 994 34912
rect 938 33768 994 33824
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 2686 32952 2742 33008
rect 938 32716 940 32736
rect 940 32716 992 32736
rect 992 32716 994 32736
rect 938 32680 994 32716
rect 1490 31592 1546 31648
rect 1214 30504 1270 30560
rect 1214 29416 1270 29472
rect 1490 29144 1546 29200
rect 1214 28328 1270 28384
rect 1214 27240 1270 27296
rect 1582 28056 1638 28112
rect 2870 30504 2926 30560
rect 2962 30368 3018 30424
rect 3330 30660 3386 30696
rect 3330 30640 3332 30660
rect 3332 30640 3384 30660
rect 3384 30640 3386 30660
rect 2318 29280 2374 29336
rect 2226 28736 2282 28792
rect 1674 27104 1730 27160
rect 3054 29416 3110 29472
rect 3330 29280 3386 29336
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4158 31864 4214 31920
rect 3606 28600 3662 28656
rect 3238 28364 3240 28384
rect 3240 28364 3292 28384
rect 3292 28364 3294 28384
rect 3238 28328 3294 28364
rect 2962 27920 3018 27976
rect 1582 26324 1584 26344
rect 1584 26324 1636 26344
rect 1636 26324 1638 26344
rect 1582 26288 1638 26324
rect 1858 26152 1914 26208
rect 1214 23976 1270 24032
rect 1214 22888 1270 22944
rect 1214 21800 1270 21856
rect 1214 20712 1270 20768
rect 1214 19624 1270 19680
rect 1582 24248 1638 24304
rect 2042 22072 2098 22128
rect 1950 21564 1952 21584
rect 1952 21564 2004 21584
rect 2004 21564 2006 21584
rect 1950 21528 2006 21564
rect 1214 18536 1270 18592
rect 1214 17448 1270 17504
rect 1214 16360 1270 16416
rect 1214 15272 1270 15328
rect 1214 14184 1270 14240
rect 2502 20984 2558 21040
rect 2502 20712 2558 20768
rect 2778 25064 2834 25120
rect 3330 26152 3386 26208
rect 3422 25200 3478 25256
rect 3054 23024 3110 23080
rect 2962 22888 3018 22944
rect 3330 23160 3386 23216
rect 3054 22616 3110 22672
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4894 30676 4896 30696
rect 4896 30676 4948 30696
rect 4948 30676 4950 30696
rect 4894 30640 4950 30676
rect 4802 30388 4858 30424
rect 4802 30368 4804 30388
rect 4804 30368 4856 30388
rect 4856 30368 4858 30388
rect 4526 30232 4582 30288
rect 5538 31320 5594 31376
rect 5170 30368 5226 30424
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4066 29688 4122 29744
rect 4986 30232 5042 30288
rect 5446 30504 5502 30560
rect 3974 28756 4030 28792
rect 3974 28736 3976 28756
rect 3976 28736 4028 28756
rect 4028 28736 4030 28756
rect 4526 29164 4582 29200
rect 4526 29144 4528 29164
rect 4528 29144 4580 29164
rect 4580 29144 4582 29164
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 3974 28192 4030 28248
rect 4434 28484 4490 28520
rect 4434 28464 4436 28484
rect 4436 28464 4488 28484
rect 4488 28464 4490 28484
rect 4802 28736 4858 28792
rect 4986 29164 5042 29200
rect 4986 29144 4988 29164
rect 4988 29144 5040 29164
rect 5040 29144 5042 29164
rect 5354 29688 5410 29744
rect 5630 28756 5686 28792
rect 5630 28736 5632 28756
rect 5632 28736 5684 28756
rect 5684 28736 5686 28756
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4342 26968 4398 27024
rect 4342 26868 4344 26888
rect 4344 26868 4396 26888
rect 4396 26868 4398 26888
rect 4342 26832 4398 26868
rect 4802 26988 4858 27024
rect 4802 26968 4804 26988
rect 4804 26968 4856 26988
rect 4856 26968 4858 26988
rect 4802 26696 4858 26752
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4434 25744 4490 25800
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 3606 21936 3662 21992
rect 3054 20304 3110 20360
rect 3054 19216 3110 19272
rect 3422 20476 3424 20496
rect 3424 20476 3476 20496
rect 3476 20476 3478 20496
rect 3422 20440 3478 20476
rect 4710 24928 4766 24984
rect 5630 28364 5632 28384
rect 5632 28364 5684 28384
rect 5684 28364 5686 28384
rect 5630 28328 5686 28364
rect 5262 27240 5318 27296
rect 5538 27784 5594 27840
rect 5538 27240 5594 27296
rect 5354 26832 5410 26888
rect 5262 26696 5318 26752
rect 5170 26460 5172 26480
rect 5172 26460 5224 26480
rect 5224 26460 5226 26480
rect 5170 26424 5226 26460
rect 5262 25900 5318 25936
rect 5262 25880 5264 25900
rect 5264 25880 5316 25900
rect 5316 25880 5318 25900
rect 5170 25472 5226 25528
rect 4618 24656 4674 24712
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4158 23840 4214 23896
rect 4526 23568 4582 23624
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4710 23296 4766 23352
rect 4250 22480 4306 22536
rect 3882 21664 3938 21720
rect 3698 20848 3754 20904
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4802 22752 4858 22808
rect 5906 34448 5962 34504
rect 6182 34176 6238 34232
rect 5906 26832 5962 26888
rect 5814 26424 5870 26480
rect 5814 25336 5870 25392
rect 4250 21936 4306 21992
rect 4158 21800 4214 21856
rect 4250 21392 4306 21448
rect 4526 21664 4582 21720
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4158 20576 4214 20632
rect 4526 20440 4582 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 5078 23840 5134 23896
rect 5262 23840 5318 23896
rect 5262 23432 5318 23488
rect 5538 24112 5594 24168
rect 5538 23568 5594 23624
rect 5170 22480 5226 22536
rect 5078 22344 5134 22400
rect 4986 22072 5042 22128
rect 4986 21956 5042 21992
rect 4986 21936 4988 21956
rect 4988 21936 5040 21956
rect 5040 21936 5042 21956
rect 4710 20712 4766 20768
rect 4894 21256 4950 21312
rect 4894 20984 4950 21040
rect 4894 20168 4950 20224
rect 5354 22752 5410 22808
rect 5354 22480 5410 22536
rect 5814 25064 5870 25120
rect 6458 30232 6514 30288
rect 6366 28736 6422 28792
rect 6366 28464 6422 28520
rect 6366 27376 6422 27432
rect 5998 25608 6054 25664
rect 5906 24384 5962 24440
rect 8298 36080 8354 36136
rect 7286 29416 7342 29472
rect 6642 27920 6698 27976
rect 6458 26016 6514 26072
rect 6366 25608 6422 25664
rect 7010 27784 7066 27840
rect 6734 27376 6790 27432
rect 7194 27104 7250 27160
rect 6734 26288 6790 26344
rect 6550 25608 6606 25664
rect 6642 25336 6698 25392
rect 6458 25100 6460 25120
rect 6460 25100 6512 25120
rect 6512 25100 6514 25120
rect 6458 25064 6514 25100
rect 6550 24928 6606 24984
rect 6274 24656 6330 24712
rect 6366 24520 6422 24576
rect 8574 34196 8630 34232
rect 8574 34176 8576 34196
rect 8576 34176 8628 34196
rect 8628 34176 8630 34196
rect 9310 36116 9312 36136
rect 9312 36116 9364 36136
rect 9364 36116 9366 36136
rect 9310 36080 9366 36116
rect 9678 35692 9734 35728
rect 9678 35672 9680 35692
rect 9680 35672 9732 35692
rect 9732 35672 9734 35692
rect 9678 35128 9734 35184
rect 7838 29588 7840 29608
rect 7840 29588 7892 29608
rect 7892 29588 7894 29608
rect 7838 29552 7894 29588
rect 7746 27276 7748 27296
rect 7748 27276 7800 27296
rect 7800 27276 7802 27296
rect 7746 27240 7802 27276
rect 7654 27004 7656 27024
rect 7656 27004 7708 27024
rect 7708 27004 7710 27024
rect 7654 26968 7710 27004
rect 7470 26152 7526 26208
rect 7378 25608 7434 25664
rect 7010 24928 7066 24984
rect 6918 23976 6974 24032
rect 5998 23296 6054 23352
rect 5814 23160 5870 23216
rect 5354 22072 5410 22128
rect 5354 21800 5410 21856
rect 6366 23024 6422 23080
rect 6090 22480 6146 22536
rect 5906 22344 5962 22400
rect 5906 22108 5908 22128
rect 5908 22108 5960 22128
rect 5960 22108 5962 22128
rect 5906 22072 5962 22108
rect 6274 22344 6330 22400
rect 5538 21664 5594 21720
rect 5262 21120 5318 21176
rect 5170 20440 5226 20496
rect 5262 20032 5318 20088
rect 4986 19896 5042 19952
rect 5262 19896 5318 19952
rect 4250 19760 4306 19816
rect 4618 19760 4674 19816
rect 5262 19796 5264 19816
rect 5264 19796 5316 19816
rect 5316 19796 5318 19816
rect 5262 19760 5318 19796
rect 3514 18808 3570 18864
rect 3606 18420 3662 18456
rect 3606 18400 3608 18420
rect 3608 18400 3660 18420
rect 3660 18400 3662 18420
rect 4066 19624 4122 19680
rect 4526 19488 4582 19544
rect 5170 19488 5226 19544
rect 4986 19372 5042 19408
rect 4986 19352 4988 19372
rect 4988 19352 5040 19372
rect 5040 19352 5042 19372
rect 5630 21528 5686 21584
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4066 17720 4122 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 5814 21120 5870 21176
rect 6734 23568 6790 23624
rect 6550 22480 6606 22536
rect 6550 21800 6606 21856
rect 6550 21392 6606 21448
rect 6274 21256 6330 21312
rect 6366 21120 6422 21176
rect 6182 20712 6238 20768
rect 6550 20576 6606 20632
rect 5906 19896 5962 19952
rect 6182 19896 6238 19952
rect 6366 19796 6368 19816
rect 6368 19796 6420 19816
rect 6420 19796 6422 19816
rect 6366 19760 6422 19796
rect 6090 19080 6146 19136
rect 7194 25064 7250 25120
rect 7102 23840 7158 23896
rect 7010 23296 7066 23352
rect 7562 26016 7618 26072
rect 6918 23024 6974 23080
rect 6918 22924 6920 22944
rect 6920 22924 6972 22944
rect 6972 22924 6974 22944
rect 6918 22888 6974 22924
rect 8298 27668 8354 27704
rect 8298 27648 8300 27668
rect 8300 27648 8352 27668
rect 8352 27648 8354 27668
rect 8298 27376 8354 27432
rect 9770 33088 9826 33144
rect 10966 36100 11022 36136
rect 10966 36080 10968 36100
rect 10968 36080 11020 36100
rect 11020 36080 11022 36100
rect 10966 34720 11022 34776
rect 10506 33924 10562 33960
rect 10506 33904 10508 33924
rect 10508 33904 10560 33924
rect 10560 33904 10562 33924
rect 10322 32836 10378 32872
rect 10322 32816 10324 32836
rect 10324 32816 10376 32836
rect 10376 32816 10378 32836
rect 8942 31340 8998 31376
rect 8942 31320 8944 31340
rect 8944 31320 8996 31340
rect 8996 31320 8998 31340
rect 8758 30232 8814 30288
rect 8206 27240 8262 27296
rect 8298 27124 8354 27160
rect 8298 27104 8300 27124
rect 8300 27104 8352 27124
rect 8352 27104 8354 27124
rect 7562 24792 7618 24848
rect 7654 24656 7710 24712
rect 7378 23296 7434 23352
rect 6918 22072 6974 22128
rect 7286 21936 7342 21992
rect 7010 21528 7066 21584
rect 6918 21140 6974 21176
rect 6918 21120 6920 21140
rect 6920 21120 6972 21140
rect 6972 21120 6974 21140
rect 7378 21256 7434 21312
rect 7562 22480 7618 22536
rect 7562 22208 7618 22264
rect 7194 20984 7250 21040
rect 6826 20748 6828 20768
rect 6828 20748 6880 20768
rect 6880 20748 6882 20768
rect 6826 20712 6882 20748
rect 6826 20576 6882 20632
rect 6918 20440 6974 20496
rect 5722 17604 5778 17640
rect 5722 17584 5724 17604
rect 5724 17584 5776 17604
rect 5776 17584 5778 17604
rect 4066 16088 4122 16144
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5998 17040 6054 17096
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1214 13096 1270 13152
rect 5906 16904 5962 16960
rect 6274 18692 6330 18728
rect 6274 18672 6276 18692
rect 6276 18672 6328 18692
rect 6328 18672 6330 18692
rect 6918 19080 6974 19136
rect 7378 20848 7434 20904
rect 7194 20712 7250 20768
rect 7562 20712 7618 20768
rect 7378 20440 7434 20496
rect 7286 19488 7342 19544
rect 7470 19796 7472 19816
rect 7472 19796 7524 19816
rect 7524 19796 7526 19816
rect 7470 19760 7526 19796
rect 7930 24148 7932 24168
rect 7932 24148 7984 24168
rect 7984 24148 7986 24168
rect 7930 24112 7986 24148
rect 8298 26016 8354 26072
rect 9126 29144 9182 29200
rect 9034 27784 9090 27840
rect 8482 25916 8484 25936
rect 8484 25916 8536 25936
rect 8536 25916 8538 25936
rect 8482 25880 8538 25916
rect 8206 25472 8262 25528
rect 8114 24148 8116 24168
rect 8116 24148 8168 24168
rect 8168 24148 8170 24168
rect 8114 24112 8170 24148
rect 8206 23976 8262 24032
rect 9126 26832 9182 26888
rect 11794 35128 11850 35184
rect 11794 34584 11850 34640
rect 12070 34720 12126 34776
rect 12162 34604 12218 34640
rect 12162 34584 12164 34604
rect 12164 34584 12216 34604
rect 12216 34584 12218 34604
rect 11702 34060 11758 34096
rect 11702 34040 11704 34060
rect 11704 34040 11756 34060
rect 11756 34040 11758 34060
rect 11334 33496 11390 33552
rect 10966 33224 11022 33280
rect 9678 31728 9734 31784
rect 9494 29164 9550 29200
rect 9494 29144 9496 29164
rect 9496 29144 9548 29164
rect 9548 29144 9550 29164
rect 10598 31592 10654 31648
rect 10046 30368 10102 30424
rect 9862 29280 9918 29336
rect 9586 27648 9642 27704
rect 8390 24520 8446 24576
rect 7930 21664 7986 21720
rect 7930 21528 7986 21584
rect 7654 20032 7710 20088
rect 7746 19896 7802 19952
rect 7746 19760 7802 19816
rect 7378 19352 7434 19408
rect 7194 19080 7250 19136
rect 6550 18264 6606 18320
rect 6458 16108 6514 16144
rect 6458 16088 6460 16108
rect 6460 16088 6512 16108
rect 6512 16088 6514 16108
rect 7286 18284 7342 18320
rect 7286 18264 7288 18284
rect 7288 18264 7340 18284
rect 7340 18264 7342 18284
rect 7102 17992 7158 18048
rect 7010 17584 7066 17640
rect 7194 17856 7250 17912
rect 7286 17448 7342 17504
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 8390 22344 8446 22400
rect 8298 22208 8354 22264
rect 8390 21800 8446 21856
rect 8114 21120 8170 21176
rect 8022 20868 8078 20904
rect 8022 20848 8024 20868
rect 8024 20848 8076 20868
rect 8076 20848 8078 20868
rect 8206 20848 8262 20904
rect 8298 20576 8354 20632
rect 7930 20440 7986 20496
rect 8390 20476 8392 20496
rect 8392 20476 8444 20496
rect 8444 20476 8446 20496
rect 8390 20440 8446 20476
rect 8574 21664 8630 21720
rect 8206 20032 8262 20088
rect 8114 19488 8170 19544
rect 7378 16496 7434 16552
rect 7746 18028 7748 18048
rect 7748 18028 7800 18048
rect 7800 18028 7802 18048
rect 7746 17992 7802 18028
rect 8482 20304 8538 20360
rect 8390 18964 8446 19000
rect 8390 18944 8392 18964
rect 8392 18944 8444 18964
rect 8444 18944 8446 18964
rect 7654 16632 7710 16688
rect 8206 17856 8262 17912
rect 8390 18572 8392 18592
rect 8392 18572 8444 18592
rect 8444 18572 8446 18592
rect 8390 18536 8446 18572
rect 8390 17992 8446 18048
rect 9034 24812 9090 24848
rect 9034 24792 9036 24812
rect 9036 24792 9088 24812
rect 9088 24792 9090 24812
rect 9034 23976 9090 24032
rect 9770 25744 9826 25800
rect 9586 25336 9642 25392
rect 9034 22636 9090 22672
rect 9034 22616 9036 22636
rect 9036 22616 9088 22636
rect 9088 22616 9090 22636
rect 9494 24384 9550 24440
rect 9862 25064 9918 25120
rect 9770 23976 9826 24032
rect 10230 29688 10286 29744
rect 10874 29164 10930 29200
rect 10874 29144 10876 29164
rect 10876 29144 10928 29164
rect 10928 29144 10930 29164
rect 10414 27396 10470 27432
rect 10414 27376 10416 27396
rect 10416 27376 10468 27396
rect 10468 27376 10470 27396
rect 10782 27104 10838 27160
rect 9586 22888 9642 22944
rect 9494 22480 9550 22536
rect 9402 22072 9458 22128
rect 8942 21664 8998 21720
rect 8942 21528 8998 21584
rect 8758 19760 8814 19816
rect 7838 15136 7894 15192
rect 1214 12008 1270 12064
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1858 10920 1914 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1214 9832 1270 9888
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3146 8880 3202 8936
rect 1214 8744 1270 8800
rect 1214 7656 1270 7712
rect 1214 6568 1270 6624
rect 1858 5480 1914 5536
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 9310 21800 9366 21856
rect 9402 21392 9458 21448
rect 9402 20984 9458 21040
rect 9402 20460 9458 20496
rect 9402 20440 9404 20460
rect 9404 20440 9456 20460
rect 9456 20440 9458 20460
rect 9310 20168 9366 20224
rect 9770 21664 9826 21720
rect 9770 20460 9826 20496
rect 9770 20440 9772 20460
rect 9772 20440 9824 20460
rect 9824 20440 9826 20460
rect 9586 19624 9642 19680
rect 9862 18808 9918 18864
rect 9126 18536 9182 18592
rect 10230 24792 10286 24848
rect 10138 22072 10194 22128
rect 10138 21800 10194 21856
rect 10690 24384 10746 24440
rect 10414 22344 10470 22400
rect 11334 30252 11390 30288
rect 11334 30232 11336 30252
rect 11336 30232 11388 30252
rect 11388 30232 11390 30252
rect 11058 29164 11114 29200
rect 11058 29144 11060 29164
rect 11060 29144 11112 29164
rect 11112 29144 11114 29164
rect 11058 27648 11114 27704
rect 11702 33360 11758 33416
rect 12438 33940 12440 33960
rect 12440 33940 12492 33960
rect 12492 33940 12494 33960
rect 12438 33904 12494 33940
rect 13266 35572 13268 35592
rect 13268 35572 13320 35592
rect 13320 35572 13322 35592
rect 13266 35536 13322 35572
rect 13266 34060 13322 34096
rect 13266 34040 13268 34060
rect 13268 34040 13320 34060
rect 13320 34040 13322 34060
rect 12254 33516 12310 33552
rect 12254 33496 12256 33516
rect 12256 33496 12308 33516
rect 12308 33496 12310 33516
rect 12254 31592 12310 31648
rect 12714 33360 12770 33416
rect 13174 33652 13230 33688
rect 13174 33632 13176 33652
rect 13176 33632 13228 33652
rect 13228 33632 13230 33652
rect 13266 33360 13322 33416
rect 12990 32136 13046 32192
rect 11886 29844 11942 29880
rect 11886 29824 11888 29844
rect 11888 29824 11940 29844
rect 11940 29824 11942 29844
rect 11886 29688 11942 29744
rect 11978 29416 12034 29472
rect 12714 29452 12716 29472
rect 12716 29452 12768 29472
rect 12768 29452 12770 29472
rect 12714 29416 12770 29452
rect 11242 26968 11298 27024
rect 11058 26016 11114 26072
rect 11150 25880 11206 25936
rect 11150 25236 11152 25256
rect 11152 25236 11204 25256
rect 11204 25236 11206 25256
rect 11150 25200 11206 25236
rect 10874 25064 10930 25120
rect 11426 26016 11482 26072
rect 11978 26988 12034 27024
rect 11978 26968 11980 26988
rect 11980 26968 12032 26988
rect 12032 26968 12034 26988
rect 10598 23160 10654 23216
rect 10598 22888 10654 22944
rect 10506 21936 10562 21992
rect 10046 20884 10048 20904
rect 10048 20884 10100 20904
rect 10100 20884 10102 20904
rect 10046 20848 10102 20884
rect 10322 20440 10378 20496
rect 9586 18128 9642 18184
rect 9126 18028 9128 18048
rect 9128 18028 9180 18048
rect 9180 18028 9182 18048
rect 9126 17992 9182 18028
rect 10414 20032 10470 20088
rect 11058 23840 11114 23896
rect 11518 25336 11574 25392
rect 11058 23060 11060 23080
rect 11060 23060 11112 23080
rect 11112 23060 11114 23080
rect 11058 23024 11114 23060
rect 10782 22636 10838 22672
rect 10782 22616 10784 22636
rect 10784 22616 10836 22636
rect 10836 22616 10838 22636
rect 11242 22752 11298 22808
rect 10874 22480 10930 22536
rect 10782 22344 10838 22400
rect 11058 21392 11114 21448
rect 11426 22344 11482 22400
rect 11702 24384 11758 24440
rect 11610 23060 11612 23080
rect 11612 23060 11664 23080
rect 11664 23060 11666 23080
rect 11610 23024 11666 23060
rect 11610 22516 11612 22536
rect 11612 22516 11664 22536
rect 11664 22516 11666 22536
rect 11610 22480 11666 22516
rect 11426 21800 11482 21856
rect 11518 21528 11574 21584
rect 11150 21120 11206 21176
rect 10782 20712 10838 20768
rect 11058 20748 11060 20768
rect 11060 20748 11112 20768
rect 11112 20748 11114 20768
rect 10690 20168 10746 20224
rect 11058 20712 11114 20748
rect 10874 20304 10930 20360
rect 10874 20032 10930 20088
rect 10506 18692 10562 18728
rect 10506 18672 10508 18692
rect 10508 18672 10560 18692
rect 10560 18672 10562 18692
rect 10874 18944 10930 19000
rect 10782 18808 10838 18864
rect 11150 20204 11152 20224
rect 11152 20204 11204 20224
rect 11204 20204 11206 20224
rect 11150 20168 11206 20204
rect 11334 21256 11390 21312
rect 11334 19896 11390 19952
rect 11058 19080 11114 19136
rect 10966 17856 11022 17912
rect 11886 25608 11942 25664
rect 12990 29824 13046 29880
rect 13174 29588 13176 29608
rect 13176 29588 13228 29608
rect 13228 29588 13230 29608
rect 13174 29552 13230 29588
rect 12622 27412 12624 27432
rect 12624 27412 12676 27432
rect 12676 27412 12678 27432
rect 12622 27376 12678 27412
rect 11886 24928 11942 24984
rect 12070 23568 12126 23624
rect 12254 25064 12310 25120
rect 12254 23840 12310 23896
rect 13082 29144 13138 29200
rect 13174 29008 13230 29064
rect 14278 36760 14334 36816
rect 13634 33224 13690 33280
rect 13634 33108 13690 33144
rect 13634 33088 13636 33108
rect 13636 33088 13688 33108
rect 13688 33088 13690 33108
rect 13634 32564 13690 32600
rect 13634 32544 13636 32564
rect 13636 32544 13688 32564
rect 13688 32544 13690 32564
rect 13542 32272 13598 32328
rect 13634 31320 13690 31376
rect 13542 29688 13598 29744
rect 13726 29552 13782 29608
rect 13082 27648 13138 27704
rect 12990 25336 13046 25392
rect 12714 24268 12770 24304
rect 12714 24248 12716 24268
rect 12716 24248 12768 24268
rect 12768 24248 12770 24268
rect 12622 23724 12678 23760
rect 13266 25764 13322 25800
rect 13266 25744 13268 25764
rect 13268 25744 13320 25764
rect 13320 25744 13322 25764
rect 12622 23704 12624 23724
rect 12624 23704 12676 23724
rect 12676 23704 12678 23724
rect 11978 22616 12034 22672
rect 11886 22208 11942 22264
rect 12530 22480 12586 22536
rect 11886 20168 11942 20224
rect 12898 21428 12900 21448
rect 12900 21428 12952 21448
rect 12952 21428 12954 21448
rect 12898 21392 12954 21428
rect 12070 20984 12126 21040
rect 12162 20440 12218 20496
rect 12070 19624 12126 19680
rect 11978 19372 12034 19408
rect 11978 19352 11980 19372
rect 11980 19352 12032 19372
rect 12032 19352 12034 19372
rect 12438 20984 12494 21040
rect 12346 20032 12402 20088
rect 13266 24384 13322 24440
rect 14922 37712 14978 37768
rect 14922 36760 14978 36816
rect 14738 36080 14794 36136
rect 15014 34720 15070 34776
rect 14922 34176 14978 34232
rect 14002 32428 14058 32464
rect 14002 32408 14004 32428
rect 14004 32408 14056 32428
rect 14056 32408 14058 32428
rect 13542 27512 13598 27568
rect 15842 37032 15898 37088
rect 14554 32000 14610 32056
rect 14370 31864 14426 31920
rect 14278 29960 14334 30016
rect 14462 30368 14518 30424
rect 14462 29708 14518 29744
rect 14462 29688 14464 29708
rect 14464 29688 14516 29708
rect 14516 29688 14518 29708
rect 14830 32272 14886 32328
rect 15382 34448 15438 34504
rect 15658 33360 15714 33416
rect 15382 33224 15438 33280
rect 15382 32544 15438 32600
rect 14646 30504 14702 30560
rect 13818 27648 13874 27704
rect 13726 24928 13782 24984
rect 13726 24812 13782 24848
rect 13726 24792 13728 24812
rect 13728 24792 13780 24812
rect 13780 24792 13782 24812
rect 13358 22888 13414 22944
rect 14186 28056 14242 28112
rect 14002 27240 14058 27296
rect 14370 27820 14372 27840
rect 14372 27820 14424 27840
rect 14424 27820 14426 27840
rect 14370 27784 14426 27820
rect 15106 28872 15162 28928
rect 13910 24248 13966 24304
rect 13634 23296 13690 23352
rect 14094 24404 14150 24440
rect 14094 24384 14096 24404
rect 14096 24384 14148 24404
rect 14148 24384 14150 24404
rect 13634 21664 13690 21720
rect 12898 20748 12900 20768
rect 12900 20748 12952 20768
rect 12952 20748 12954 20768
rect 12898 20712 12954 20748
rect 13082 20440 13138 20496
rect 13174 20304 13230 20360
rect 13358 21120 13414 21176
rect 12990 20168 13046 20224
rect 12622 18672 12678 18728
rect 11702 16632 11758 16688
rect 12070 16632 12126 16688
rect 12622 17720 12678 17776
rect 12162 16496 12218 16552
rect 13174 17856 13230 17912
rect 13542 19760 13598 19816
rect 13450 18148 13506 18184
rect 13450 18128 13452 18148
rect 13452 18128 13504 18148
rect 13504 18128 13506 18148
rect 13910 21936 13966 21992
rect 14278 24520 14334 24576
rect 13726 18944 13782 19000
rect 13818 18264 13874 18320
rect 13634 17604 13690 17640
rect 13634 17584 13636 17604
rect 13636 17584 13688 17604
rect 13688 17584 13690 17604
rect 13450 17332 13506 17368
rect 13450 17312 13452 17332
rect 13452 17312 13504 17332
rect 13504 17312 13506 17332
rect 13634 17176 13690 17232
rect 13542 17040 13598 17096
rect 13174 15564 13230 15600
rect 13174 15544 13176 15564
rect 13176 15544 13228 15564
rect 13228 15544 13230 15564
rect 14002 21292 14004 21312
rect 14004 21292 14056 21312
rect 14056 21292 14058 21312
rect 14002 21256 14058 21292
rect 14738 25608 14794 25664
rect 14646 24928 14702 24984
rect 15014 27240 15070 27296
rect 15474 32136 15530 32192
rect 16762 34620 16764 34640
rect 16764 34620 16816 34640
rect 16816 34620 16818 34640
rect 16762 34584 16818 34620
rect 16026 32544 16082 32600
rect 15842 31728 15898 31784
rect 15474 30932 15530 30968
rect 15474 30912 15476 30932
rect 15476 30912 15528 30932
rect 15528 30912 15530 30932
rect 15474 30252 15530 30288
rect 15474 30232 15476 30252
rect 15476 30232 15528 30252
rect 15528 30232 15530 30252
rect 15474 29724 15476 29744
rect 15476 29724 15528 29744
rect 15528 29724 15530 29744
rect 15474 29688 15530 29724
rect 15106 27104 15162 27160
rect 15106 24520 15162 24576
rect 14922 23160 14978 23216
rect 14094 19896 14150 19952
rect 14186 19488 14242 19544
rect 14002 17196 14058 17232
rect 14002 17176 14004 17196
rect 14004 17176 14056 17196
rect 14056 17176 14058 17196
rect 14278 18844 14280 18864
rect 14280 18844 14332 18864
rect 14332 18844 14334 18864
rect 14278 18808 14334 18844
rect 14278 18264 14334 18320
rect 14462 20032 14518 20088
rect 15934 30252 15990 30288
rect 15934 30232 15936 30252
rect 15936 30232 15988 30252
rect 15988 30232 15990 30252
rect 17222 37732 17278 37768
rect 17222 37712 17224 37732
rect 17224 37712 17276 37732
rect 17276 37712 17278 37732
rect 17222 37204 17224 37224
rect 17224 37204 17276 37224
rect 17276 37204 17278 37224
rect 17222 37168 17278 37204
rect 17038 37032 17094 37088
rect 17130 35536 17186 35592
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 17498 36100 17554 36136
rect 17498 36080 17500 36100
rect 17500 36080 17552 36100
rect 17552 36080 17554 36100
rect 16762 32444 16764 32464
rect 16764 32444 16816 32464
rect 16816 32444 16818 32464
rect 16762 32408 16818 32444
rect 16118 29688 16174 29744
rect 16302 29416 16358 29472
rect 16210 27104 16266 27160
rect 16026 26968 16082 27024
rect 15658 26152 15714 26208
rect 15382 25100 15384 25120
rect 15384 25100 15436 25120
rect 15436 25100 15438 25120
rect 15382 25064 15438 25100
rect 16026 26424 16082 26480
rect 15014 22344 15070 22400
rect 15014 21972 15016 21992
rect 15016 21972 15068 21992
rect 15068 21972 15070 21992
rect 15014 21936 15070 21972
rect 14922 21664 14978 21720
rect 15106 21392 15162 21448
rect 14186 16632 14242 16688
rect 13818 16496 13874 16552
rect 14554 18420 14610 18456
rect 14554 18400 14556 18420
rect 14556 18400 14608 18420
rect 14608 18400 14610 18420
rect 14830 21256 14886 21312
rect 14830 20304 14886 20360
rect 15842 25608 15898 25664
rect 15934 25472 15990 25528
rect 16118 26016 16174 26072
rect 15750 24112 15806 24168
rect 14646 18148 14702 18184
rect 14646 18128 14648 18148
rect 14648 18128 14700 18148
rect 14700 18128 14702 18148
rect 15382 19252 15384 19272
rect 15384 19252 15436 19272
rect 15436 19252 15438 19272
rect 15382 19216 15438 19252
rect 15106 19080 15162 19136
rect 15290 18284 15346 18320
rect 15290 18264 15292 18284
rect 15292 18264 15344 18284
rect 15344 18264 15346 18284
rect 15198 18128 15254 18184
rect 14830 17720 14886 17776
rect 15290 17756 15292 17776
rect 15292 17756 15344 17776
rect 15344 17756 15346 17776
rect 15290 17720 15346 17756
rect 15106 17176 15162 17232
rect 15014 16904 15070 16960
rect 15382 16532 15384 16552
rect 15384 16532 15436 16552
rect 15436 16532 15438 16552
rect 15382 16496 15438 16532
rect 15658 21120 15714 21176
rect 15750 20848 15806 20904
rect 16486 30132 16488 30152
rect 16488 30132 16540 30152
rect 16540 30132 16542 30152
rect 16486 30096 16542 30132
rect 16486 28076 16542 28112
rect 16486 28056 16488 28076
rect 16488 28056 16540 28076
rect 16540 28056 16542 28076
rect 16394 26560 16450 26616
rect 16762 27956 16764 27976
rect 16764 27956 16816 27976
rect 16816 27956 16818 27976
rect 16762 27920 16818 27956
rect 16762 27512 16818 27568
rect 16762 27240 16818 27296
rect 16394 25780 16396 25800
rect 16396 25780 16448 25800
rect 16448 25780 16450 25800
rect 16394 25744 16450 25780
rect 15934 22480 15990 22536
rect 15658 19780 15714 19816
rect 15658 19760 15660 19780
rect 15660 19760 15712 19780
rect 15712 19760 15714 19780
rect 16302 23296 16358 23352
rect 17406 30912 17462 30968
rect 18050 31900 18052 31920
rect 18052 31900 18104 31920
rect 18104 31900 18106 31920
rect 18050 31864 18106 31900
rect 17682 31184 17738 31240
rect 17314 30676 17316 30696
rect 17316 30676 17368 30696
rect 17368 30676 17370 30696
rect 17314 30640 17370 30676
rect 17038 29280 17094 29336
rect 17038 27240 17094 27296
rect 17958 30368 18014 30424
rect 17314 27920 17370 27976
rect 17958 30252 18014 30288
rect 17958 30232 17960 30252
rect 17960 30232 18012 30252
rect 18012 30232 18014 30252
rect 17866 29824 17922 29880
rect 17774 27512 17830 27568
rect 17406 27276 17408 27296
rect 17408 27276 17460 27296
rect 17460 27276 17462 27296
rect 17406 27240 17462 27276
rect 17406 26832 17462 26888
rect 17314 26308 17370 26344
rect 17314 26288 17316 26308
rect 17316 26288 17368 26308
rect 17368 26288 17370 26308
rect 16670 24928 16726 24984
rect 16854 24248 16910 24304
rect 16486 22072 16542 22128
rect 16578 21548 16634 21584
rect 16578 21528 16580 21548
rect 16580 21528 16632 21548
rect 16632 21528 16634 21548
rect 16486 21256 16542 21312
rect 16762 21392 16818 21448
rect 16578 20848 16634 20904
rect 16118 18964 16174 19000
rect 16118 18944 16120 18964
rect 16120 18944 16172 18964
rect 16172 18944 16174 18964
rect 16118 18808 16174 18864
rect 16026 18400 16082 18456
rect 15750 17040 15806 17096
rect 16394 19896 16450 19952
rect 16578 20748 16580 20768
rect 16580 20748 16632 20768
rect 16632 20748 16634 20768
rect 16578 20712 16634 20748
rect 16486 18420 16542 18456
rect 16486 18400 16488 18420
rect 16488 18400 16540 18420
rect 16540 18400 16542 18420
rect 17590 27240 17646 27296
rect 18142 29552 18198 29608
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 18510 34584 18566 34640
rect 18510 32680 18566 32736
rect 18694 32000 18750 32056
rect 18602 31048 18658 31104
rect 18510 30912 18566 30968
rect 19246 37188 19302 37224
rect 19246 37168 19248 37188
rect 19248 37168 19300 37188
rect 19300 37168 19302 37188
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 21178 38548 21234 38584
rect 21178 38528 21180 38548
rect 21180 38528 21232 38548
rect 21232 38528 21234 38548
rect 20718 38412 20774 38448
rect 20718 38392 20720 38412
rect 20720 38392 20772 38412
rect 20772 38392 20774 38412
rect 21270 38120 21326 38176
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19982 34856 20038 34912
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 18878 32816 18934 32872
rect 18326 30504 18382 30560
rect 18602 29416 18658 29472
rect 18142 28192 18198 28248
rect 17222 24928 17278 24984
rect 17222 24284 17224 24304
rect 17224 24284 17276 24304
rect 17276 24284 17278 24304
rect 17222 24248 17278 24284
rect 17314 23704 17370 23760
rect 17038 23160 17094 23216
rect 17222 23160 17278 23216
rect 16946 22072 17002 22128
rect 17314 23024 17370 23080
rect 17314 22924 17316 22944
rect 17316 22924 17368 22944
rect 17368 22924 17370 22944
rect 17314 22888 17370 22924
rect 17222 22636 17278 22672
rect 17222 22616 17224 22636
rect 17224 22616 17276 22636
rect 17276 22616 17278 22636
rect 16762 18808 16818 18864
rect 17130 21412 17186 21448
rect 17130 21392 17132 21412
rect 17132 21392 17184 21412
rect 17184 21392 17186 21412
rect 17498 25200 17554 25256
rect 18050 26288 18106 26344
rect 18234 27784 18290 27840
rect 18602 28636 18604 28656
rect 18604 28636 18656 28656
rect 18656 28636 18658 28656
rect 18602 28600 18658 28636
rect 18602 27784 18658 27840
rect 18326 26560 18382 26616
rect 18142 25744 18198 25800
rect 18510 25336 18566 25392
rect 17866 23976 17922 24032
rect 17682 23432 17738 23488
rect 17774 23160 17830 23216
rect 17406 22480 17462 22536
rect 17314 20576 17370 20632
rect 16394 18128 16450 18184
rect 16302 17856 16358 17912
rect 16210 17584 16266 17640
rect 16578 16904 16634 16960
rect 16854 17620 16856 17640
rect 16856 17620 16908 17640
rect 16908 17620 16910 17640
rect 16854 17584 16910 17620
rect 17314 19216 17370 19272
rect 17590 22380 17592 22400
rect 17592 22380 17644 22400
rect 17644 22380 17646 22400
rect 17590 22344 17646 22380
rect 17498 21800 17554 21856
rect 17498 21392 17554 21448
rect 18050 23160 18106 23216
rect 17866 21800 17922 21856
rect 17590 19216 17646 19272
rect 17590 18264 17646 18320
rect 18050 21004 18106 21040
rect 18050 20984 18052 21004
rect 18052 20984 18104 21004
rect 18104 20984 18106 21004
rect 18602 24148 18604 24168
rect 18604 24148 18656 24168
rect 18656 24148 18658 24168
rect 18602 24112 18658 24148
rect 18510 23296 18566 23352
rect 18326 23044 18382 23080
rect 18326 23024 18328 23044
rect 18328 23024 18380 23044
rect 18380 23024 18382 23044
rect 18326 22208 18382 22264
rect 18050 19216 18106 19272
rect 18510 22208 18566 22264
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19154 31340 19210 31376
rect 19154 31320 19156 31340
rect 19156 31320 19208 31340
rect 19208 31320 19210 31340
rect 19154 31204 19210 31240
rect 19154 31184 19156 31204
rect 19156 31184 19208 31204
rect 19208 31184 19210 31204
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19522 30776 19578 30832
rect 19154 30232 19210 30288
rect 19154 29960 19210 30016
rect 20166 31320 20222 31376
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 18878 26968 18934 27024
rect 18786 25472 18842 25528
rect 19338 28464 19394 28520
rect 20166 30504 20222 30560
rect 19890 28636 19892 28656
rect 19892 28636 19944 28656
rect 19944 28636 19946 28656
rect 20166 29416 20222 29472
rect 19890 28600 19946 28636
rect 19798 28464 19854 28520
rect 19154 27784 19210 27840
rect 19062 27240 19118 27296
rect 19246 26696 19302 26752
rect 19062 26152 19118 26208
rect 18970 24656 19026 24712
rect 19062 24384 19118 24440
rect 19062 23976 19118 24032
rect 18786 22888 18842 22944
rect 18878 22752 18934 22808
rect 18510 21664 18566 21720
rect 18970 22344 19026 22400
rect 18970 22208 19026 22264
rect 18418 20596 18474 20632
rect 18418 20576 18420 20596
rect 18420 20576 18472 20596
rect 18472 20576 18474 20596
rect 18326 19896 18382 19952
rect 18418 18944 18474 19000
rect 18418 18536 18474 18592
rect 17406 17992 17462 18048
rect 17314 17312 17370 17368
rect 17590 17756 17592 17776
rect 17592 17756 17644 17776
rect 17644 17756 17646 17776
rect 17590 17720 17646 17756
rect 18694 20848 18750 20904
rect 18602 19624 18658 19680
rect 18970 21800 19026 21856
rect 18970 21664 19026 21720
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19798 27376 19854 27432
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 20166 28600 20222 28656
rect 19614 26696 19670 26752
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19798 25336 19854 25392
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19338 23976 19394 24032
rect 19706 24656 19762 24712
rect 20166 25064 20222 25120
rect 20074 24928 20130 24984
rect 21638 38392 21694 38448
rect 21914 38528 21970 38584
rect 21270 34604 21326 34640
rect 21270 34584 21272 34604
rect 21272 34584 21324 34604
rect 21324 34584 21326 34604
rect 21178 33768 21234 33824
rect 20718 30796 20774 30832
rect 20718 30776 20720 30796
rect 20720 30776 20772 30796
rect 20772 30776 20774 30796
rect 20534 30540 20536 30560
rect 20536 30540 20588 30560
rect 20588 30540 20590 30560
rect 20534 30504 20590 30540
rect 23110 36624 23166 36680
rect 21546 33224 21602 33280
rect 21362 32952 21418 33008
rect 20442 30268 20444 30288
rect 20444 30268 20496 30288
rect 20496 30268 20498 30288
rect 20442 30232 20498 30268
rect 20810 30232 20866 30288
rect 20350 29552 20406 29608
rect 21362 31184 21418 31240
rect 21270 30368 21326 30424
rect 21362 30096 21418 30152
rect 21546 30096 21602 30152
rect 22374 34584 22430 34640
rect 23018 34584 23074 34640
rect 21822 30504 21878 30560
rect 21730 29688 21786 29744
rect 21178 29416 21234 29472
rect 21454 29416 21510 29472
rect 21454 29280 21510 29336
rect 22374 30912 22430 30968
rect 22650 30640 22706 30696
rect 22098 29280 22154 29336
rect 20442 29008 20498 29064
rect 20810 28056 20866 28112
rect 20534 26424 20590 26480
rect 20718 25900 20774 25936
rect 20718 25880 20720 25900
rect 20720 25880 20772 25900
rect 20772 25880 20774 25900
rect 21270 27820 21272 27840
rect 21272 27820 21324 27840
rect 21324 27820 21326 27840
rect 21270 27784 21326 27820
rect 20902 25880 20958 25936
rect 20902 25608 20958 25664
rect 20626 25336 20682 25392
rect 20350 25064 20406 25120
rect 20442 24928 20498 24984
rect 19982 23976 20038 24032
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19430 23840 19486 23896
rect 19890 23316 19946 23352
rect 19890 23296 19892 23316
rect 19892 23296 19944 23316
rect 19944 23296 19946 23316
rect 21546 26016 21602 26072
rect 22190 27396 22246 27432
rect 22190 27376 22192 27396
rect 22192 27376 22244 27396
rect 22244 27376 22246 27396
rect 22190 27104 22246 27160
rect 22558 29144 22614 29200
rect 22650 28908 22652 28928
rect 22652 28908 22704 28928
rect 22704 28908 22706 28928
rect 22650 28872 22706 28908
rect 22098 26988 22154 27024
rect 22098 26968 22100 26988
rect 22100 26968 22152 26988
rect 22152 26968 22154 26988
rect 22650 26696 22706 26752
rect 22466 26152 22522 26208
rect 21546 24948 21602 24984
rect 21546 24928 21548 24948
rect 21548 24928 21600 24948
rect 21600 24928 21602 24948
rect 20902 24676 20958 24712
rect 20902 24656 20904 24676
rect 20904 24656 20956 24676
rect 20956 24656 20958 24676
rect 21270 24656 21326 24712
rect 21178 24384 21234 24440
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20258 22888 20314 22944
rect 19614 22652 19616 22672
rect 19616 22652 19668 22672
rect 19668 22652 19670 22672
rect 19614 22616 19670 22652
rect 19798 22616 19854 22672
rect 19246 22480 19302 22536
rect 19154 21800 19210 21856
rect 20626 22752 20682 22808
rect 21086 23976 21142 24032
rect 21178 23840 21234 23896
rect 22466 25236 22468 25256
rect 22468 25236 22520 25256
rect 22520 25236 22522 25256
rect 22466 25200 22522 25236
rect 21546 24148 21548 24168
rect 21548 24148 21600 24168
rect 21600 24148 21602 24168
rect 21546 24112 21602 24148
rect 20074 22344 20130 22400
rect 20534 22380 20536 22400
rect 20536 22380 20588 22400
rect 20588 22380 20590 22400
rect 20534 22344 20590 22380
rect 20350 22208 20406 22264
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 18786 20440 18842 20496
rect 18970 19760 19026 19816
rect 18786 18420 18842 18456
rect 18786 18400 18788 18420
rect 18788 18400 18840 18420
rect 18840 18400 18842 18420
rect 18418 17584 18474 17640
rect 19246 21120 19302 21176
rect 20166 22072 20222 22128
rect 20534 22072 20590 22128
rect 20442 21936 20498 21992
rect 20350 21800 20406 21856
rect 20258 21664 20314 21720
rect 19798 21292 19800 21312
rect 19800 21292 19852 21312
rect 19852 21292 19854 21312
rect 19798 21256 19854 21292
rect 19982 20984 20038 21040
rect 19890 20884 19892 20904
rect 19892 20884 19944 20904
rect 19944 20884 19946 20904
rect 19890 20848 19946 20884
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19430 20576 19486 20632
rect 19246 20168 19302 20224
rect 20258 20984 20314 21040
rect 20166 20712 20222 20768
rect 19982 20304 20038 20360
rect 19706 19760 19762 19816
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 19388 19892 19408
rect 19892 19388 19944 19408
rect 19944 19388 19946 19408
rect 19890 19352 19946 19388
rect 19706 18808 19762 18864
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18510 16496 18566 16552
rect 15014 15580 15016 15600
rect 15016 15580 15068 15600
rect 15068 15580 15070 15600
rect 15014 15544 15070 15580
rect 19522 17856 19578 17912
rect 20350 20576 20406 20632
rect 20350 19216 20406 19272
rect 21178 22092 21234 22128
rect 21178 22072 21180 22092
rect 21180 22072 21232 22092
rect 21232 22072 21234 22092
rect 21086 21548 21142 21584
rect 21086 21528 21088 21548
rect 21088 21528 21140 21548
rect 21140 21528 21142 21548
rect 20166 17584 20222 17640
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19890 17196 19946 17232
rect 19890 17176 19892 17196
rect 19892 17176 19944 17196
rect 19944 17176 19946 17196
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20810 20576 20866 20632
rect 20810 18944 20866 19000
rect 20534 17856 20590 17912
rect 21086 20204 21088 20224
rect 21088 20204 21140 20224
rect 21140 20204 21142 20224
rect 21086 20168 21142 20204
rect 21638 22616 21694 22672
rect 21546 22344 21602 22400
rect 21914 24812 21970 24848
rect 21914 24792 21916 24812
rect 21916 24792 21968 24812
rect 21968 24792 21970 24812
rect 22006 24384 22062 24440
rect 21914 23840 21970 23896
rect 22006 23704 22062 23760
rect 21914 23316 21970 23352
rect 21914 23296 21916 23316
rect 21916 23296 21968 23316
rect 21968 23296 21970 23316
rect 21822 22344 21878 22400
rect 21638 21664 21694 21720
rect 21086 17720 21142 17776
rect 20902 17584 20958 17640
rect 21454 21256 21510 21312
rect 21914 21548 21970 21584
rect 21914 21528 21916 21548
rect 21916 21528 21968 21548
rect 21968 21528 21970 21548
rect 22282 23296 22338 23352
rect 22190 22888 22246 22944
rect 21914 21256 21970 21312
rect 21822 20984 21878 21040
rect 21454 19624 21510 19680
rect 21454 19080 21510 19136
rect 21362 18944 21418 19000
rect 21730 18844 21732 18864
rect 21732 18844 21784 18864
rect 21784 18844 21786 18864
rect 21730 18808 21786 18844
rect 21362 18672 21418 18728
rect 22006 19624 22062 19680
rect 21914 19352 21970 19408
rect 22282 18944 22338 19000
rect 22098 18708 22100 18728
rect 22100 18708 22152 18728
rect 22152 18708 22154 18728
rect 22098 18672 22154 18708
rect 21362 17604 21418 17640
rect 21362 17584 21364 17604
rect 21364 17584 21416 17604
rect 21416 17584 21418 17604
rect 21454 17448 21510 17504
rect 21362 17212 21364 17232
rect 21364 17212 21416 17232
rect 21416 17212 21418 17232
rect 21362 17176 21418 17212
rect 22190 18572 22192 18592
rect 22192 18572 22244 18592
rect 22244 18572 22246 18592
rect 22190 18536 22246 18572
rect 21638 17176 21694 17232
rect 21822 17856 21878 17912
rect 22006 18028 22008 18048
rect 22008 18028 22060 18048
rect 22060 18028 22062 18048
rect 22006 17992 22062 18028
rect 22558 23976 22614 24032
rect 23478 35148 23534 35184
rect 23478 35128 23480 35148
rect 23480 35128 23532 35148
rect 23532 35128 23534 35148
rect 23294 33496 23350 33552
rect 22926 30640 22982 30696
rect 22926 30096 22982 30152
rect 23110 30368 23166 30424
rect 23202 29824 23258 29880
rect 23110 29552 23166 29608
rect 22926 29044 22928 29064
rect 22928 29044 22980 29064
rect 22980 29044 22982 29064
rect 22926 29008 22982 29044
rect 22742 24948 22798 24984
rect 22742 24928 22744 24948
rect 22744 24928 22796 24948
rect 22796 24928 22798 24948
rect 25410 38120 25466 38176
rect 24214 37188 24270 37224
rect 24214 37168 24216 37188
rect 24216 37168 24268 37188
rect 24268 37168 24270 37188
rect 23662 32952 23718 33008
rect 24030 33632 24086 33688
rect 23938 32000 23994 32056
rect 24030 31592 24086 31648
rect 23662 31048 23718 31104
rect 23846 30676 23848 30696
rect 23848 30676 23900 30696
rect 23900 30676 23902 30696
rect 23846 30640 23902 30676
rect 23570 29572 23626 29608
rect 23570 29552 23572 29572
rect 23572 29552 23624 29572
rect 23624 29552 23626 29572
rect 23846 29300 23902 29336
rect 23846 29280 23848 29300
rect 23848 29280 23900 29300
rect 23900 29280 23902 29300
rect 23294 27512 23350 27568
rect 23294 27104 23350 27160
rect 23202 26424 23258 26480
rect 23478 27512 23534 27568
rect 23386 26288 23442 26344
rect 22834 24556 22836 24576
rect 22836 24556 22888 24576
rect 22888 24556 22890 24576
rect 22834 24520 22890 24556
rect 22834 23976 22890 24032
rect 23386 25200 23442 25256
rect 23754 26832 23810 26888
rect 24122 29960 24178 30016
rect 24674 33904 24730 33960
rect 25410 35944 25466 36000
rect 26422 36352 26478 36408
rect 25962 35808 26018 35864
rect 25042 34176 25098 34232
rect 24858 33768 24914 33824
rect 24950 33360 25006 33416
rect 25594 34176 25650 34232
rect 25686 34040 25742 34096
rect 25502 33632 25558 33688
rect 24674 32136 24730 32192
rect 24306 31320 24362 31376
rect 24582 31048 24638 31104
rect 24306 30776 24362 30832
rect 24950 31456 25006 31512
rect 25226 32000 25282 32056
rect 24766 31048 24822 31104
rect 24674 30232 24730 30288
rect 24950 30912 25006 30968
rect 25594 32172 25596 32192
rect 25596 32172 25648 32192
rect 25648 32172 25650 32192
rect 25594 32136 25650 32172
rect 28078 38392 28134 38448
rect 28814 38004 28870 38040
rect 28814 37984 28816 38004
rect 28816 37984 28868 38004
rect 28868 37984 28870 38004
rect 28354 36780 28410 36816
rect 28354 36760 28356 36780
rect 28356 36760 28408 36780
rect 28408 36760 28410 36780
rect 26238 33516 26294 33552
rect 26238 33496 26240 33516
rect 26240 33496 26292 33516
rect 26292 33496 26294 33516
rect 26514 32408 26570 32464
rect 26330 32172 26332 32192
rect 26332 32172 26384 32192
rect 26384 32172 26386 32192
rect 26330 32136 26386 32172
rect 25318 30252 25374 30288
rect 25318 30232 25320 30252
rect 25320 30232 25372 30252
rect 25372 30232 25374 30252
rect 25410 30116 25466 30152
rect 25410 30096 25412 30116
rect 25412 30096 25464 30116
rect 25464 30096 25466 30116
rect 26054 31456 26110 31512
rect 25962 31320 26018 31376
rect 25962 31048 26018 31104
rect 25870 30912 25926 30968
rect 25778 30504 25834 30560
rect 26330 30912 26386 30968
rect 25870 30232 25926 30288
rect 25778 30116 25834 30152
rect 25778 30096 25780 30116
rect 25780 30096 25832 30116
rect 25832 30096 25834 30116
rect 25226 29844 25282 29880
rect 25226 29824 25228 29844
rect 25228 29824 25280 29844
rect 25280 29824 25282 29844
rect 24950 29416 25006 29472
rect 25042 29164 25098 29200
rect 25042 29144 25044 29164
rect 25044 29144 25096 29164
rect 25096 29144 25098 29164
rect 24674 29008 24730 29064
rect 24674 28736 24730 28792
rect 24306 27240 24362 27296
rect 23662 25608 23718 25664
rect 25318 27920 25374 27976
rect 23570 24556 23572 24576
rect 23572 24556 23624 24576
rect 23624 24556 23626 24576
rect 23570 24520 23626 24556
rect 23018 22752 23074 22808
rect 22558 21836 22560 21856
rect 22560 21836 22612 21856
rect 22612 21836 22614 21856
rect 22558 21800 22614 21836
rect 22466 20032 22522 20088
rect 22926 21800 22982 21856
rect 22650 21392 22706 21448
rect 23110 21800 23166 21856
rect 22834 21256 22890 21312
rect 22742 21120 22798 21176
rect 22834 20848 22890 20904
rect 22742 20712 22798 20768
rect 22190 17856 22246 17912
rect 23018 20440 23074 20496
rect 22926 19624 22982 19680
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 22558 16532 22560 16552
rect 22560 16532 22612 16552
rect 22612 16532 22614 16552
rect 22558 16496 22614 16532
rect 23110 19760 23166 19816
rect 22834 18128 22890 18184
rect 24214 25744 24270 25800
rect 24306 25064 24362 25120
rect 24582 24948 24638 24984
rect 24582 24928 24584 24948
rect 24584 24928 24636 24948
rect 24636 24928 24638 24948
rect 25226 25780 25228 25800
rect 25228 25780 25280 25800
rect 25280 25780 25282 25800
rect 25226 25744 25282 25780
rect 25870 27648 25926 27704
rect 23386 22072 23442 22128
rect 23294 21256 23350 21312
rect 23294 20032 23350 20088
rect 24030 21956 24086 21992
rect 24030 21936 24032 21956
rect 24032 21936 24084 21956
rect 24084 21936 24086 21956
rect 23938 21528 23994 21584
rect 24398 24656 24454 24712
rect 24306 23432 24362 23488
rect 23662 20984 23718 21040
rect 23662 20848 23718 20904
rect 24582 23160 24638 23216
rect 24398 22636 24454 22672
rect 24398 22616 24400 22636
rect 24400 22616 24452 22636
rect 24452 22616 24454 22636
rect 24858 23160 24914 23216
rect 24766 22072 24822 22128
rect 24674 21800 24730 21856
rect 23846 20712 23902 20768
rect 24030 20712 24086 20768
rect 23938 20576 23994 20632
rect 23294 19216 23350 19272
rect 23570 19760 23626 19816
rect 24030 20440 24086 20496
rect 24214 20304 24270 20360
rect 25410 23024 25466 23080
rect 25042 20984 25098 21040
rect 25318 21528 25374 21584
rect 26698 33940 26700 33960
rect 26700 33940 26752 33960
rect 26752 33940 26754 33960
rect 26698 33904 26754 33940
rect 26698 33632 26754 33688
rect 26882 34856 26938 34912
rect 27986 36352 28042 36408
rect 27986 36080 28042 36136
rect 27894 35536 27950 35592
rect 27158 34176 27214 34232
rect 26882 32136 26938 32192
rect 26974 32000 27030 32056
rect 27802 34312 27858 34368
rect 27618 34076 27620 34096
rect 27620 34076 27672 34096
rect 27672 34076 27674 34096
rect 27618 34040 27674 34076
rect 28354 36216 28410 36272
rect 28906 37168 28962 37224
rect 28722 36896 28778 36952
rect 28630 36488 28686 36544
rect 28814 36352 28870 36408
rect 29090 36524 29092 36544
rect 29092 36524 29144 36544
rect 29144 36524 29146 36544
rect 28538 35808 28594 35864
rect 27986 34060 28042 34096
rect 27986 34040 27988 34060
rect 27988 34040 28040 34060
rect 28040 34040 28042 34060
rect 28262 34312 28318 34368
rect 27618 33804 27620 33824
rect 27620 33804 27672 33824
rect 27672 33804 27674 33824
rect 27618 33768 27674 33804
rect 26514 30252 26570 30288
rect 26514 30232 26516 30252
rect 26516 30232 26568 30252
rect 26568 30232 26570 30252
rect 26422 28756 26478 28792
rect 26422 28736 26424 28756
rect 26424 28736 26476 28756
rect 26476 28736 26478 28756
rect 27066 31456 27122 31512
rect 26974 30368 27030 30424
rect 26054 26832 26110 26888
rect 25870 26288 25926 26344
rect 26514 27512 26570 27568
rect 26514 27240 26570 27296
rect 26146 25744 26202 25800
rect 26238 25608 26294 25664
rect 26514 25064 26570 25120
rect 27066 29824 27122 29880
rect 27342 31048 27398 31104
rect 27894 33224 27950 33280
rect 27802 33088 27858 33144
rect 28078 33652 28134 33688
rect 28078 33632 28080 33652
rect 28080 33632 28132 33652
rect 28132 33632 28134 33652
rect 29090 36488 29146 36524
rect 29090 36116 29092 36136
rect 29092 36116 29144 36136
rect 29144 36116 29146 36136
rect 29090 36080 29146 36116
rect 29458 36780 29514 36816
rect 29458 36760 29460 36780
rect 29460 36760 29512 36780
rect 29512 36760 29514 36780
rect 29826 37032 29882 37088
rect 29458 36624 29514 36680
rect 29090 35708 29092 35728
rect 29092 35708 29144 35728
rect 29144 35708 29146 35728
rect 29090 35672 29146 35708
rect 29274 35536 29330 35592
rect 28354 33768 28410 33824
rect 27342 29416 27398 29472
rect 27710 30504 27766 30560
rect 27342 29164 27398 29200
rect 27342 29144 27344 29164
rect 27344 29144 27396 29164
rect 27396 29144 27398 29164
rect 26790 27784 26846 27840
rect 27710 28872 27766 28928
rect 28170 30932 28226 30968
rect 28170 30912 28172 30932
rect 28172 30912 28224 30932
rect 28224 30912 28226 30932
rect 27802 28736 27858 28792
rect 27710 28328 27766 28384
rect 27250 27648 27306 27704
rect 27526 27512 27582 27568
rect 27250 27240 27306 27296
rect 26698 26152 26754 26208
rect 25778 24112 25834 24168
rect 25778 23840 25834 23896
rect 25962 23976 26018 24032
rect 26146 23840 26202 23896
rect 25594 22108 25596 22128
rect 25596 22108 25648 22128
rect 25648 22108 25650 22128
rect 25594 22072 25650 22108
rect 25594 21972 25596 21992
rect 25596 21972 25648 21992
rect 25648 21972 25650 21992
rect 25594 21936 25650 21972
rect 24582 19896 24638 19952
rect 23294 18536 23350 18592
rect 25134 20168 25190 20224
rect 24398 18944 24454 19000
rect 24122 18284 24178 18320
rect 24122 18264 24124 18284
rect 24124 18264 24176 18284
rect 24176 18264 24178 18284
rect 23846 17992 23902 18048
rect 23662 17604 23718 17640
rect 23662 17584 23664 17604
rect 23664 17584 23716 17604
rect 23716 17584 23718 17604
rect 23570 17196 23626 17232
rect 23570 17176 23572 17196
rect 23572 17176 23624 17196
rect 23624 17176 23626 17196
rect 25134 18808 25190 18864
rect 24766 18264 24822 18320
rect 25870 22500 25926 22536
rect 25870 22480 25872 22500
rect 25872 22480 25924 22500
rect 25924 22480 25926 22500
rect 26054 23432 26110 23488
rect 26330 23160 26386 23216
rect 25962 22208 26018 22264
rect 25778 21548 25834 21584
rect 25778 21528 25780 21548
rect 25780 21528 25832 21548
rect 25832 21528 25834 21548
rect 26238 21936 26294 21992
rect 25502 18672 25558 18728
rect 25686 17856 25742 17912
rect 25962 19624 26018 19680
rect 25962 18944 26018 19000
rect 26238 20324 26294 20360
rect 26238 20304 26240 20324
rect 26240 20304 26292 20324
rect 26292 20304 26294 20324
rect 26422 20984 26478 21040
rect 26882 24112 26938 24168
rect 27342 26288 27398 26344
rect 27250 25744 27306 25800
rect 27158 23432 27214 23488
rect 26514 20848 26570 20904
rect 26606 20576 26662 20632
rect 26882 20712 26938 20768
rect 28814 32716 28816 32736
rect 28816 32716 28868 32736
rect 28868 32716 28870 32736
rect 28814 32680 28870 32716
rect 28722 30812 28724 30832
rect 28724 30812 28776 30832
rect 28776 30812 28778 30832
rect 28722 30776 28778 30812
rect 29274 32972 29330 33008
rect 29734 36372 29790 36408
rect 29734 36352 29736 36372
rect 29736 36352 29788 36372
rect 29788 36352 29790 36372
rect 29918 36216 29974 36272
rect 30102 35672 30158 35728
rect 30286 36488 30342 36544
rect 31114 36080 31170 36136
rect 29274 32952 29276 32972
rect 29276 32952 29328 32972
rect 29328 32952 29330 32972
rect 28722 30096 28778 30152
rect 28538 29280 28594 29336
rect 28814 29416 28870 29472
rect 28630 28872 28686 28928
rect 29090 29960 29146 30016
rect 29366 29824 29422 29880
rect 29274 29280 29330 29336
rect 28170 27784 28226 27840
rect 28078 26832 28134 26888
rect 27158 20440 27214 20496
rect 26238 19080 26294 19136
rect 25594 17448 25650 17504
rect 27342 20032 27398 20088
rect 27986 25356 28042 25392
rect 27986 25336 27988 25356
rect 27988 25336 28040 25356
rect 28040 25336 28042 25356
rect 27894 23296 27950 23352
rect 27894 22752 27950 22808
rect 27342 19760 27398 19816
rect 26698 17720 26754 17776
rect 28262 26696 28318 26752
rect 28170 24520 28226 24576
rect 28630 26288 28686 26344
rect 28446 23704 28502 23760
rect 29458 29164 29514 29200
rect 29458 29144 29460 29164
rect 29460 29144 29512 29164
rect 29512 29144 29514 29164
rect 29550 29008 29606 29064
rect 29274 26424 29330 26480
rect 29918 31592 29974 31648
rect 30194 29688 30250 29744
rect 31666 30640 31722 30696
rect 30562 29688 30618 29744
rect 30102 29044 30104 29064
rect 30104 29044 30156 29064
rect 30156 29044 30158 29064
rect 30102 29008 30158 29044
rect 32310 37984 32366 38040
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 32218 37032 32274 37088
rect 32126 36896 32182 36952
rect 31942 35980 31944 36000
rect 31944 35980 31996 36000
rect 31996 35980 31998 36000
rect 31942 35944 31998 35980
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 33322 37168 33378 37224
rect 32310 36100 32366 36136
rect 32310 36080 32312 36100
rect 32312 36080 32364 36100
rect 32364 36080 32366 36100
rect 32126 31864 32182 31920
rect 31942 29552 31998 29608
rect 31482 28600 31538 28656
rect 31390 28500 31392 28520
rect 31392 28500 31444 28520
rect 31444 28500 31446 28520
rect 31390 28464 31446 28500
rect 30746 27240 30802 27296
rect 30378 26968 30434 27024
rect 30102 26560 30158 26616
rect 28906 26152 28962 26208
rect 28630 25744 28686 25800
rect 28538 23024 28594 23080
rect 28262 22888 28318 22944
rect 28354 22480 28410 22536
rect 28538 22344 28594 22400
rect 28262 20460 28318 20496
rect 28262 20440 28264 20460
rect 28264 20440 28316 20460
rect 28316 20440 28318 20460
rect 28078 20204 28080 20224
rect 28080 20204 28132 20224
rect 28132 20204 28134 20224
rect 28078 20168 28134 20204
rect 28538 21528 28594 21584
rect 30010 25236 30012 25256
rect 30012 25236 30064 25256
rect 30064 25236 30066 25256
rect 30010 25200 30066 25236
rect 29734 25064 29790 25120
rect 31758 27548 31760 27568
rect 31760 27548 31812 27568
rect 31812 27548 31814 27568
rect 31758 27512 31814 27548
rect 31758 27104 31814 27160
rect 30930 25880 30986 25936
rect 32678 27240 32734 27296
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 33046 27548 33048 27568
rect 33048 27548 33100 27568
rect 33100 27548 33102 27568
rect 33046 27512 33102 27548
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 32494 25880 32550 25936
rect 32954 25492 33010 25528
rect 32954 25472 32956 25492
rect 32956 25472 33008 25492
rect 33008 25472 33010 25492
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 42154 31184 42210 31240
rect 43810 39208 43866 39264
rect 43810 28076 43866 28112
rect 43810 28056 43812 28076
rect 43812 28056 43864 28076
rect 43864 28056 43866 28076
rect 40682 27376 40738 27432
rect 31482 23568 31538 23624
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 30194 21664 30250 21720
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 29642 19760 29698 19816
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 29090 18964 29146 19000
rect 29090 18944 29092 18964
rect 29092 18944 29144 18964
rect 29144 18944 29146 18964
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 43166 16904 43222 16960
rect 40682 5752 40738 5808
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 1214 4392 1270 4448
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 3146 3984 3202 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 1214 3304 1270 3360
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 24674 2644 24730 2680
rect 24674 2624 24676 2644
rect 24676 2624 24728 2644
rect 24728 2624 24730 2644
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 0 41442 800 41472
rect 933 41442 999 41445
rect 0 41440 999 41442
rect 0 41384 938 41440
rect 994 41384 999 41440
rect 0 41382 999 41384
rect 0 41352 800 41382
rect 933 41379 999 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 0 40354 800 40384
rect 933 40354 999 40357
rect 0 40352 999 40354
rect 0 40296 938 40352
rect 994 40296 999 40352
rect 0 40294 999 40296
rect 0 40264 800 40294
rect 933 40291 999 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39266 800 39296
rect 1209 39266 1275 39269
rect 0 39264 1275 39266
rect 0 39208 1214 39264
rect 1270 39208 1275 39264
rect 0 39206 1275 39208
rect 0 39176 800 39206
rect 1209 39203 1275 39206
rect 43805 39266 43871 39269
rect 44200 39266 45000 39296
rect 43805 39264 45000 39266
rect 43805 39208 43810 39264
rect 43866 39208 45000 39264
rect 43805 39206 45000 39208
rect 43805 39203 43871 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 44200 39176 45000 39206
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 21173 38586 21239 38589
rect 21909 38586 21975 38589
rect 21173 38584 21975 38586
rect 21173 38528 21178 38584
rect 21234 38528 21914 38584
rect 21970 38528 21975 38584
rect 21173 38526 21975 38528
rect 21173 38523 21239 38526
rect 21909 38523 21975 38526
rect 10358 38388 10364 38452
rect 10428 38450 10434 38452
rect 20713 38450 20779 38453
rect 10428 38448 20779 38450
rect 10428 38392 20718 38448
rect 20774 38392 20779 38448
rect 10428 38390 20779 38392
rect 10428 38388 10434 38390
rect 20713 38387 20779 38390
rect 21633 38450 21699 38453
rect 28073 38450 28139 38453
rect 21633 38448 28139 38450
rect 21633 38392 21638 38448
rect 21694 38392 28078 38448
rect 28134 38392 28139 38448
rect 21633 38390 28139 38392
rect 21633 38387 21699 38390
rect 28073 38387 28139 38390
rect 0 38178 800 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 800 38118
rect 1209 38115 1275 38118
rect 21265 38178 21331 38181
rect 25405 38178 25471 38181
rect 21265 38176 25471 38178
rect 21265 38120 21270 38176
rect 21326 38120 25410 38176
rect 25466 38120 25471 38176
rect 21265 38118 25471 38120
rect 21265 38115 21331 38118
rect 25405 38115 25471 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 28809 38042 28875 38045
rect 32305 38042 32371 38045
rect 28809 38040 32371 38042
rect 28809 37984 28814 38040
rect 28870 37984 32310 38040
rect 32366 37984 32371 38040
rect 28809 37982 32371 37984
rect 28809 37979 28875 37982
rect 32305 37979 32371 37982
rect 14917 37770 14983 37773
rect 17217 37770 17283 37773
rect 14917 37768 17283 37770
rect 14917 37712 14922 37768
rect 14978 37712 17222 37768
rect 17278 37712 17283 37768
rect 14917 37710 17283 37712
rect 14917 37707 14983 37710
rect 17217 37707 17283 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 17217 37226 17283 37229
rect 19241 37226 19307 37229
rect 17217 37224 19307 37226
rect 17217 37168 17222 37224
rect 17278 37168 19246 37224
rect 19302 37168 19307 37224
rect 17217 37166 19307 37168
rect 17217 37163 17283 37166
rect 19241 37163 19307 37166
rect 24209 37226 24275 37229
rect 28901 37226 28967 37229
rect 33317 37226 33383 37229
rect 24209 37224 33383 37226
rect 24209 37168 24214 37224
rect 24270 37168 28906 37224
rect 28962 37168 33322 37224
rect 33378 37168 33383 37224
rect 24209 37166 33383 37168
rect 24209 37163 24275 37166
rect 28901 37163 28967 37166
rect 33317 37163 33383 37166
rect 0 37090 800 37120
rect 1209 37090 1275 37093
rect 0 37088 1275 37090
rect 0 37032 1214 37088
rect 1270 37032 1275 37088
rect 0 37030 1275 37032
rect 0 37000 800 37030
rect 1209 37027 1275 37030
rect 15837 37090 15903 37093
rect 17033 37090 17099 37093
rect 15837 37088 17099 37090
rect 15837 37032 15842 37088
rect 15898 37032 17038 37088
rect 17094 37032 17099 37088
rect 15837 37030 17099 37032
rect 15837 37027 15903 37030
rect 17033 37027 17099 37030
rect 29821 37090 29887 37093
rect 32213 37090 32279 37093
rect 29821 37088 32279 37090
rect 29821 37032 29826 37088
rect 29882 37032 32218 37088
rect 32274 37032 32279 37088
rect 29821 37030 32279 37032
rect 29821 37027 29887 37030
rect 32213 37027 32279 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 28717 36954 28783 36957
rect 32121 36954 32187 36957
rect 28717 36952 32187 36954
rect 28717 36896 28722 36952
rect 28778 36896 32126 36952
rect 32182 36896 32187 36952
rect 28717 36894 32187 36896
rect 28717 36891 28783 36894
rect 32121 36891 32187 36894
rect 14273 36818 14339 36821
rect 14917 36818 14983 36821
rect 14273 36816 14983 36818
rect 14273 36760 14278 36816
rect 14334 36760 14922 36816
rect 14978 36760 14983 36816
rect 14273 36758 14983 36760
rect 14273 36755 14339 36758
rect 14917 36755 14983 36758
rect 28349 36818 28415 36821
rect 29453 36818 29519 36821
rect 28349 36816 29519 36818
rect 28349 36760 28354 36816
rect 28410 36760 29458 36816
rect 29514 36760 29519 36816
rect 28349 36758 29519 36760
rect 28349 36755 28415 36758
rect 29453 36755 29519 36758
rect 23105 36682 23171 36685
rect 29453 36682 29519 36685
rect 23105 36680 29519 36682
rect 23105 36624 23110 36680
rect 23166 36624 29458 36680
rect 29514 36624 29519 36680
rect 23105 36622 29519 36624
rect 23105 36619 23171 36622
rect 29453 36619 29519 36622
rect 28625 36546 28691 36549
rect 11102 36544 28691 36546
rect 11102 36488 28630 36544
rect 28686 36488 28691 36544
rect 11102 36486 28691 36488
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 8293 36138 8359 36141
rect 9305 36138 9371 36141
rect 10961 36138 11027 36141
rect 11102 36138 11162 36486
rect 28625 36483 28691 36486
rect 29085 36546 29151 36549
rect 30281 36546 30347 36549
rect 29085 36544 30347 36546
rect 29085 36488 29090 36544
rect 29146 36488 30286 36544
rect 30342 36488 30347 36544
rect 29085 36486 30347 36488
rect 29085 36483 29151 36486
rect 30281 36483 30347 36486
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 26417 36410 26483 36413
rect 27981 36410 28047 36413
rect 26417 36408 28047 36410
rect 26417 36352 26422 36408
rect 26478 36352 27986 36408
rect 28042 36352 28047 36408
rect 26417 36350 28047 36352
rect 26417 36347 26483 36350
rect 27981 36347 28047 36350
rect 28809 36410 28875 36413
rect 29729 36410 29795 36413
rect 28809 36408 29795 36410
rect 28809 36352 28814 36408
rect 28870 36352 29734 36408
rect 29790 36352 29795 36408
rect 28809 36350 29795 36352
rect 28809 36347 28875 36350
rect 29729 36347 29795 36350
rect 28349 36274 28415 36277
rect 29913 36274 29979 36277
rect 8212 36136 10794 36138
rect 8212 36080 8298 36136
rect 8354 36080 9310 36136
rect 9366 36080 10794 36136
rect 8212 36078 10794 36080
rect 8293 36075 8402 36078
rect 9305 36075 9371 36078
rect 0 36002 800 36032
rect 933 36002 999 36005
rect 8342 36004 8402 36075
rect 0 36000 999 36002
rect 0 35944 938 36000
rect 994 35944 999 36000
rect 0 35942 999 35944
rect 0 35912 800 35942
rect 933 35939 999 35942
rect 8334 35940 8340 36004
rect 8404 35940 8410 36004
rect 10734 36002 10794 36078
rect 10961 36136 11162 36138
rect 10961 36080 10966 36136
rect 11022 36080 11162 36136
rect 10961 36078 11162 36080
rect 12390 36272 31770 36274
rect 12390 36216 28354 36272
rect 28410 36216 29918 36272
rect 29974 36216 31770 36272
rect 12390 36214 31770 36216
rect 10961 36075 11027 36078
rect 12390 36002 12450 36214
rect 28349 36211 28415 36214
rect 29913 36211 29979 36214
rect 14733 36138 14799 36141
rect 17493 36138 17559 36141
rect 14733 36136 17559 36138
rect 14733 36080 14738 36136
rect 14794 36080 17498 36136
rect 17554 36080 17559 36136
rect 14733 36078 17559 36080
rect 14733 36075 14799 36078
rect 17493 36075 17559 36078
rect 27981 36138 28047 36141
rect 29085 36138 29151 36141
rect 31109 36138 31175 36141
rect 27981 36136 28090 36138
rect 27981 36080 27986 36136
rect 28042 36080 28090 36136
rect 27981 36075 28090 36080
rect 29085 36136 31175 36138
rect 29085 36080 29090 36136
rect 29146 36080 31114 36136
rect 31170 36080 31175 36136
rect 29085 36078 31175 36080
rect 31710 36138 31770 36214
rect 32305 36138 32371 36141
rect 31710 36136 32371 36138
rect 31710 36080 32310 36136
rect 32366 36080 32371 36136
rect 31710 36078 32371 36080
rect 29085 36075 29151 36078
rect 31109 36075 31175 36078
rect 32305 36075 32371 36078
rect 10734 35942 12450 36002
rect 25405 36002 25471 36005
rect 25630 36002 25636 36004
rect 25405 36000 25636 36002
rect 25405 35944 25410 36000
rect 25466 35944 25636 36000
rect 25405 35942 25636 35944
rect 25405 35939 25471 35942
rect 25630 35940 25636 35942
rect 25700 35940 25706 36004
rect 28030 36002 28090 36075
rect 31937 36002 32003 36005
rect 28030 36000 32003 36002
rect 28030 35944 31942 36000
rect 31998 35944 32003 36000
rect 28030 35942 32003 35944
rect 31937 35939 32003 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 25957 35866 26023 35869
rect 28533 35866 28599 35869
rect 25957 35864 28599 35866
rect 25957 35808 25962 35864
rect 26018 35808 28538 35864
rect 28594 35808 28599 35864
rect 25957 35806 28599 35808
rect 25957 35803 26023 35806
rect 28533 35803 28599 35806
rect 9673 35730 9739 35733
rect 29085 35730 29151 35733
rect 30097 35730 30163 35733
rect 9673 35728 30163 35730
rect 9673 35672 9678 35728
rect 9734 35672 29090 35728
rect 29146 35672 30102 35728
rect 30158 35672 30163 35728
rect 9673 35670 30163 35672
rect 9673 35667 9739 35670
rect 29085 35667 29151 35670
rect 30097 35667 30163 35670
rect 13261 35594 13327 35597
rect 17125 35594 17191 35597
rect 13261 35592 17191 35594
rect 13261 35536 13266 35592
rect 13322 35536 17130 35592
rect 17186 35536 17191 35592
rect 13261 35534 17191 35536
rect 13261 35531 13327 35534
rect 17125 35531 17191 35534
rect 27889 35594 27955 35597
rect 29269 35594 29335 35597
rect 27889 35592 29335 35594
rect 27889 35536 27894 35592
rect 27950 35536 29274 35592
rect 29330 35536 29335 35592
rect 27889 35534 29335 35536
rect 27889 35531 27955 35534
rect 29269 35531 29335 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 9438 35124 9444 35188
rect 9508 35186 9514 35188
rect 9673 35186 9739 35189
rect 9508 35184 9739 35186
rect 9508 35128 9678 35184
rect 9734 35128 9739 35184
rect 9508 35126 9739 35128
rect 9508 35124 9514 35126
rect 9673 35123 9739 35126
rect 11789 35186 11855 35189
rect 23473 35186 23539 35189
rect 11789 35184 23539 35186
rect 11789 35128 11794 35184
rect 11850 35128 23478 35184
rect 23534 35128 23539 35184
rect 11789 35126 23539 35128
rect 11789 35123 11855 35126
rect 23473 35123 23539 35126
rect 0 34914 800 34944
rect 933 34914 999 34917
rect 0 34912 999 34914
rect 0 34856 938 34912
rect 994 34856 999 34912
rect 0 34854 999 34856
rect 0 34824 800 34854
rect 933 34851 999 34854
rect 19977 34914 20043 34917
rect 26877 34914 26943 34917
rect 19977 34912 26943 34914
rect 19977 34856 19982 34912
rect 20038 34856 26882 34912
rect 26938 34856 26943 34912
rect 19977 34854 26943 34856
rect 19977 34851 20043 34854
rect 26877 34851 26943 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 8150 34716 8156 34780
rect 8220 34778 8226 34780
rect 10961 34778 11027 34781
rect 8220 34776 11027 34778
rect 8220 34720 10966 34776
rect 11022 34720 11027 34776
rect 8220 34718 11027 34720
rect 8220 34716 8226 34718
rect 10961 34715 11027 34718
rect 12065 34778 12131 34781
rect 15009 34778 15075 34781
rect 12065 34776 15075 34778
rect 12065 34720 12070 34776
rect 12126 34720 15014 34776
rect 15070 34720 15075 34776
rect 12065 34718 15075 34720
rect 12065 34715 12131 34718
rect 15009 34715 15075 34718
rect 11462 34580 11468 34644
rect 11532 34642 11538 34644
rect 11789 34642 11855 34645
rect 11532 34640 11855 34642
rect 11532 34584 11794 34640
rect 11850 34584 11855 34640
rect 11532 34582 11855 34584
rect 11532 34580 11538 34582
rect 11789 34579 11855 34582
rect 12157 34642 12223 34645
rect 16757 34642 16823 34645
rect 18505 34642 18571 34645
rect 12157 34640 15394 34642
rect 12157 34584 12162 34640
rect 12218 34584 15394 34640
rect 12157 34582 15394 34584
rect 12157 34579 12223 34582
rect 15334 34509 15394 34582
rect 16757 34640 18571 34642
rect 16757 34584 16762 34640
rect 16818 34584 18510 34640
rect 18566 34584 18571 34640
rect 16757 34582 18571 34584
rect 16757 34579 16823 34582
rect 18505 34579 18571 34582
rect 21265 34642 21331 34645
rect 22369 34642 22435 34645
rect 23013 34642 23079 34645
rect 21265 34640 23079 34642
rect 21265 34584 21270 34640
rect 21326 34584 22374 34640
rect 22430 34584 23018 34640
rect 23074 34584 23079 34640
rect 21265 34582 23079 34584
rect 21265 34579 21331 34582
rect 22369 34579 22435 34582
rect 23013 34579 23079 34582
rect 5901 34506 5967 34509
rect 11830 34506 11836 34508
rect 5901 34504 11836 34506
rect 5901 34448 5906 34504
rect 5962 34448 11836 34504
rect 5901 34446 11836 34448
rect 5901 34443 5967 34446
rect 11830 34444 11836 34446
rect 11900 34444 11906 34508
rect 15334 34504 15443 34509
rect 15334 34448 15382 34504
rect 15438 34448 15443 34504
rect 15334 34446 15443 34448
rect 15377 34443 15443 34446
rect 27797 34370 27863 34373
rect 28257 34370 28323 34373
rect 27797 34368 28323 34370
rect 27797 34312 27802 34368
rect 27858 34312 28262 34368
rect 28318 34312 28323 34368
rect 27797 34310 28323 34312
rect 27797 34307 27863 34310
rect 28257 34307 28323 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 6177 34234 6243 34237
rect 8569 34234 8635 34237
rect 6177 34232 8635 34234
rect 6177 34176 6182 34232
rect 6238 34176 8574 34232
rect 8630 34176 8635 34232
rect 6177 34174 8635 34176
rect 6177 34171 6243 34174
rect 8569 34171 8635 34174
rect 14917 34234 14983 34237
rect 25037 34234 25103 34237
rect 14917 34232 25103 34234
rect 14917 34176 14922 34232
rect 14978 34176 25042 34232
rect 25098 34176 25103 34232
rect 14917 34174 25103 34176
rect 14917 34171 14983 34174
rect 25037 34171 25103 34174
rect 25446 34172 25452 34236
rect 25516 34234 25522 34236
rect 25589 34234 25655 34237
rect 27153 34234 27219 34237
rect 25516 34232 27219 34234
rect 25516 34176 25594 34232
rect 25650 34176 27158 34232
rect 27214 34176 27219 34232
rect 25516 34174 27219 34176
rect 25516 34172 25522 34174
rect 25589 34171 25655 34174
rect 27153 34171 27219 34174
rect 11697 34098 11763 34101
rect 13261 34098 13327 34101
rect 25681 34098 25747 34101
rect 11697 34096 25747 34098
rect 11697 34040 11702 34096
rect 11758 34040 13266 34096
rect 13322 34040 25686 34096
rect 25742 34040 25747 34096
rect 11697 34038 25747 34040
rect 11697 34035 11763 34038
rect 13261 34035 13327 34038
rect 25681 34035 25747 34038
rect 27613 34098 27679 34101
rect 27981 34098 28047 34101
rect 27613 34096 28047 34098
rect 27613 34040 27618 34096
rect 27674 34040 27986 34096
rect 28042 34040 28047 34096
rect 27613 34038 28047 34040
rect 27613 34035 27679 34038
rect 27981 34035 28047 34038
rect 10501 33962 10567 33965
rect 12433 33962 12499 33965
rect 10501 33960 12499 33962
rect 10501 33904 10506 33960
rect 10562 33904 12438 33960
rect 12494 33904 12499 33960
rect 10501 33902 12499 33904
rect 10501 33899 10567 33902
rect 12433 33899 12499 33902
rect 24669 33962 24735 33965
rect 26693 33962 26759 33965
rect 24669 33960 26759 33962
rect 24669 33904 24674 33960
rect 24730 33904 26698 33960
rect 26754 33904 26759 33960
rect 24669 33902 26759 33904
rect 24669 33899 24735 33902
rect 26693 33899 26759 33902
rect 0 33826 800 33856
rect 933 33826 999 33829
rect 0 33824 999 33826
rect 0 33768 938 33824
rect 994 33768 999 33824
rect 0 33766 999 33768
rect 0 33736 800 33766
rect 933 33763 999 33766
rect 21173 33826 21239 33829
rect 24853 33826 24919 33829
rect 21173 33824 24919 33826
rect 21173 33768 21178 33824
rect 21234 33768 24858 33824
rect 24914 33768 24919 33824
rect 21173 33766 24919 33768
rect 21173 33763 21239 33766
rect 24853 33763 24919 33766
rect 27613 33826 27679 33829
rect 28349 33826 28415 33829
rect 27613 33824 28415 33826
rect 27613 33768 27618 33824
rect 27674 33768 28354 33824
rect 28410 33768 28415 33824
rect 27613 33766 28415 33768
rect 27613 33763 27679 33766
rect 28349 33763 28415 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 13169 33690 13235 33693
rect 12252 33688 13235 33690
rect 12252 33632 13174 33688
rect 13230 33632 13235 33688
rect 12252 33630 13235 33632
rect 12252 33557 12312 33630
rect 13169 33627 13235 33630
rect 24025 33690 24091 33693
rect 25497 33690 25563 33693
rect 24025 33688 25563 33690
rect 24025 33632 24030 33688
rect 24086 33632 25502 33688
rect 25558 33632 25563 33688
rect 24025 33630 25563 33632
rect 24025 33627 24091 33630
rect 25497 33627 25563 33630
rect 26693 33690 26759 33693
rect 28073 33690 28139 33693
rect 26693 33688 28139 33690
rect 26693 33632 26698 33688
rect 26754 33632 28078 33688
rect 28134 33632 28139 33688
rect 26693 33630 28139 33632
rect 26693 33627 26759 33630
rect 28073 33627 28139 33630
rect 11329 33554 11395 33557
rect 12249 33554 12315 33557
rect 11329 33552 12315 33554
rect 11329 33496 11334 33552
rect 11390 33496 12254 33552
rect 12310 33496 12315 33552
rect 11329 33494 12315 33496
rect 11329 33491 11395 33494
rect 12249 33491 12315 33494
rect 23289 33554 23355 33557
rect 26233 33554 26299 33557
rect 26366 33554 26372 33556
rect 23289 33552 26372 33554
rect 23289 33496 23294 33552
rect 23350 33496 26238 33552
rect 26294 33496 26372 33552
rect 23289 33494 26372 33496
rect 23289 33491 23355 33494
rect 26233 33491 26299 33494
rect 26366 33492 26372 33494
rect 26436 33492 26442 33556
rect 11697 33418 11763 33421
rect 12709 33418 12775 33421
rect 11697 33416 12775 33418
rect 11697 33360 11702 33416
rect 11758 33360 12714 33416
rect 12770 33360 12775 33416
rect 11697 33358 12775 33360
rect 11697 33355 11763 33358
rect 12709 33355 12775 33358
rect 13261 33418 13327 33421
rect 15653 33418 15719 33421
rect 24945 33420 25011 33421
rect 13261 33416 15719 33418
rect 13261 33360 13266 33416
rect 13322 33360 15658 33416
rect 15714 33360 15719 33416
rect 13261 33358 15719 33360
rect 13261 33355 13327 33358
rect 15653 33355 15719 33358
rect 24894 33356 24900 33420
rect 24964 33418 25011 33420
rect 24964 33416 25056 33418
rect 25006 33360 25056 33416
rect 24964 33358 25056 33360
rect 24964 33356 25011 33358
rect 24945 33355 25011 33356
rect 10961 33282 11027 33285
rect 13629 33282 13695 33285
rect 15377 33282 15443 33285
rect 10961 33280 15443 33282
rect 10961 33224 10966 33280
rect 11022 33224 13634 33280
rect 13690 33224 15382 33280
rect 15438 33224 15443 33280
rect 10961 33222 15443 33224
rect 10961 33219 11027 33222
rect 13629 33219 13695 33222
rect 15377 33219 15443 33222
rect 21541 33282 21607 33285
rect 27889 33282 27955 33285
rect 21541 33280 27955 33282
rect 21541 33224 21546 33280
rect 21602 33224 27894 33280
rect 27950 33224 27955 33280
rect 21541 33222 27955 33224
rect 21541 33219 21607 33222
rect 27889 33219 27955 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 9765 33146 9831 33149
rect 13629 33146 13695 33149
rect 9765 33144 13695 33146
rect 9765 33088 9770 33144
rect 9826 33088 13634 33144
rect 13690 33088 13695 33144
rect 9765 33086 13695 33088
rect 9765 33083 9831 33086
rect 13629 33083 13695 33086
rect 27654 33084 27660 33148
rect 27724 33146 27730 33148
rect 27797 33146 27863 33149
rect 27724 33144 27863 33146
rect 27724 33088 27802 33144
rect 27858 33088 27863 33144
rect 27724 33086 27863 33088
rect 27724 33084 27730 33086
rect 27797 33083 27863 33086
rect 2681 33010 2747 33013
rect 21357 33010 21423 33013
rect 2681 33008 21423 33010
rect 2681 32952 2686 33008
rect 2742 32952 21362 33008
rect 21418 32952 21423 33008
rect 2681 32950 21423 32952
rect 2681 32947 2747 32950
rect 21357 32947 21423 32950
rect 23657 33010 23723 33013
rect 29269 33010 29335 33013
rect 23657 33008 29335 33010
rect 23657 32952 23662 33008
rect 23718 32952 29274 33008
rect 29330 32952 29335 33008
rect 23657 32950 29335 32952
rect 23657 32947 23723 32950
rect 29269 32947 29335 32950
rect 10317 32874 10383 32877
rect 18873 32874 18939 32877
rect 10317 32872 18939 32874
rect 10317 32816 10322 32872
rect 10378 32816 18878 32872
rect 18934 32816 18939 32872
rect 10317 32814 18939 32816
rect 10317 32811 10383 32814
rect 18873 32811 18939 32814
rect 0 32738 800 32768
rect 933 32738 999 32741
rect 18505 32740 18571 32741
rect 18454 32738 18460 32740
rect 0 32736 999 32738
rect 0 32680 938 32736
rect 994 32680 999 32736
rect 0 32678 999 32680
rect 18414 32678 18460 32738
rect 18524 32736 18571 32740
rect 18566 32680 18571 32736
rect 0 32648 800 32678
rect 933 32675 999 32678
rect 18454 32676 18460 32678
rect 18524 32676 18571 32680
rect 28574 32676 28580 32740
rect 28644 32738 28650 32740
rect 28809 32738 28875 32741
rect 28644 32736 28875 32738
rect 28644 32680 28814 32736
rect 28870 32680 28875 32736
rect 28644 32678 28875 32680
rect 28644 32676 28650 32678
rect 18505 32675 18571 32676
rect 28809 32675 28875 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 13629 32602 13695 32605
rect 15377 32602 15443 32605
rect 16021 32602 16087 32605
rect 13629 32600 16087 32602
rect 13629 32544 13634 32600
rect 13690 32544 15382 32600
rect 15438 32544 16026 32600
rect 16082 32544 16087 32600
rect 13629 32542 16087 32544
rect 13629 32539 13695 32542
rect 15377 32539 15443 32542
rect 16021 32539 16087 32542
rect 13997 32466 14063 32469
rect 16757 32466 16823 32469
rect 26509 32466 26575 32469
rect 13997 32464 16823 32466
rect 13997 32408 14002 32464
rect 14058 32408 16762 32464
rect 16818 32408 16823 32464
rect 13997 32406 16823 32408
rect 13997 32403 14063 32406
rect 16757 32403 16823 32406
rect 26374 32464 26575 32466
rect 26374 32408 26514 32464
rect 26570 32408 26575 32464
rect 26374 32406 26575 32408
rect 13537 32330 13603 32333
rect 14825 32330 14891 32333
rect 26374 32330 26434 32406
rect 26509 32403 26575 32406
rect 13537 32328 14891 32330
rect 13537 32272 13542 32328
rect 13598 32272 14830 32328
rect 14886 32272 14891 32328
rect 13537 32270 14891 32272
rect 13537 32267 13603 32270
rect 14825 32267 14891 32270
rect 26190 32270 26434 32330
rect 12985 32194 13051 32197
rect 15469 32194 15535 32197
rect 12985 32192 15535 32194
rect 12985 32136 12990 32192
rect 13046 32136 15474 32192
rect 15530 32136 15535 32192
rect 12985 32134 15535 32136
rect 12985 32131 13051 32134
rect 15469 32131 15535 32134
rect 24669 32194 24735 32197
rect 25589 32194 25655 32197
rect 24669 32192 25655 32194
rect 24669 32136 24674 32192
rect 24730 32136 25594 32192
rect 25650 32136 25655 32192
rect 24669 32134 25655 32136
rect 24669 32131 24735 32134
rect 25589 32131 25655 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 6126 31996 6132 32060
rect 6196 32058 6202 32060
rect 14549 32058 14615 32061
rect 6196 32056 14615 32058
rect 6196 32000 14554 32056
rect 14610 32000 14615 32056
rect 6196 31998 14615 32000
rect 6196 31996 6202 31998
rect 4153 31922 4219 31925
rect 6134 31922 6194 31996
rect 14549 31995 14615 31998
rect 18689 32058 18755 32061
rect 23933 32058 23999 32061
rect 18689 32056 23999 32058
rect 18689 32000 18694 32056
rect 18750 32000 23938 32056
rect 23994 32000 23999 32056
rect 18689 31998 23999 32000
rect 18689 31995 18755 31998
rect 23933 31995 23999 31998
rect 25221 32058 25287 32061
rect 25814 32058 25820 32060
rect 25221 32056 25820 32058
rect 25221 32000 25226 32056
rect 25282 32000 25820 32056
rect 25221 31998 25820 32000
rect 25221 31995 25287 31998
rect 25814 31996 25820 31998
rect 25884 31996 25890 32060
rect 26190 32058 26250 32270
rect 26325 32194 26391 32197
rect 26877 32194 26943 32197
rect 26325 32192 26943 32194
rect 26325 32136 26330 32192
rect 26386 32136 26882 32192
rect 26938 32136 26943 32192
rect 26325 32134 26943 32136
rect 26325 32131 26391 32134
rect 26877 32131 26943 32134
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 26969 32058 27035 32061
rect 26190 32056 27035 32058
rect 26190 32000 26974 32056
rect 27030 32000 27035 32056
rect 26190 31998 27035 32000
rect 26969 31995 27035 31998
rect 4153 31920 6194 31922
rect 4153 31864 4158 31920
rect 4214 31864 6194 31920
rect 4153 31862 6194 31864
rect 14365 31922 14431 31925
rect 18045 31922 18111 31925
rect 32121 31922 32187 31925
rect 14365 31920 32187 31922
rect 14365 31864 14370 31920
rect 14426 31864 18050 31920
rect 18106 31864 32126 31920
rect 32182 31864 32187 31920
rect 14365 31862 32187 31864
rect 4153 31859 4219 31862
rect 14365 31859 14431 31862
rect 18045 31859 18111 31862
rect 32121 31859 32187 31862
rect 9673 31786 9739 31789
rect 15837 31786 15903 31789
rect 9673 31784 15903 31786
rect 9673 31728 9678 31784
rect 9734 31728 15842 31784
rect 15898 31728 15903 31784
rect 9673 31726 15903 31728
rect 9673 31723 9739 31726
rect 15837 31723 15903 31726
rect 0 31650 800 31680
rect 1485 31650 1551 31653
rect 0 31648 1551 31650
rect 0 31592 1490 31648
rect 1546 31592 1551 31648
rect 0 31590 1551 31592
rect 0 31560 800 31590
rect 1485 31587 1551 31590
rect 10593 31650 10659 31653
rect 12249 31650 12315 31653
rect 10593 31648 12315 31650
rect 10593 31592 10598 31648
rect 10654 31592 12254 31648
rect 12310 31592 12315 31648
rect 10593 31590 12315 31592
rect 10593 31587 10659 31590
rect 12249 31587 12315 31590
rect 24025 31650 24091 31653
rect 29913 31650 29979 31653
rect 24025 31648 29979 31650
rect 24025 31592 24030 31648
rect 24086 31592 29918 31648
rect 29974 31592 29979 31648
rect 24025 31590 29979 31592
rect 24025 31587 24091 31590
rect 29913 31587 29979 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 24945 31514 25011 31517
rect 25262 31514 25268 31516
rect 24945 31512 25268 31514
rect 24945 31456 24950 31512
rect 25006 31456 25268 31512
rect 24945 31454 25268 31456
rect 24945 31451 25011 31454
rect 25262 31452 25268 31454
rect 25332 31514 25338 31516
rect 26049 31514 26115 31517
rect 27061 31514 27127 31517
rect 25332 31512 27127 31514
rect 25332 31456 26054 31512
rect 26110 31456 27066 31512
rect 27122 31456 27127 31512
rect 25332 31454 27127 31456
rect 25332 31452 25338 31454
rect 26049 31451 26115 31454
rect 27061 31451 27127 31454
rect 5533 31378 5599 31381
rect 8937 31378 9003 31381
rect 5533 31376 9003 31378
rect 5533 31320 5538 31376
rect 5594 31320 8942 31376
rect 8998 31320 9003 31376
rect 5533 31318 9003 31320
rect 5533 31315 5599 31318
rect 8937 31315 9003 31318
rect 13629 31378 13695 31381
rect 18086 31378 18092 31380
rect 13629 31376 18092 31378
rect 13629 31320 13634 31376
rect 13690 31320 18092 31376
rect 13629 31318 18092 31320
rect 13629 31315 13695 31318
rect 18086 31316 18092 31318
rect 18156 31378 18162 31380
rect 19149 31378 19215 31381
rect 20161 31378 20227 31381
rect 18156 31376 20227 31378
rect 18156 31320 19154 31376
rect 19210 31320 20166 31376
rect 20222 31320 20227 31376
rect 18156 31318 20227 31320
rect 18156 31316 18162 31318
rect 19149 31315 19215 31318
rect 20161 31315 20227 31318
rect 24301 31378 24367 31381
rect 25957 31378 26023 31381
rect 24301 31376 26023 31378
rect 24301 31320 24306 31376
rect 24362 31320 25962 31376
rect 26018 31320 26023 31376
rect 24301 31318 26023 31320
rect 24301 31315 24367 31318
rect 25957 31315 26023 31318
rect 17677 31242 17743 31245
rect 19149 31242 19215 31245
rect 17677 31240 19215 31242
rect 17677 31184 17682 31240
rect 17738 31184 19154 31240
rect 19210 31184 19215 31240
rect 17677 31182 19215 31184
rect 17677 31179 17743 31182
rect 19149 31179 19215 31182
rect 21357 31242 21423 31245
rect 42149 31242 42215 31245
rect 21357 31240 42215 31242
rect 21357 31184 21362 31240
rect 21418 31184 42154 31240
rect 42210 31184 42215 31240
rect 21357 31182 42215 31184
rect 21357 31179 21423 31182
rect 42149 31179 42215 31182
rect 18597 31106 18663 31109
rect 23657 31106 23723 31109
rect 24577 31106 24643 31109
rect 18597 31104 24643 31106
rect 18597 31048 18602 31104
rect 18658 31048 23662 31104
rect 23718 31048 24582 31104
rect 24638 31048 24643 31104
rect 18597 31046 24643 31048
rect 18597 31043 18663 31046
rect 23657 31043 23723 31046
rect 24577 31043 24643 31046
rect 24761 31106 24827 31109
rect 25446 31106 25452 31108
rect 24761 31104 25452 31106
rect 24761 31048 24766 31104
rect 24822 31048 25452 31104
rect 24761 31046 25452 31048
rect 24761 31043 24827 31046
rect 25446 31044 25452 31046
rect 25516 31044 25522 31108
rect 25814 31044 25820 31108
rect 25884 31106 25890 31108
rect 25957 31106 26023 31109
rect 27337 31106 27403 31109
rect 25884 31104 26023 31106
rect 25884 31048 25962 31104
rect 26018 31048 26023 31104
rect 25884 31046 26023 31048
rect 25884 31044 25890 31046
rect 25957 31043 26023 31046
rect 26190 31104 27403 31106
rect 26190 31048 27342 31104
rect 27398 31048 27403 31104
rect 26190 31046 27403 31048
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 15469 30970 15535 30973
rect 17401 30970 17467 30973
rect 18505 30970 18571 30973
rect 22369 30970 22435 30973
rect 24945 30970 25011 30973
rect 15469 30968 21098 30970
rect 15469 30912 15474 30968
rect 15530 30912 17406 30968
rect 17462 30912 18510 30968
rect 18566 30912 21098 30968
rect 15469 30910 21098 30912
rect 15469 30907 15535 30910
rect 17401 30907 17467 30910
rect 18505 30907 18571 30910
rect 19517 30834 19583 30837
rect 20713 30834 20779 30837
rect 21038 30836 21098 30910
rect 22369 30968 25011 30970
rect 22369 30912 22374 30968
rect 22430 30912 24950 30968
rect 25006 30912 25011 30968
rect 22369 30910 25011 30912
rect 22369 30907 22435 30910
rect 24945 30907 25011 30910
rect 25865 30970 25931 30973
rect 26190 30972 26250 31046
rect 27337 31043 27403 31046
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 26182 30970 26188 30972
rect 25865 30968 26188 30970
rect 25865 30912 25870 30968
rect 25926 30912 26188 30968
rect 25865 30910 26188 30912
rect 25865 30907 25931 30910
rect 26182 30908 26188 30910
rect 26252 30908 26258 30972
rect 26325 30970 26391 30973
rect 28165 30970 28231 30973
rect 26325 30968 28231 30970
rect 26325 30912 26330 30968
rect 26386 30912 28170 30968
rect 28226 30912 28231 30968
rect 26325 30910 28231 30912
rect 26325 30907 26391 30910
rect 28165 30907 28231 30910
rect 19517 30832 20779 30834
rect 19517 30776 19522 30832
rect 19578 30776 20718 30832
rect 20774 30776 20779 30832
rect 19517 30774 20779 30776
rect 19517 30771 19583 30774
rect 20713 30771 20779 30774
rect 21030 30772 21036 30836
rect 21100 30772 21106 30836
rect 24301 30834 24367 30837
rect 28717 30834 28783 30837
rect 24301 30832 28783 30834
rect 24301 30776 24306 30832
rect 24362 30776 28722 30832
rect 28778 30776 28783 30832
rect 24301 30774 28783 30776
rect 24301 30771 24367 30774
rect 28717 30771 28783 30774
rect 3325 30698 3391 30701
rect 4889 30698 4955 30701
rect 3325 30696 4955 30698
rect 3325 30640 3330 30696
rect 3386 30640 4894 30696
rect 4950 30640 4955 30696
rect 3325 30638 4955 30640
rect 3325 30635 3391 30638
rect 4889 30635 4955 30638
rect 17309 30698 17375 30701
rect 22645 30698 22711 30701
rect 17309 30696 22711 30698
rect 17309 30640 17314 30696
rect 17370 30640 22650 30696
rect 22706 30640 22711 30696
rect 17309 30638 22711 30640
rect 17309 30635 17375 30638
rect 22645 30635 22711 30638
rect 22921 30698 22987 30701
rect 23841 30698 23907 30701
rect 31661 30698 31727 30701
rect 22921 30696 31727 30698
rect 22921 30640 22926 30696
rect 22982 30640 23846 30696
rect 23902 30640 31666 30696
rect 31722 30640 31727 30696
rect 22921 30638 31727 30640
rect 22921 30635 22987 30638
rect 23841 30635 23907 30638
rect 31661 30635 31727 30638
rect 0 30562 800 30592
rect 1209 30562 1275 30565
rect 0 30560 1275 30562
rect 0 30504 1214 30560
rect 1270 30504 1275 30560
rect 0 30502 1275 30504
rect 0 30472 800 30502
rect 1209 30499 1275 30502
rect 2865 30562 2931 30565
rect 5441 30562 5507 30565
rect 2865 30560 5507 30562
rect 2865 30504 2870 30560
rect 2926 30504 5446 30560
rect 5502 30504 5507 30560
rect 2865 30502 5507 30504
rect 2865 30499 2931 30502
rect 5441 30499 5507 30502
rect 9622 30500 9628 30564
rect 9692 30562 9698 30564
rect 14641 30562 14707 30565
rect 9692 30560 14707 30562
rect 9692 30504 14646 30560
rect 14702 30504 14707 30560
rect 9692 30502 14707 30504
rect 9692 30500 9698 30502
rect 14641 30499 14707 30502
rect 16430 30500 16436 30564
rect 16500 30562 16506 30564
rect 18321 30562 18387 30565
rect 16500 30560 18387 30562
rect 16500 30504 18326 30560
rect 18382 30504 18387 30560
rect 16500 30502 18387 30504
rect 16500 30500 16506 30502
rect 18321 30499 18387 30502
rect 20161 30562 20227 30565
rect 20529 30562 20595 30565
rect 21817 30562 21883 30565
rect 25773 30562 25839 30565
rect 20161 30560 21883 30562
rect 20161 30504 20166 30560
rect 20222 30504 20534 30560
rect 20590 30504 21822 30560
rect 21878 30504 21883 30560
rect 20161 30502 21883 30504
rect 20161 30499 20227 30502
rect 20529 30499 20595 30502
rect 21817 30499 21883 30502
rect 23108 30560 25839 30562
rect 23108 30504 25778 30560
rect 25834 30504 25839 30560
rect 23108 30502 25839 30504
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 23108 30429 23168 30502
rect 25773 30499 25839 30502
rect 26550 30500 26556 30564
rect 26620 30562 26626 30564
rect 27705 30562 27771 30565
rect 26620 30560 27771 30562
rect 26620 30504 27710 30560
rect 27766 30504 27771 30560
rect 26620 30502 27771 30504
rect 26620 30500 26626 30502
rect 27705 30499 27771 30502
rect 2957 30426 3023 30429
rect 4797 30426 4863 30429
rect 5165 30428 5231 30429
rect 5165 30426 5212 30428
rect 2957 30424 4863 30426
rect 2957 30368 2962 30424
rect 3018 30368 4802 30424
rect 4858 30368 4863 30424
rect 2957 30366 4863 30368
rect 5120 30424 5212 30426
rect 5120 30368 5170 30424
rect 5120 30366 5212 30368
rect 2957 30363 3023 30366
rect 4797 30363 4863 30366
rect 5165 30364 5212 30366
rect 5276 30364 5282 30428
rect 10041 30426 10107 30429
rect 10910 30426 10916 30428
rect 10041 30424 10916 30426
rect 10041 30368 10046 30424
rect 10102 30368 10916 30424
rect 10041 30366 10916 30368
rect 5165 30363 5231 30364
rect 10041 30363 10107 30366
rect 10910 30364 10916 30366
rect 10980 30364 10986 30428
rect 14457 30426 14523 30429
rect 14590 30426 14596 30428
rect 14457 30424 14596 30426
rect 14457 30368 14462 30424
rect 14518 30368 14596 30424
rect 14457 30366 14596 30368
rect 14457 30363 14523 30366
rect 14590 30364 14596 30366
rect 14660 30364 14666 30428
rect 14958 30364 14964 30428
rect 15028 30426 15034 30428
rect 17953 30426 18019 30429
rect 15028 30424 18019 30426
rect 15028 30368 17958 30424
rect 18014 30368 18019 30424
rect 15028 30366 18019 30368
rect 15028 30364 15034 30366
rect 17953 30363 18019 30366
rect 21265 30426 21331 30429
rect 23105 30426 23171 30429
rect 21265 30424 23171 30426
rect 21265 30368 21270 30424
rect 21326 30368 23110 30424
rect 23166 30368 23171 30424
rect 21265 30366 23171 30368
rect 21265 30363 21331 30366
rect 23105 30363 23171 30366
rect 26366 30364 26372 30428
rect 26436 30426 26442 30428
rect 26969 30426 27035 30429
rect 26436 30424 27035 30426
rect 26436 30368 26974 30424
rect 27030 30368 27035 30424
rect 26436 30366 27035 30368
rect 26436 30364 26442 30366
rect 26969 30363 27035 30366
rect 4521 30290 4587 30293
rect 4981 30290 5047 30293
rect 4521 30288 5047 30290
rect 4521 30232 4526 30288
rect 4582 30232 4986 30288
rect 5042 30232 5047 30288
rect 4521 30230 5047 30232
rect 4521 30227 4587 30230
rect 4981 30227 5047 30230
rect 6453 30290 6519 30293
rect 8753 30290 8819 30293
rect 11329 30290 11395 30293
rect 15469 30290 15535 30293
rect 6453 30288 15535 30290
rect 6453 30232 6458 30288
rect 6514 30232 8758 30288
rect 8814 30232 11334 30288
rect 11390 30232 15474 30288
rect 15530 30232 15535 30288
rect 6453 30230 15535 30232
rect 6453 30227 6519 30230
rect 8753 30227 8819 30230
rect 11329 30227 11395 30230
rect 15469 30227 15535 30230
rect 15929 30290 15995 30293
rect 17953 30290 18019 30293
rect 15929 30288 18019 30290
rect 15929 30232 15934 30288
rect 15990 30232 17958 30288
rect 18014 30232 18019 30288
rect 15929 30230 18019 30232
rect 15929 30227 15995 30230
rect 17953 30227 18019 30230
rect 19149 30290 19215 30293
rect 20437 30290 20503 30293
rect 19149 30288 20503 30290
rect 19149 30232 19154 30288
rect 19210 30232 20442 30288
rect 20498 30232 20503 30288
rect 19149 30230 20503 30232
rect 19149 30227 19215 30230
rect 20437 30227 20503 30230
rect 20805 30290 20871 30293
rect 24669 30290 24735 30293
rect 20805 30288 24735 30290
rect 20805 30232 20810 30288
rect 20866 30232 24674 30288
rect 24730 30232 24735 30288
rect 20805 30230 24735 30232
rect 20805 30227 20871 30230
rect 24669 30227 24735 30230
rect 25313 30290 25379 30293
rect 25865 30290 25931 30293
rect 26509 30290 26575 30293
rect 25313 30288 26575 30290
rect 25313 30232 25318 30288
rect 25374 30232 25870 30288
rect 25926 30232 26514 30288
rect 26570 30232 26575 30288
rect 25313 30230 26575 30232
rect 25313 30227 25379 30230
rect 25865 30227 25931 30230
rect 26509 30227 26575 30230
rect 16481 30154 16547 30157
rect 21357 30154 21423 30157
rect 16481 30152 21423 30154
rect 16481 30096 16486 30152
rect 16542 30096 21362 30152
rect 21418 30096 21423 30152
rect 16481 30094 21423 30096
rect 16481 30091 16547 30094
rect 21357 30091 21423 30094
rect 21541 30154 21607 30157
rect 22921 30154 22987 30157
rect 25262 30154 25268 30156
rect 21541 30152 25268 30154
rect 21541 30096 21546 30152
rect 21602 30096 22926 30152
rect 22982 30096 25268 30152
rect 21541 30094 25268 30096
rect 21541 30091 21607 30094
rect 22921 30091 22987 30094
rect 25262 30092 25268 30094
rect 25332 30154 25338 30156
rect 25405 30154 25471 30157
rect 25332 30152 25471 30154
rect 25332 30096 25410 30152
rect 25466 30096 25471 30152
rect 25332 30094 25471 30096
rect 25332 30092 25338 30094
rect 25405 30091 25471 30094
rect 25773 30154 25839 30157
rect 28717 30154 28783 30157
rect 25773 30152 28783 30154
rect 25773 30096 25778 30152
rect 25834 30096 28722 30152
rect 28778 30096 28783 30152
rect 25773 30094 28783 30096
rect 25773 30091 25839 30094
rect 28717 30091 28783 30094
rect 14273 30018 14339 30021
rect 19149 30018 19215 30021
rect 14273 30016 19215 30018
rect 14273 29960 14278 30016
rect 14334 29960 19154 30016
rect 19210 29960 19215 30016
rect 14273 29958 19215 29960
rect 14273 29955 14339 29958
rect 19149 29955 19215 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 11881 29882 11947 29885
rect 12985 29882 13051 29885
rect 11881 29880 13051 29882
rect 11881 29824 11886 29880
rect 11942 29824 12990 29880
rect 13046 29824 13051 29880
rect 11881 29822 13051 29824
rect 11881 29819 11947 29822
rect 12985 29819 13051 29822
rect 17861 29882 17927 29885
rect 21544 29882 21604 30091
rect 24117 30018 24183 30021
rect 29085 30018 29151 30021
rect 24117 30016 29151 30018
rect 24117 29960 24122 30016
rect 24178 29960 29090 30016
rect 29146 29960 29151 30016
rect 24117 29958 29151 29960
rect 24117 29955 24183 29958
rect 29085 29955 29151 29958
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 17861 29880 21604 29882
rect 17861 29824 17866 29880
rect 17922 29824 21604 29880
rect 17861 29822 21604 29824
rect 23197 29882 23263 29885
rect 25221 29882 25287 29885
rect 23197 29880 25287 29882
rect 23197 29824 23202 29880
rect 23258 29824 25226 29880
rect 25282 29824 25287 29880
rect 23197 29822 25287 29824
rect 17861 29819 17927 29822
rect 23197 29819 23263 29822
rect 25221 29819 25287 29822
rect 27061 29882 27127 29885
rect 29361 29882 29427 29885
rect 27061 29880 29427 29882
rect 27061 29824 27066 29880
rect 27122 29824 29366 29880
rect 29422 29824 29427 29880
rect 27061 29822 29427 29824
rect 27061 29819 27127 29822
rect 29361 29819 29427 29822
rect 4061 29746 4127 29749
rect 5349 29746 5415 29749
rect 4061 29744 5415 29746
rect 4061 29688 4066 29744
rect 4122 29688 5354 29744
rect 5410 29688 5415 29744
rect 4061 29686 5415 29688
rect 4061 29683 4127 29686
rect 5349 29683 5415 29686
rect 10225 29746 10291 29749
rect 11881 29746 11947 29749
rect 13537 29746 13603 29749
rect 10225 29744 13603 29746
rect 10225 29688 10230 29744
rect 10286 29688 11886 29744
rect 11942 29688 13542 29744
rect 13598 29688 13603 29744
rect 10225 29686 13603 29688
rect 10225 29683 10291 29686
rect 11881 29683 11947 29686
rect 13537 29683 13603 29686
rect 14457 29746 14523 29749
rect 15469 29746 15535 29749
rect 14457 29744 15535 29746
rect 14457 29688 14462 29744
rect 14518 29688 15474 29744
rect 15530 29688 15535 29744
rect 14457 29686 15535 29688
rect 14457 29683 14523 29686
rect 15469 29683 15535 29686
rect 16113 29746 16179 29749
rect 21725 29746 21791 29749
rect 16113 29744 21791 29746
rect 16113 29688 16118 29744
rect 16174 29688 21730 29744
rect 21786 29688 21791 29744
rect 16113 29686 21791 29688
rect 16113 29683 16179 29686
rect 21725 29683 21791 29686
rect 30189 29746 30255 29749
rect 30557 29746 30623 29749
rect 30189 29744 30623 29746
rect 30189 29688 30194 29744
rect 30250 29688 30562 29744
rect 30618 29688 30623 29744
rect 30189 29686 30623 29688
rect 30189 29683 30255 29686
rect 30557 29683 30623 29686
rect 7833 29610 7899 29613
rect 13169 29610 13235 29613
rect 7833 29608 13235 29610
rect 7833 29552 7838 29608
rect 7894 29552 13174 29608
rect 13230 29552 13235 29608
rect 7833 29550 13235 29552
rect 7833 29547 7899 29550
rect 13169 29547 13235 29550
rect 13721 29610 13787 29613
rect 18137 29610 18203 29613
rect 20345 29610 20411 29613
rect 23105 29610 23171 29613
rect 13721 29608 20224 29610
rect 13721 29552 13726 29608
rect 13782 29552 18142 29608
rect 18198 29552 20224 29608
rect 13721 29550 20224 29552
rect 13721 29547 13787 29550
rect 18137 29547 18203 29550
rect 0 29474 800 29504
rect 20164 29477 20224 29550
rect 20345 29608 23171 29610
rect 20345 29552 20350 29608
rect 20406 29552 23110 29608
rect 23166 29552 23171 29608
rect 20345 29550 23171 29552
rect 20345 29547 20411 29550
rect 23105 29547 23171 29550
rect 23565 29610 23631 29613
rect 31937 29610 32003 29613
rect 23565 29608 32003 29610
rect 23565 29552 23570 29608
rect 23626 29552 31942 29608
rect 31998 29552 32003 29608
rect 23565 29550 32003 29552
rect 23565 29547 23631 29550
rect 31937 29547 32003 29550
rect 1209 29474 1275 29477
rect 0 29472 1275 29474
rect 0 29416 1214 29472
rect 1270 29416 1275 29472
rect 0 29414 1275 29416
rect 0 29384 800 29414
rect 1209 29411 1275 29414
rect 3049 29474 3115 29477
rect 7281 29474 7347 29477
rect 3049 29472 7347 29474
rect 3049 29416 3054 29472
rect 3110 29416 7286 29472
rect 7342 29416 7347 29472
rect 3049 29414 7347 29416
rect 3049 29411 3115 29414
rect 7281 29411 7347 29414
rect 11973 29474 12039 29477
rect 12709 29474 12775 29477
rect 11973 29472 12775 29474
rect 11973 29416 11978 29472
rect 12034 29416 12714 29472
rect 12770 29416 12775 29472
rect 11973 29414 12775 29416
rect 11973 29411 12039 29414
rect 12709 29411 12775 29414
rect 16297 29474 16363 29477
rect 18597 29474 18663 29477
rect 20161 29474 20227 29477
rect 21173 29474 21239 29477
rect 16297 29472 18663 29474
rect 16297 29416 16302 29472
rect 16358 29416 18602 29472
rect 18658 29416 18663 29472
rect 16297 29414 18663 29416
rect 20070 29472 21239 29474
rect 20070 29416 20166 29472
rect 20222 29416 21178 29472
rect 21234 29416 21239 29472
rect 20070 29414 21239 29416
rect 16297 29411 16363 29414
rect 18597 29411 18663 29414
rect 20161 29411 20227 29414
rect 21173 29411 21239 29414
rect 21449 29474 21515 29477
rect 24945 29474 25011 29477
rect 27337 29474 27403 29477
rect 28809 29474 28875 29477
rect 21449 29472 28875 29474
rect 21449 29416 21454 29472
rect 21510 29416 24950 29472
rect 25006 29416 27342 29472
rect 27398 29416 28814 29472
rect 28870 29416 28875 29472
rect 21449 29414 28875 29416
rect 21449 29411 21515 29414
rect 24945 29411 25011 29414
rect 27337 29411 27403 29414
rect 28809 29411 28875 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 2313 29338 2379 29341
rect 3325 29338 3391 29341
rect 2313 29336 3391 29338
rect 2313 29280 2318 29336
rect 2374 29280 3330 29336
rect 3386 29280 3391 29336
rect 2313 29278 3391 29280
rect 2313 29275 2379 29278
rect 3325 29275 3391 29278
rect 9857 29338 9923 29341
rect 17033 29338 17099 29341
rect 9857 29336 17099 29338
rect 9857 29280 9862 29336
rect 9918 29280 17038 29336
rect 17094 29280 17099 29336
rect 9857 29278 17099 29280
rect 9857 29275 9923 29278
rect 17033 29275 17099 29278
rect 21449 29338 21515 29341
rect 22093 29338 22159 29341
rect 23841 29338 23907 29341
rect 21449 29336 23907 29338
rect 21449 29280 21454 29336
rect 21510 29280 22098 29336
rect 22154 29280 23846 29336
rect 23902 29280 23907 29336
rect 21449 29278 23907 29280
rect 21449 29275 21515 29278
rect 22093 29275 22159 29278
rect 23841 29275 23907 29278
rect 28533 29338 28599 29341
rect 29269 29338 29335 29341
rect 28533 29336 29335 29338
rect 28533 29280 28538 29336
rect 28594 29280 29274 29336
rect 29330 29280 29335 29336
rect 28533 29278 29335 29280
rect 28533 29275 28599 29278
rect 29269 29275 29335 29278
rect 1485 29202 1551 29205
rect 4521 29202 4587 29205
rect 1485 29200 4587 29202
rect 1485 29144 1490 29200
rect 1546 29144 4526 29200
rect 4582 29144 4587 29200
rect 1485 29142 4587 29144
rect 1485 29139 1551 29142
rect 4521 29139 4587 29142
rect 4981 29200 5047 29205
rect 4981 29144 4986 29200
rect 5042 29144 5047 29200
rect 4981 29139 5047 29144
rect 9121 29202 9187 29205
rect 9489 29202 9555 29205
rect 10869 29202 10935 29205
rect 9121 29200 10935 29202
rect 9121 29144 9126 29200
rect 9182 29144 9494 29200
rect 9550 29144 10874 29200
rect 10930 29144 10935 29200
rect 9121 29142 10935 29144
rect 9121 29139 9187 29142
rect 9489 29139 9555 29142
rect 10869 29139 10935 29142
rect 11053 29202 11119 29205
rect 13077 29202 13143 29205
rect 11053 29200 13143 29202
rect 11053 29144 11058 29200
rect 11114 29144 13082 29200
rect 13138 29144 13143 29200
rect 11053 29142 13143 29144
rect 11053 29139 11119 29142
rect 13077 29139 13143 29142
rect 17902 29140 17908 29204
rect 17972 29202 17978 29204
rect 22553 29202 22619 29205
rect 25037 29202 25103 29205
rect 17972 29200 25103 29202
rect 17972 29144 22558 29200
rect 22614 29144 25042 29200
rect 25098 29144 25103 29200
rect 17972 29142 25103 29144
rect 17972 29140 17978 29142
rect 22553 29139 22619 29142
rect 25037 29139 25103 29142
rect 27337 29202 27403 29205
rect 29453 29202 29519 29205
rect 27337 29200 29519 29202
rect 27337 29144 27342 29200
rect 27398 29144 29458 29200
rect 29514 29144 29519 29200
rect 27337 29142 29519 29144
rect 27337 29139 27403 29142
rect 29453 29139 29519 29142
rect 4984 29066 5044 29139
rect 13169 29066 13235 29069
rect 20437 29066 20503 29069
rect 4984 29064 20503 29066
rect 4984 29008 13174 29064
rect 13230 29008 20442 29064
rect 20498 29008 20503 29064
rect 4984 29006 20503 29008
rect 13169 29003 13235 29006
rect 20437 29003 20503 29006
rect 22921 29066 22987 29069
rect 23238 29066 23244 29068
rect 22921 29064 23244 29066
rect 22921 29008 22926 29064
rect 22982 29008 23244 29064
rect 22921 29006 23244 29008
rect 22921 29003 22987 29006
rect 23238 29004 23244 29006
rect 23308 29004 23314 29068
rect 24669 29066 24735 29069
rect 29545 29066 29611 29069
rect 30097 29066 30163 29069
rect 24669 29064 30163 29066
rect 24669 29008 24674 29064
rect 24730 29008 29550 29064
rect 29606 29008 30102 29064
rect 30158 29008 30163 29064
rect 24669 29006 30163 29008
rect 24669 29003 24735 29006
rect 29545 29003 29611 29006
rect 30097 29003 30163 29006
rect 9254 28868 9260 28932
rect 9324 28930 9330 28932
rect 9622 28930 9628 28932
rect 9324 28870 9628 28930
rect 9324 28868 9330 28870
rect 9622 28868 9628 28870
rect 9692 28868 9698 28932
rect 15101 28930 15167 28933
rect 22645 28930 22711 28933
rect 26550 28930 26556 28932
rect 15101 28928 22711 28930
rect 15101 28872 15106 28928
rect 15162 28872 22650 28928
rect 22706 28872 22711 28928
rect 15101 28870 22711 28872
rect 15101 28867 15167 28870
rect 22645 28867 22711 28870
rect 24534 28870 26556 28930
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 2221 28794 2287 28797
rect 3969 28794 4035 28797
rect 2221 28792 4035 28794
rect 2221 28736 2226 28792
rect 2282 28736 3974 28792
rect 4030 28736 4035 28792
rect 2221 28734 4035 28736
rect 2221 28731 2287 28734
rect 3969 28731 4035 28734
rect 4797 28794 4863 28797
rect 5625 28794 5691 28797
rect 4797 28792 5691 28794
rect 4797 28736 4802 28792
rect 4858 28736 5630 28792
rect 5686 28736 5691 28792
rect 4797 28734 5691 28736
rect 4797 28731 4863 28734
rect 5625 28731 5691 28734
rect 6361 28794 6427 28797
rect 8150 28794 8156 28796
rect 6361 28792 8156 28794
rect 6361 28736 6366 28792
rect 6422 28736 8156 28792
rect 6361 28734 8156 28736
rect 6361 28731 6427 28734
rect 8150 28732 8156 28734
rect 8220 28732 8226 28796
rect 16246 28732 16252 28796
rect 16316 28794 16322 28796
rect 24534 28794 24594 28870
rect 26550 28868 26556 28870
rect 26620 28868 26626 28932
rect 27705 28930 27771 28933
rect 28625 28930 28691 28933
rect 27705 28928 28691 28930
rect 27705 28872 27710 28928
rect 27766 28872 28630 28928
rect 28686 28872 28691 28928
rect 27705 28870 28691 28872
rect 27705 28867 27771 28870
rect 28625 28867 28691 28870
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 16316 28734 24594 28794
rect 24669 28794 24735 28797
rect 24894 28794 24900 28796
rect 24669 28792 24900 28794
rect 24669 28736 24674 28792
rect 24730 28736 24900 28792
rect 24669 28734 24900 28736
rect 16316 28732 16322 28734
rect 24669 28731 24735 28734
rect 24894 28732 24900 28734
rect 24964 28732 24970 28796
rect 26417 28794 26483 28797
rect 27797 28794 27863 28797
rect 26417 28792 27863 28794
rect 26417 28736 26422 28792
rect 26478 28736 27802 28792
rect 27858 28736 27863 28792
rect 26417 28734 27863 28736
rect 26417 28731 26483 28734
rect 27797 28731 27863 28734
rect 3601 28658 3667 28661
rect 4800 28658 4860 28731
rect 3601 28656 4860 28658
rect 3601 28600 3606 28656
rect 3662 28600 4860 28656
rect 3601 28598 4860 28600
rect 18597 28658 18663 28661
rect 19885 28658 19951 28661
rect 18597 28656 19951 28658
rect 18597 28600 18602 28656
rect 18658 28600 19890 28656
rect 19946 28600 19951 28656
rect 18597 28598 19951 28600
rect 3601 28595 3667 28598
rect 18597 28595 18663 28598
rect 19885 28595 19951 28598
rect 20161 28658 20227 28661
rect 31477 28658 31543 28661
rect 20161 28656 31543 28658
rect 20161 28600 20166 28656
rect 20222 28600 31482 28656
rect 31538 28600 31543 28656
rect 20161 28598 31543 28600
rect 20161 28595 20227 28598
rect 31477 28595 31543 28598
rect 4429 28522 4495 28525
rect 6361 28522 6427 28525
rect 4429 28520 6427 28522
rect 4429 28464 4434 28520
rect 4490 28464 6366 28520
rect 6422 28464 6427 28520
rect 4429 28462 6427 28464
rect 4429 28459 4495 28462
rect 6361 28459 6427 28462
rect 19333 28522 19399 28525
rect 19793 28522 19859 28525
rect 31385 28522 31451 28525
rect 19333 28520 31451 28522
rect 19333 28464 19338 28520
rect 19394 28464 19798 28520
rect 19854 28464 31390 28520
rect 31446 28464 31451 28520
rect 19333 28462 31451 28464
rect 19333 28459 19399 28462
rect 19793 28459 19859 28462
rect 31385 28459 31451 28462
rect 0 28386 800 28416
rect 1209 28386 1275 28389
rect 0 28384 1275 28386
rect 0 28328 1214 28384
rect 1270 28328 1275 28384
rect 0 28326 1275 28328
rect 0 28296 800 28326
rect 1209 28323 1275 28326
rect 3233 28386 3299 28389
rect 5625 28386 5691 28389
rect 27705 28388 27771 28389
rect 3233 28384 5691 28386
rect 3233 28328 3238 28384
rect 3294 28328 5630 28384
rect 5686 28328 5691 28384
rect 3233 28326 5691 28328
rect 3233 28323 3299 28326
rect 5625 28323 5691 28326
rect 27654 28324 27660 28388
rect 27724 28386 27771 28388
rect 27724 28384 27816 28386
rect 27766 28328 27816 28384
rect 27724 28326 27816 28328
rect 27724 28324 27771 28326
rect 27705 28323 27771 28324
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 3969 28250 4035 28253
rect 18137 28250 18203 28253
rect 3969 28248 18203 28250
rect 3969 28192 3974 28248
rect 4030 28192 18142 28248
rect 18198 28192 18203 28248
rect 3969 28190 18203 28192
rect 3969 28187 4035 28190
rect 18137 28187 18203 28190
rect 1577 28114 1643 28117
rect 7046 28114 7052 28116
rect 1577 28112 7052 28114
rect 1577 28056 1582 28112
rect 1638 28056 7052 28112
rect 1577 28054 7052 28056
rect 1577 28051 1643 28054
rect 7046 28052 7052 28054
rect 7116 28052 7122 28116
rect 14181 28114 14247 28117
rect 8250 28112 14247 28114
rect 8250 28056 14186 28112
rect 14242 28056 14247 28112
rect 8250 28054 14247 28056
rect 2957 27978 3023 27981
rect 5574 27978 5580 27980
rect 2957 27976 5580 27978
rect 2957 27920 2962 27976
rect 3018 27920 5580 27976
rect 2957 27918 5580 27920
rect 2957 27915 3023 27918
rect 5574 27916 5580 27918
rect 5644 27916 5650 27980
rect 6637 27978 6703 27981
rect 8250 27978 8310 28054
rect 14181 28051 14247 28054
rect 16481 28114 16547 28117
rect 20805 28114 20871 28117
rect 16481 28112 20871 28114
rect 16481 28056 16486 28112
rect 16542 28056 20810 28112
rect 20866 28056 20871 28112
rect 16481 28054 20871 28056
rect 16481 28051 16547 28054
rect 20805 28051 20871 28054
rect 43805 28114 43871 28117
rect 44200 28114 45000 28144
rect 43805 28112 45000 28114
rect 43805 28056 43810 28112
rect 43866 28056 45000 28112
rect 43805 28054 45000 28056
rect 43805 28051 43871 28054
rect 44200 28024 45000 28054
rect 6637 27976 8310 27978
rect 6637 27920 6642 27976
rect 6698 27920 8310 27976
rect 6637 27918 8310 27920
rect 6637 27915 6703 27918
rect 16614 27916 16620 27980
rect 16684 27978 16690 27980
rect 16757 27978 16823 27981
rect 16684 27976 16823 27978
rect 16684 27920 16762 27976
rect 16818 27920 16823 27976
rect 16684 27918 16823 27920
rect 16684 27916 16690 27918
rect 16757 27915 16823 27918
rect 17309 27978 17375 27981
rect 25313 27978 25379 27981
rect 17309 27976 25379 27978
rect 17309 27920 17314 27976
rect 17370 27920 25318 27976
rect 25374 27920 25379 27976
rect 17309 27918 25379 27920
rect 17309 27915 17375 27918
rect 25313 27915 25379 27918
rect 5533 27842 5599 27845
rect 7005 27842 7071 27845
rect 5533 27840 7071 27842
rect 5533 27784 5538 27840
rect 5594 27784 7010 27840
rect 7066 27784 7071 27840
rect 5533 27782 7071 27784
rect 5533 27779 5599 27782
rect 7005 27779 7071 27782
rect 7598 27780 7604 27844
rect 7668 27842 7674 27844
rect 9029 27842 9095 27845
rect 14365 27842 14431 27845
rect 7668 27840 14431 27842
rect 7668 27784 9034 27840
rect 9090 27784 14370 27840
rect 14426 27784 14431 27840
rect 7668 27782 14431 27784
rect 7668 27780 7674 27782
rect 9029 27779 9095 27782
rect 14365 27779 14431 27782
rect 18229 27842 18295 27845
rect 18597 27842 18663 27845
rect 18229 27840 18663 27842
rect 18229 27784 18234 27840
rect 18290 27784 18602 27840
rect 18658 27784 18663 27840
rect 18229 27782 18663 27784
rect 18229 27779 18295 27782
rect 18597 27779 18663 27782
rect 19149 27842 19215 27845
rect 21265 27842 21331 27845
rect 19149 27840 21331 27842
rect 19149 27784 19154 27840
rect 19210 27784 21270 27840
rect 21326 27784 21331 27840
rect 19149 27782 21331 27784
rect 19149 27779 19215 27782
rect 21265 27779 21331 27782
rect 26785 27842 26851 27845
rect 28165 27842 28231 27845
rect 26785 27840 28231 27842
rect 26785 27784 26790 27840
rect 26846 27784 28170 27840
rect 28226 27784 28231 27840
rect 26785 27782 28231 27784
rect 26785 27779 26851 27782
rect 28165 27779 28231 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 8293 27706 8359 27709
rect 9581 27706 9647 27709
rect 8293 27704 9647 27706
rect 8293 27648 8298 27704
rect 8354 27648 9586 27704
rect 9642 27648 9647 27704
rect 8293 27646 9647 27648
rect 8293 27643 8359 27646
rect 9581 27643 9647 27646
rect 11053 27706 11119 27709
rect 13077 27706 13143 27709
rect 13813 27706 13879 27709
rect 25865 27706 25931 27709
rect 27245 27706 27311 27709
rect 11053 27704 13879 27706
rect 11053 27648 11058 27704
rect 11114 27648 13082 27704
rect 13138 27648 13818 27704
rect 13874 27648 13879 27704
rect 11053 27646 13879 27648
rect 11053 27643 11119 27646
rect 13077 27643 13143 27646
rect 13813 27643 13879 27646
rect 17542 27646 20316 27706
rect 13537 27570 13603 27573
rect 9630 27568 13603 27570
rect 9630 27512 13542 27568
rect 13598 27512 13603 27568
rect 9630 27510 13603 27512
rect 6361 27434 6427 27437
rect 6729 27434 6795 27437
rect 8293 27434 8359 27437
rect 9630 27434 9690 27510
rect 13537 27507 13603 27510
rect 16757 27570 16823 27573
rect 17542 27570 17602 27646
rect 16757 27568 17602 27570
rect 16757 27512 16762 27568
rect 16818 27512 17602 27568
rect 16757 27510 17602 27512
rect 17769 27570 17835 27573
rect 17902 27570 17908 27572
rect 17769 27568 17908 27570
rect 17769 27512 17774 27568
rect 17830 27512 17908 27568
rect 17769 27510 17908 27512
rect 16757 27507 16823 27510
rect 17769 27507 17835 27510
rect 17902 27508 17908 27510
rect 17972 27508 17978 27572
rect 20256 27570 20316 27646
rect 25865 27704 27311 27706
rect 25865 27648 25870 27704
rect 25926 27648 27250 27704
rect 27306 27648 27311 27704
rect 25865 27646 27311 27648
rect 25865 27643 25931 27646
rect 27245 27643 27311 27646
rect 23289 27570 23355 27573
rect 19244 27510 20178 27570
rect 20256 27568 23355 27570
rect 20256 27512 23294 27568
rect 23350 27512 23355 27568
rect 20256 27510 23355 27512
rect 6361 27432 9690 27434
rect 6361 27376 6366 27432
rect 6422 27376 6734 27432
rect 6790 27376 8298 27432
rect 8354 27376 9690 27432
rect 6361 27374 9690 27376
rect 10409 27434 10475 27437
rect 12617 27434 12683 27437
rect 19244 27434 19304 27510
rect 19793 27434 19859 27437
rect 10409 27432 12683 27434
rect 10409 27376 10414 27432
rect 10470 27376 12622 27432
rect 12678 27376 12683 27432
rect 10409 27374 12683 27376
rect 6361 27371 6427 27374
rect 6729 27371 6795 27374
rect 8293 27371 8359 27374
rect 10409 27371 10475 27374
rect 12617 27371 12683 27374
rect 14598 27374 19304 27434
rect 19382 27432 19859 27434
rect 19382 27376 19798 27432
rect 19854 27376 19859 27432
rect 19382 27374 19859 27376
rect 0 27298 800 27328
rect 1209 27298 1275 27301
rect 0 27296 1275 27298
rect 0 27240 1214 27296
rect 1270 27240 1275 27296
rect 0 27238 1275 27240
rect 0 27208 800 27238
rect 1209 27235 1275 27238
rect 5257 27298 5323 27301
rect 5533 27298 5599 27301
rect 5257 27296 5599 27298
rect 5257 27240 5262 27296
rect 5318 27240 5538 27296
rect 5594 27240 5599 27296
rect 5257 27238 5599 27240
rect 5257 27235 5323 27238
rect 5533 27235 5599 27238
rect 7741 27298 7807 27301
rect 8201 27298 8267 27301
rect 7741 27296 8267 27298
rect 7741 27240 7746 27296
rect 7802 27240 8206 27296
rect 8262 27240 8267 27296
rect 7741 27238 8267 27240
rect 7741 27235 7807 27238
rect 8201 27235 8267 27238
rect 13854 27236 13860 27300
rect 13924 27298 13930 27300
rect 13997 27298 14063 27301
rect 14598 27300 14658 27374
rect 13924 27296 14063 27298
rect 13924 27240 14002 27296
rect 14058 27240 14063 27296
rect 13924 27238 14063 27240
rect 13924 27236 13930 27238
rect 13997 27235 14063 27238
rect 14590 27236 14596 27300
rect 14660 27236 14666 27300
rect 15009 27298 15075 27301
rect 16757 27298 16823 27301
rect 15009 27296 16823 27298
rect 15009 27240 15014 27296
rect 15070 27240 16762 27296
rect 16818 27240 16823 27296
rect 15009 27238 16823 27240
rect 15009 27235 15075 27238
rect 16757 27235 16823 27238
rect 17033 27298 17099 27301
rect 17401 27298 17467 27301
rect 17033 27296 17467 27298
rect 17033 27240 17038 27296
rect 17094 27240 17406 27296
rect 17462 27240 17467 27296
rect 17033 27238 17467 27240
rect 17033 27235 17099 27238
rect 17401 27235 17467 27238
rect 17585 27298 17651 27301
rect 19057 27298 19123 27301
rect 19382 27298 19442 27374
rect 19793 27371 19859 27374
rect 17585 27296 19442 27298
rect 17585 27240 17590 27296
rect 17646 27240 19062 27296
rect 19118 27240 19442 27296
rect 17585 27238 19442 27240
rect 20118 27298 20178 27510
rect 23289 27507 23355 27510
rect 23473 27570 23539 27573
rect 25630 27570 25636 27572
rect 23473 27568 25636 27570
rect 23473 27512 23478 27568
rect 23534 27512 25636 27568
rect 23473 27510 25636 27512
rect 23473 27507 23539 27510
rect 25630 27508 25636 27510
rect 25700 27508 25706 27572
rect 26509 27570 26575 27573
rect 27521 27570 27587 27573
rect 26509 27568 27587 27570
rect 26509 27512 26514 27568
rect 26570 27512 27526 27568
rect 27582 27512 27587 27568
rect 26509 27510 27587 27512
rect 26509 27507 26575 27510
rect 27521 27507 27587 27510
rect 31753 27570 31819 27573
rect 33041 27570 33107 27573
rect 31753 27568 33107 27570
rect 31753 27512 31758 27568
rect 31814 27512 33046 27568
rect 33102 27512 33107 27568
rect 31753 27510 33107 27512
rect 31753 27507 31819 27510
rect 33041 27507 33107 27510
rect 22185 27434 22251 27437
rect 40677 27434 40743 27437
rect 22185 27432 40743 27434
rect 22185 27376 22190 27432
rect 22246 27376 40682 27432
rect 40738 27376 40743 27432
rect 22185 27374 40743 27376
rect 22185 27371 22251 27374
rect 40677 27371 40743 27374
rect 24301 27298 24367 27301
rect 20118 27296 24367 27298
rect 20118 27240 24306 27296
rect 24362 27240 24367 27296
rect 20118 27238 24367 27240
rect 17585 27235 17651 27238
rect 19057 27235 19123 27238
rect 24301 27235 24367 27238
rect 26182 27236 26188 27300
rect 26252 27298 26258 27300
rect 26509 27298 26575 27301
rect 27245 27298 27311 27301
rect 26252 27296 27311 27298
rect 26252 27240 26514 27296
rect 26570 27240 27250 27296
rect 27306 27240 27311 27296
rect 26252 27238 27311 27240
rect 26252 27236 26258 27238
rect 26509 27235 26575 27238
rect 27245 27235 27311 27238
rect 30741 27298 30807 27301
rect 32673 27298 32739 27301
rect 30741 27296 32739 27298
rect 30741 27240 30746 27296
rect 30802 27240 32678 27296
rect 32734 27240 32739 27296
rect 30741 27238 32739 27240
rect 30741 27235 30807 27238
rect 32673 27235 32739 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 1669 27162 1735 27165
rect 7189 27162 7255 27165
rect 8293 27164 8359 27165
rect 8293 27162 8340 27164
rect 1669 27160 7255 27162
rect 1669 27104 1674 27160
rect 1730 27104 7194 27160
rect 7250 27104 7255 27160
rect 1669 27102 7255 27104
rect 8248 27160 8340 27162
rect 8248 27104 8298 27160
rect 8248 27102 8340 27104
rect 1669 27099 1735 27102
rect 7189 27099 7255 27102
rect 8293 27100 8340 27102
rect 8404 27100 8410 27164
rect 10777 27162 10843 27165
rect 15101 27162 15167 27165
rect 10777 27160 15167 27162
rect 10777 27104 10782 27160
rect 10838 27104 15106 27160
rect 15162 27104 15167 27160
rect 10777 27102 15167 27104
rect 8293 27099 8359 27100
rect 10777 27099 10843 27102
rect 15101 27099 15167 27102
rect 16205 27162 16271 27165
rect 22185 27162 22251 27165
rect 16205 27160 19350 27162
rect 16205 27104 16210 27160
rect 16266 27104 19350 27160
rect 16205 27102 19350 27104
rect 16205 27099 16271 27102
rect 4337 27026 4403 27029
rect 4797 27026 4863 27029
rect 7649 27026 7715 27029
rect 4337 27024 7715 27026
rect 4337 26968 4342 27024
rect 4398 26968 4802 27024
rect 4858 26968 7654 27024
rect 7710 26968 7715 27024
rect 4337 26966 7715 26968
rect 4337 26963 4403 26966
rect 4797 26963 4863 26966
rect 7649 26963 7715 26966
rect 11237 27026 11303 27029
rect 11973 27026 12039 27029
rect 16021 27026 16087 27029
rect 18873 27026 18939 27029
rect 11237 27024 18939 27026
rect 11237 26968 11242 27024
rect 11298 26968 11978 27024
rect 12034 26968 16026 27024
rect 16082 26968 18878 27024
rect 18934 26968 18939 27024
rect 11237 26966 18939 26968
rect 19290 27026 19350 27102
rect 20118 27160 22251 27162
rect 20118 27104 22190 27160
rect 22246 27104 22251 27160
rect 20118 27102 22251 27104
rect 20118 27026 20178 27102
rect 22185 27099 22251 27102
rect 23289 27162 23355 27165
rect 26918 27162 26924 27164
rect 23289 27160 26924 27162
rect 23289 27104 23294 27160
rect 23350 27104 26924 27160
rect 23289 27102 26924 27104
rect 23289 27099 23355 27102
rect 26918 27100 26924 27102
rect 26988 27100 26994 27164
rect 31753 27162 31819 27165
rect 31710 27160 31819 27162
rect 31710 27104 31758 27160
rect 31814 27104 31819 27160
rect 31710 27099 31819 27104
rect 19290 26966 20178 27026
rect 22093 27026 22159 27029
rect 30373 27026 30439 27029
rect 31710 27026 31770 27099
rect 22093 27024 31770 27026
rect 22093 26968 22098 27024
rect 22154 26968 30378 27024
rect 30434 26968 31770 27024
rect 22093 26966 31770 26968
rect 11237 26963 11303 26966
rect 11973 26963 12039 26966
rect 16021 26963 16087 26966
rect 18873 26963 18939 26966
rect 22093 26963 22159 26966
rect 30373 26963 30439 26966
rect 4337 26890 4403 26893
rect 5349 26890 5415 26893
rect 4337 26888 5415 26890
rect 4337 26832 4342 26888
rect 4398 26832 5354 26888
rect 5410 26832 5415 26888
rect 4337 26830 5415 26832
rect 4337 26827 4403 26830
rect 5349 26827 5415 26830
rect 5901 26890 5967 26893
rect 6494 26890 6500 26892
rect 5901 26888 6500 26890
rect 5901 26832 5906 26888
rect 5962 26832 6500 26888
rect 5901 26830 6500 26832
rect 5901 26827 5967 26830
rect 6494 26828 6500 26830
rect 6564 26890 6570 26892
rect 9121 26890 9187 26893
rect 6564 26888 9187 26890
rect 6564 26832 9126 26888
rect 9182 26832 9187 26888
rect 6564 26830 9187 26832
rect 6564 26828 6570 26830
rect 9121 26827 9187 26830
rect 17401 26890 17467 26893
rect 23749 26890 23815 26893
rect 17401 26888 23815 26890
rect 17401 26832 17406 26888
rect 17462 26832 23754 26888
rect 23810 26832 23815 26888
rect 17401 26830 23815 26832
rect 17401 26827 17467 26830
rect 23749 26827 23815 26830
rect 26049 26890 26115 26893
rect 28073 26890 28139 26893
rect 26049 26888 28139 26890
rect 26049 26832 26054 26888
rect 26110 26832 28078 26888
rect 28134 26832 28139 26888
rect 26049 26830 28139 26832
rect 26049 26827 26115 26830
rect 28073 26827 28139 26830
rect 4797 26754 4863 26757
rect 5257 26754 5323 26757
rect 4797 26752 5323 26754
rect 4797 26696 4802 26752
rect 4858 26696 5262 26752
rect 5318 26696 5323 26752
rect 4797 26694 5323 26696
rect 4797 26691 4863 26694
rect 5257 26691 5323 26694
rect 13670 26692 13676 26756
rect 13740 26754 13746 26756
rect 19241 26754 19307 26757
rect 13740 26752 19307 26754
rect 13740 26696 19246 26752
rect 19302 26696 19307 26752
rect 13740 26694 19307 26696
rect 13740 26692 13746 26694
rect 19241 26691 19307 26694
rect 19609 26754 19675 26757
rect 20662 26754 20668 26756
rect 19609 26752 20668 26754
rect 19609 26696 19614 26752
rect 19670 26696 20668 26752
rect 19609 26694 20668 26696
rect 19609 26691 19675 26694
rect 20662 26692 20668 26694
rect 20732 26692 20738 26756
rect 22645 26754 22711 26757
rect 28257 26754 28323 26757
rect 22645 26752 28323 26754
rect 22645 26696 22650 26752
rect 22706 26696 28262 26752
rect 28318 26696 28323 26752
rect 22645 26694 28323 26696
rect 22645 26691 22711 26694
rect 28257 26691 28323 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 16389 26620 16455 26621
rect 16389 26618 16436 26620
rect 16344 26616 16436 26618
rect 16344 26560 16394 26616
rect 16344 26558 16436 26560
rect 16389 26556 16436 26558
rect 16500 26556 16506 26620
rect 18321 26618 18387 26621
rect 30097 26618 30163 26621
rect 18321 26616 30163 26618
rect 18321 26560 18326 26616
rect 18382 26560 30102 26616
rect 30158 26560 30163 26616
rect 18321 26558 30163 26560
rect 16389 26555 16455 26556
rect 18321 26555 18387 26558
rect 30097 26555 30163 26558
rect 5165 26482 5231 26485
rect 5809 26482 5875 26485
rect 5165 26480 5875 26482
rect 5165 26424 5170 26480
rect 5226 26424 5814 26480
rect 5870 26424 5875 26480
rect 5165 26422 5875 26424
rect 5165 26419 5231 26422
rect 5809 26419 5875 26422
rect 16021 26482 16087 26485
rect 20529 26482 20595 26485
rect 16021 26480 20595 26482
rect 16021 26424 16026 26480
rect 16082 26424 20534 26480
rect 20590 26424 20595 26480
rect 16021 26422 20595 26424
rect 16021 26419 16087 26422
rect 20529 26419 20595 26422
rect 23197 26482 23263 26485
rect 29269 26482 29335 26485
rect 23197 26480 29335 26482
rect 23197 26424 23202 26480
rect 23258 26424 29274 26480
rect 29330 26424 29335 26480
rect 23197 26422 29335 26424
rect 23197 26419 23263 26422
rect 1577 26346 1643 26349
rect 6729 26346 6795 26349
rect 17309 26348 17375 26349
rect 17309 26346 17356 26348
rect 1577 26344 6795 26346
rect 1577 26288 1582 26344
rect 1638 26288 6734 26344
rect 6790 26288 6795 26344
rect 1577 26286 6795 26288
rect 17264 26344 17356 26346
rect 17264 26288 17314 26344
rect 17264 26286 17356 26288
rect 1577 26283 1643 26286
rect 6729 26283 6795 26286
rect 17309 26284 17356 26286
rect 17420 26284 17426 26348
rect 18045 26346 18111 26349
rect 23381 26346 23447 26349
rect 18045 26344 23447 26346
rect 18045 26288 18050 26344
rect 18106 26288 23386 26344
rect 23442 26288 23447 26344
rect 18045 26286 23447 26288
rect 17309 26283 17375 26284
rect 18045 26283 18111 26286
rect 23381 26283 23447 26286
rect 0 26210 800 26240
rect 1853 26210 1919 26213
rect 0 26208 1919 26210
rect 0 26152 1858 26208
rect 1914 26152 1919 26208
rect 0 26150 1919 26152
rect 0 26120 800 26150
rect 1853 26147 1919 26150
rect 3325 26210 3391 26213
rect 7465 26210 7531 26213
rect 3325 26208 7531 26210
rect 3325 26152 3330 26208
rect 3386 26152 7470 26208
rect 7526 26152 7531 26208
rect 3325 26150 7531 26152
rect 3325 26147 3391 26150
rect 7465 26147 7531 26150
rect 15653 26210 15719 26213
rect 19057 26210 19123 26213
rect 15653 26208 19123 26210
rect 15653 26152 15658 26208
rect 15714 26152 19062 26208
rect 19118 26152 19123 26208
rect 15653 26150 19123 26152
rect 15653 26147 15719 26150
rect 19057 26147 19123 26150
rect 20294 26148 20300 26212
rect 20364 26210 20370 26212
rect 22461 26210 22527 26213
rect 25270 26212 25330 26422
rect 29269 26419 29335 26422
rect 25865 26346 25931 26349
rect 27337 26346 27403 26349
rect 25865 26344 27403 26346
rect 25865 26288 25870 26344
rect 25926 26288 27342 26344
rect 27398 26288 27403 26344
rect 25865 26286 27403 26288
rect 25865 26283 25931 26286
rect 27337 26283 27403 26286
rect 27654 26284 27660 26348
rect 27724 26346 27730 26348
rect 28625 26346 28691 26349
rect 27724 26344 28691 26346
rect 27724 26288 28630 26344
rect 28686 26288 28691 26344
rect 27724 26286 28691 26288
rect 27724 26284 27730 26286
rect 28625 26283 28691 26286
rect 20364 26208 22527 26210
rect 20364 26152 22466 26208
rect 22522 26152 22527 26208
rect 20364 26150 22527 26152
rect 20364 26148 20370 26150
rect 22461 26147 22527 26150
rect 25262 26148 25268 26212
rect 25332 26148 25338 26212
rect 26693 26210 26759 26213
rect 28901 26210 28967 26213
rect 26693 26208 28967 26210
rect 26693 26152 26698 26208
rect 26754 26152 28906 26208
rect 28962 26152 28967 26208
rect 26693 26150 28967 26152
rect 26693 26147 26759 26150
rect 28901 26147 28967 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 6453 26074 6519 26077
rect 7557 26074 7623 26077
rect 6453 26072 7623 26074
rect 6453 26016 6458 26072
rect 6514 26016 7562 26072
rect 7618 26016 7623 26072
rect 6453 26014 7623 26016
rect 6453 26011 6519 26014
rect 7557 26011 7623 26014
rect 8293 26074 8359 26077
rect 9438 26074 9444 26076
rect 8293 26072 9444 26074
rect 8293 26016 8298 26072
rect 8354 26016 9444 26072
rect 8293 26014 9444 26016
rect 8293 26011 8359 26014
rect 9438 26012 9444 26014
rect 9508 26012 9514 26076
rect 11053 26074 11119 26077
rect 11421 26074 11487 26077
rect 11053 26072 11487 26074
rect 11053 26016 11058 26072
rect 11114 26016 11426 26072
rect 11482 26016 11487 26072
rect 11053 26014 11487 26016
rect 11053 26011 11119 26014
rect 11421 26011 11487 26014
rect 16113 26074 16179 26077
rect 16430 26074 16436 26076
rect 16113 26072 16436 26074
rect 16113 26016 16118 26072
rect 16174 26016 16436 26072
rect 16113 26014 16436 26016
rect 16113 26011 16179 26014
rect 16430 26012 16436 26014
rect 16500 26012 16506 26076
rect 21541 26074 21607 26077
rect 24158 26074 24164 26076
rect 21541 26072 24164 26074
rect 21541 26016 21546 26072
rect 21602 26016 24164 26072
rect 21541 26014 24164 26016
rect 21541 26011 21607 26014
rect 24158 26012 24164 26014
rect 24228 26074 24234 26076
rect 24228 26014 31770 26074
rect 24228 26012 24234 26014
rect 5257 25938 5323 25941
rect 7966 25938 7972 25940
rect 5257 25936 7972 25938
rect 5257 25880 5262 25936
rect 5318 25880 7972 25936
rect 5257 25878 7972 25880
rect 5257 25875 5323 25878
rect 7966 25876 7972 25878
rect 8036 25938 8042 25940
rect 8477 25938 8543 25941
rect 8036 25936 8543 25938
rect 8036 25880 8482 25936
rect 8538 25880 8543 25936
rect 8036 25878 8543 25880
rect 8036 25876 8042 25878
rect 8477 25875 8543 25878
rect 11145 25938 11211 25941
rect 20713 25938 20779 25941
rect 11145 25936 20779 25938
rect 11145 25880 11150 25936
rect 11206 25880 20718 25936
rect 20774 25880 20779 25936
rect 11145 25878 20779 25880
rect 11145 25875 11211 25878
rect 20713 25875 20779 25878
rect 20897 25938 20963 25941
rect 30925 25938 30991 25941
rect 20897 25936 30991 25938
rect 20897 25880 20902 25936
rect 20958 25880 30930 25936
rect 30986 25880 30991 25936
rect 20897 25878 30991 25880
rect 31710 25938 31770 26014
rect 32489 25938 32555 25941
rect 31710 25936 32555 25938
rect 31710 25880 32494 25936
rect 32550 25880 32555 25936
rect 31710 25878 32555 25880
rect 20897 25875 20963 25878
rect 30925 25875 30991 25878
rect 32489 25875 32555 25878
rect 4429 25802 4495 25805
rect 9765 25802 9831 25805
rect 4429 25800 9831 25802
rect 4429 25744 4434 25800
rect 4490 25744 9770 25800
rect 9826 25744 9831 25800
rect 4429 25742 9831 25744
rect 4429 25739 4495 25742
rect 9765 25739 9831 25742
rect 13261 25802 13327 25805
rect 16389 25802 16455 25805
rect 13261 25800 16455 25802
rect 13261 25744 13266 25800
rect 13322 25744 16394 25800
rect 16450 25744 16455 25800
rect 13261 25742 16455 25744
rect 13261 25739 13327 25742
rect 16389 25739 16455 25742
rect 18137 25802 18203 25805
rect 24209 25802 24275 25805
rect 25221 25802 25287 25805
rect 18137 25800 25287 25802
rect 18137 25744 18142 25800
rect 18198 25744 24214 25800
rect 24270 25744 25226 25800
rect 25282 25744 25287 25800
rect 18137 25742 25287 25744
rect 18137 25739 18203 25742
rect 24209 25739 24275 25742
rect 25221 25739 25287 25742
rect 26141 25802 26207 25805
rect 26366 25802 26372 25804
rect 26141 25800 26372 25802
rect 26141 25744 26146 25800
rect 26202 25744 26372 25800
rect 26141 25742 26372 25744
rect 26141 25739 26207 25742
rect 26366 25740 26372 25742
rect 26436 25740 26442 25804
rect 27245 25802 27311 25805
rect 28625 25802 28691 25805
rect 27245 25800 28691 25802
rect 27245 25744 27250 25800
rect 27306 25744 28630 25800
rect 28686 25744 28691 25800
rect 27245 25742 28691 25744
rect 27245 25739 27311 25742
rect 28625 25739 28691 25742
rect 5993 25666 6059 25669
rect 6361 25666 6427 25669
rect 5993 25664 6427 25666
rect 5993 25608 5998 25664
rect 6054 25608 6366 25664
rect 6422 25608 6427 25664
rect 5993 25606 6427 25608
rect 5993 25603 6059 25606
rect 6361 25603 6427 25606
rect 6545 25666 6611 25669
rect 6862 25666 6868 25668
rect 6545 25664 6868 25666
rect 6545 25608 6550 25664
rect 6606 25608 6868 25664
rect 6545 25606 6868 25608
rect 6545 25603 6611 25606
rect 6862 25604 6868 25606
rect 6932 25604 6938 25668
rect 7230 25604 7236 25668
rect 7300 25666 7306 25668
rect 7373 25666 7439 25669
rect 11881 25668 11947 25669
rect 7300 25664 7439 25666
rect 7300 25608 7378 25664
rect 7434 25608 7439 25664
rect 7300 25606 7439 25608
rect 7300 25604 7306 25606
rect 7373 25603 7439 25606
rect 11830 25604 11836 25668
rect 11900 25666 11947 25668
rect 14733 25666 14799 25669
rect 11900 25664 14799 25666
rect 11942 25608 14738 25664
rect 14794 25608 14799 25664
rect 11900 25606 14799 25608
rect 11900 25604 11947 25606
rect 11881 25603 11947 25604
rect 14733 25603 14799 25606
rect 15837 25666 15903 25669
rect 20897 25666 20963 25669
rect 15837 25664 20963 25666
rect 15837 25608 15842 25664
rect 15898 25608 20902 25664
rect 20958 25608 20963 25664
rect 15837 25606 20963 25608
rect 15837 25603 15903 25606
rect 20897 25603 20963 25606
rect 23657 25666 23723 25669
rect 26233 25666 26299 25669
rect 26550 25666 26556 25668
rect 23657 25664 26556 25666
rect 23657 25608 23662 25664
rect 23718 25608 26238 25664
rect 26294 25608 26556 25664
rect 23657 25606 26556 25608
rect 23657 25603 23723 25606
rect 26233 25603 26299 25606
rect 26550 25604 26556 25606
rect 26620 25604 26626 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 5165 25530 5231 25533
rect 8201 25530 8267 25533
rect 5165 25528 8267 25530
rect 5165 25472 5170 25528
rect 5226 25472 8206 25528
rect 8262 25472 8267 25528
rect 5165 25470 8267 25472
rect 5165 25467 5231 25470
rect 8201 25467 8267 25470
rect 15929 25530 15995 25533
rect 18781 25530 18847 25533
rect 15929 25528 18847 25530
rect 15929 25472 15934 25528
rect 15990 25472 18786 25528
rect 18842 25472 18847 25528
rect 15929 25470 18847 25472
rect 15929 25467 15995 25470
rect 18781 25467 18847 25470
rect 19290 25470 26250 25530
rect 5809 25394 5875 25397
rect 6637 25394 6703 25397
rect 5809 25392 6703 25394
rect 5809 25336 5814 25392
rect 5870 25336 6642 25392
rect 6698 25336 6703 25392
rect 5809 25334 6703 25336
rect 5809 25331 5875 25334
rect 6637 25331 6703 25334
rect 9254 25332 9260 25396
rect 9324 25394 9330 25396
rect 9581 25394 9647 25397
rect 11513 25396 11579 25397
rect 9324 25392 9647 25394
rect 9324 25336 9586 25392
rect 9642 25336 9647 25392
rect 9324 25334 9647 25336
rect 9324 25332 9330 25334
rect 9581 25331 9647 25334
rect 11462 25332 11468 25396
rect 11532 25394 11579 25396
rect 12985 25394 13051 25397
rect 16614 25394 16620 25396
rect 11532 25392 11624 25394
rect 11574 25336 11624 25392
rect 11532 25334 11624 25336
rect 12985 25392 16620 25394
rect 12985 25336 12990 25392
rect 13046 25336 16620 25392
rect 12985 25334 16620 25336
rect 11532 25332 11579 25334
rect 11513 25331 11579 25332
rect 12985 25331 13051 25334
rect 16614 25332 16620 25334
rect 16684 25394 16690 25396
rect 18505 25394 18571 25397
rect 19290 25394 19350 25470
rect 16684 25392 19350 25394
rect 16684 25336 18510 25392
rect 18566 25336 19350 25392
rect 16684 25334 19350 25336
rect 19793 25394 19859 25397
rect 20294 25394 20300 25396
rect 19793 25392 20300 25394
rect 19793 25336 19798 25392
rect 19854 25336 20300 25392
rect 19793 25334 20300 25336
rect 16684 25332 16690 25334
rect 18505 25331 18571 25334
rect 19793 25331 19859 25334
rect 20294 25332 20300 25334
rect 20364 25332 20370 25396
rect 20621 25394 20687 25397
rect 26190 25394 26250 25470
rect 26918 25468 26924 25532
rect 26988 25530 26994 25532
rect 32949 25530 33015 25533
rect 26988 25528 33015 25530
rect 26988 25472 32954 25528
rect 33010 25472 33015 25528
rect 26988 25470 33015 25472
rect 26988 25468 26994 25470
rect 32949 25467 33015 25470
rect 27981 25394 28047 25397
rect 20621 25392 23122 25394
rect 20621 25336 20626 25392
rect 20682 25336 23122 25392
rect 20621 25334 23122 25336
rect 26190 25392 28047 25394
rect 26190 25336 27986 25392
rect 28042 25336 28047 25392
rect 26190 25334 28047 25336
rect 20621 25331 20687 25334
rect 3417 25258 3483 25261
rect 11145 25258 11211 25261
rect 17493 25260 17559 25261
rect 16246 25258 16252 25260
rect 3417 25256 11211 25258
rect 3417 25200 3422 25256
rect 3478 25200 11150 25256
rect 11206 25200 11211 25256
rect 3417 25198 11211 25200
rect 3417 25195 3483 25198
rect 11145 25195 11211 25198
rect 15518 25198 16252 25258
rect 0 25122 800 25152
rect 2773 25122 2839 25125
rect 0 25120 2839 25122
rect 0 25064 2778 25120
rect 2834 25064 2839 25120
rect 0 25062 2839 25064
rect 0 25032 800 25062
rect 2773 25059 2839 25062
rect 5809 25122 5875 25125
rect 6453 25122 6519 25125
rect 7189 25124 7255 25125
rect 7189 25122 7236 25124
rect 5809 25120 6519 25122
rect 5809 25064 5814 25120
rect 5870 25064 6458 25120
rect 6514 25064 6519 25120
rect 5809 25062 6519 25064
rect 7144 25120 7236 25122
rect 7144 25064 7194 25120
rect 7144 25062 7236 25064
rect 5809 25059 5875 25062
rect 6453 25059 6519 25062
rect 7189 25060 7236 25062
rect 7300 25060 7306 25124
rect 9857 25122 9923 25125
rect 10869 25122 10935 25125
rect 12249 25122 12315 25125
rect 9857 25120 12315 25122
rect 9857 25064 9862 25120
rect 9918 25064 10874 25120
rect 10930 25064 12254 25120
rect 12310 25064 12315 25120
rect 9857 25062 12315 25064
rect 7189 25059 7255 25060
rect 9857 25059 9923 25062
rect 10869 25059 10935 25062
rect 12249 25059 12315 25062
rect 15377 25122 15443 25125
rect 15518 25124 15578 25198
rect 16246 25196 16252 25198
rect 16316 25196 16322 25260
rect 17493 25258 17540 25260
rect 17452 25256 17540 25258
rect 17604 25258 17610 25260
rect 22461 25258 22527 25261
rect 23062 25260 23122 25334
rect 27981 25331 28047 25334
rect 17604 25256 22527 25258
rect 17452 25200 17498 25256
rect 17604 25200 22466 25256
rect 22522 25200 22527 25256
rect 17452 25198 17540 25200
rect 17493 25196 17540 25198
rect 17604 25198 22527 25200
rect 17604 25196 17610 25198
rect 17493 25195 17559 25196
rect 22461 25195 22527 25198
rect 23054 25196 23060 25260
rect 23124 25258 23130 25260
rect 23381 25258 23447 25261
rect 23124 25256 23447 25258
rect 23124 25200 23386 25256
rect 23442 25200 23447 25256
rect 23124 25198 23447 25200
rect 27984 25258 28044 25331
rect 30005 25258 30071 25261
rect 27984 25256 30071 25258
rect 27984 25200 30010 25256
rect 30066 25200 30071 25256
rect 27984 25198 30071 25200
rect 23124 25196 23130 25198
rect 23381 25195 23447 25198
rect 30005 25195 30071 25198
rect 20161 25124 20227 25125
rect 15510 25122 15516 25124
rect 15377 25120 15516 25122
rect 15377 25064 15382 25120
rect 15438 25064 15516 25120
rect 15377 25062 15516 25064
rect 15377 25059 15443 25062
rect 15510 25060 15516 25062
rect 15580 25060 15586 25124
rect 20110 25122 20116 25124
rect 20034 25062 20116 25122
rect 20180 25122 20227 25124
rect 20345 25122 20411 25125
rect 24301 25122 24367 25125
rect 20180 25120 24367 25122
rect 20222 25064 20350 25120
rect 20406 25064 24306 25120
rect 24362 25064 24367 25120
rect 20110 25060 20116 25062
rect 20180 25062 24367 25064
rect 20180 25060 20227 25062
rect 20161 25059 20227 25060
rect 20345 25059 20411 25062
rect 24301 25059 24367 25062
rect 26509 25122 26575 25125
rect 29729 25122 29795 25125
rect 26509 25120 29795 25122
rect 26509 25064 26514 25120
rect 26570 25064 29734 25120
rect 29790 25064 29795 25120
rect 26509 25062 29795 25064
rect 26509 25059 26575 25062
rect 29729 25059 29795 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4705 24986 4771 24989
rect 6545 24986 6611 24989
rect 4705 24984 6611 24986
rect 4705 24928 4710 24984
rect 4766 24928 6550 24984
rect 6606 24928 6611 24984
rect 4705 24926 6611 24928
rect 4705 24923 4771 24926
rect 6545 24923 6611 24926
rect 6678 24924 6684 24988
rect 6748 24986 6754 24988
rect 7005 24986 7071 24989
rect 6748 24984 7071 24986
rect 6748 24928 7010 24984
rect 7066 24928 7071 24984
rect 6748 24926 7071 24928
rect 6748 24924 6754 24926
rect 7005 24923 7071 24926
rect 11881 24986 11947 24989
rect 13721 24986 13787 24989
rect 14406 24986 14412 24988
rect 11881 24984 14412 24986
rect 11881 24928 11886 24984
rect 11942 24928 13726 24984
rect 13782 24928 14412 24984
rect 11881 24926 14412 24928
rect 11881 24923 11947 24926
rect 13721 24923 13787 24926
rect 14406 24924 14412 24926
rect 14476 24924 14482 24988
rect 14641 24986 14707 24989
rect 16665 24986 16731 24989
rect 17217 24988 17283 24989
rect 14641 24984 16731 24986
rect 14641 24928 14646 24984
rect 14702 24928 16670 24984
rect 16726 24928 16731 24984
rect 14641 24926 16731 24928
rect 14641 24923 14707 24926
rect 16665 24923 16731 24926
rect 17166 24924 17172 24988
rect 17236 24986 17283 24988
rect 20069 24986 20135 24989
rect 20437 24988 20503 24989
rect 20294 24986 20300 24988
rect 17236 24984 17328 24986
rect 17278 24928 17328 24984
rect 17236 24926 17328 24928
rect 20069 24984 20300 24986
rect 20069 24928 20074 24984
rect 20130 24928 20300 24984
rect 20069 24926 20300 24928
rect 17236 24924 17283 24926
rect 17217 24923 17283 24924
rect 20069 24923 20135 24926
rect 20294 24924 20300 24926
rect 20364 24924 20370 24988
rect 20437 24984 20484 24988
rect 20548 24986 20554 24988
rect 20437 24928 20442 24984
rect 20437 24924 20484 24928
rect 20548 24926 20594 24986
rect 20548 24924 20554 24926
rect 21398 24924 21404 24988
rect 21468 24986 21474 24988
rect 21541 24986 21607 24989
rect 21468 24984 21607 24986
rect 21468 24928 21546 24984
rect 21602 24928 21607 24984
rect 21468 24926 21607 24928
rect 21468 24924 21474 24926
rect 20437 24923 20503 24924
rect 21541 24923 21607 24926
rect 22737 24986 22803 24989
rect 24577 24986 24643 24989
rect 22737 24984 24643 24986
rect 22737 24928 22742 24984
rect 22798 24928 24582 24984
rect 24638 24928 24643 24984
rect 22737 24926 24643 24928
rect 22737 24923 22803 24926
rect 24577 24923 24643 24926
rect 5574 24788 5580 24852
rect 5644 24788 5650 24852
rect 7046 24788 7052 24852
rect 7116 24850 7122 24852
rect 7557 24850 7623 24853
rect 7116 24848 7623 24850
rect 7116 24792 7562 24848
rect 7618 24792 7623 24848
rect 7116 24790 7623 24792
rect 7116 24788 7122 24790
rect 4613 24714 4679 24717
rect 5582 24714 5642 24788
rect 7557 24787 7623 24790
rect 9029 24850 9095 24853
rect 10225 24850 10291 24853
rect 9029 24848 10291 24850
rect 9029 24792 9034 24848
rect 9090 24792 10230 24848
rect 10286 24792 10291 24848
rect 9029 24790 10291 24792
rect 9029 24787 9095 24790
rect 10225 24787 10291 24790
rect 13721 24850 13787 24853
rect 21909 24850 21975 24853
rect 13721 24848 21975 24850
rect 13721 24792 13726 24848
rect 13782 24792 21914 24848
rect 21970 24792 21975 24848
rect 13721 24790 21975 24792
rect 13721 24787 13787 24790
rect 21909 24787 21975 24790
rect 6269 24714 6335 24717
rect 7649 24716 7715 24717
rect 4613 24712 5090 24714
rect 4613 24656 4618 24712
rect 4674 24656 5090 24712
rect 4613 24654 5090 24656
rect 5582 24712 6335 24714
rect 5582 24656 6274 24712
rect 6330 24656 6335 24712
rect 5582 24654 6335 24656
rect 4613 24651 4679 24654
rect 5030 24578 5090 24654
rect 6269 24651 6335 24654
rect 7598 24652 7604 24716
rect 7668 24714 7715 24716
rect 18965 24716 19031 24717
rect 7668 24712 7760 24714
rect 7710 24656 7760 24712
rect 7668 24654 7760 24656
rect 18965 24712 19012 24716
rect 19076 24714 19082 24716
rect 19701 24714 19767 24717
rect 20897 24714 20963 24717
rect 18965 24656 18970 24712
rect 7668 24652 7715 24654
rect 7649 24651 7715 24652
rect 18965 24652 19012 24656
rect 19076 24654 19122 24714
rect 19701 24712 20963 24714
rect 19701 24656 19706 24712
rect 19762 24656 20902 24712
rect 20958 24656 20963 24712
rect 19701 24654 20963 24656
rect 19076 24652 19082 24654
rect 18965 24651 19031 24652
rect 19701 24651 19767 24654
rect 20897 24651 20963 24654
rect 21265 24714 21331 24717
rect 24393 24714 24459 24717
rect 21265 24712 24459 24714
rect 21265 24656 21270 24712
rect 21326 24656 24398 24712
rect 24454 24656 24459 24712
rect 21265 24654 24459 24656
rect 21265 24651 21331 24654
rect 24393 24651 24459 24654
rect 6361 24578 6427 24581
rect 5030 24576 6427 24578
rect 5030 24520 6366 24576
rect 6422 24520 6427 24576
rect 5030 24518 6427 24520
rect 6361 24515 6427 24518
rect 8385 24578 8451 24581
rect 14273 24578 14339 24581
rect 8385 24576 14339 24578
rect 8385 24520 8390 24576
rect 8446 24520 14278 24576
rect 14334 24520 14339 24576
rect 8385 24518 14339 24520
rect 8385 24515 8451 24518
rect 14273 24515 14339 24518
rect 15101 24578 15167 24581
rect 22829 24578 22895 24581
rect 15101 24576 22895 24578
rect 15101 24520 15106 24576
rect 15162 24520 22834 24576
rect 22890 24520 22895 24576
rect 15101 24518 22895 24520
rect 15101 24515 15167 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 5901 24442 5967 24445
rect 9489 24442 9555 24445
rect 5901 24440 9555 24442
rect 5901 24384 5906 24440
rect 5962 24384 9494 24440
rect 9550 24384 9555 24440
rect 5901 24382 9555 24384
rect 5901 24379 5967 24382
rect 9489 24379 9555 24382
rect 10685 24442 10751 24445
rect 11697 24442 11763 24445
rect 10685 24440 11763 24442
rect 10685 24384 10690 24440
rect 10746 24384 11702 24440
rect 11758 24384 11763 24440
rect 10685 24382 11763 24384
rect 10685 24379 10751 24382
rect 11697 24379 11763 24382
rect 13261 24442 13327 24445
rect 14089 24442 14155 24445
rect 13261 24440 14155 24442
rect 13261 24384 13266 24440
rect 13322 24384 14094 24440
rect 14150 24384 14155 24440
rect 13261 24382 14155 24384
rect 13261 24379 13327 24382
rect 14089 24379 14155 24382
rect 19057 24442 19123 24445
rect 21173 24442 21239 24445
rect 22001 24442 22067 24445
rect 19057 24440 22067 24442
rect 19057 24384 19062 24440
rect 19118 24384 21178 24440
rect 21234 24384 22006 24440
rect 22062 24384 22067 24440
rect 19057 24382 22067 24384
rect 19057 24379 19123 24382
rect 21173 24379 21239 24382
rect 22001 24379 22067 24382
rect 1577 24306 1643 24309
rect 12709 24306 12775 24309
rect 1577 24304 12775 24306
rect 1577 24248 1582 24304
rect 1638 24248 12714 24304
rect 12770 24248 12775 24304
rect 1577 24246 12775 24248
rect 1577 24243 1643 24246
rect 12709 24243 12775 24246
rect 13905 24306 13971 24309
rect 16849 24306 16915 24309
rect 13905 24304 16915 24306
rect 13905 24248 13910 24304
rect 13966 24248 16854 24304
rect 16910 24248 16915 24304
rect 13905 24246 16915 24248
rect 13905 24243 13971 24246
rect 16849 24243 16915 24246
rect 17217 24306 17283 24309
rect 17217 24304 21834 24306
rect 17217 24248 17222 24304
rect 17278 24248 21834 24304
rect 17217 24246 21834 24248
rect 17217 24243 17283 24246
rect 5533 24172 5599 24173
rect 5533 24170 5580 24172
rect 5492 24168 5580 24170
rect 5644 24170 5650 24172
rect 7925 24170 7991 24173
rect 5644 24168 7991 24170
rect 5492 24112 5538 24168
rect 5644 24112 7930 24168
rect 7986 24112 7991 24168
rect 5492 24110 5580 24112
rect 5533 24108 5580 24110
rect 5644 24110 7991 24112
rect 5644 24108 5650 24110
rect 5533 24107 5599 24108
rect 7925 24107 7991 24110
rect 8109 24170 8175 24173
rect 15745 24170 15811 24173
rect 8109 24168 15811 24170
rect 8109 24112 8114 24168
rect 8170 24112 15750 24168
rect 15806 24112 15811 24168
rect 8109 24110 15811 24112
rect 8109 24107 8175 24110
rect 15745 24107 15811 24110
rect 18597 24170 18663 24173
rect 20846 24170 20852 24172
rect 18597 24168 20852 24170
rect 18597 24112 18602 24168
rect 18658 24112 20852 24168
rect 18597 24110 20852 24112
rect 18597 24107 18663 24110
rect 20846 24108 20852 24110
rect 20916 24170 20922 24172
rect 21541 24170 21607 24173
rect 20916 24168 21607 24170
rect 20916 24112 21546 24168
rect 21602 24112 21607 24168
rect 20916 24110 21607 24112
rect 21774 24170 21834 24246
rect 21774 24110 22110 24170
rect 20916 24108 20922 24110
rect 21541 24107 21607 24110
rect 0 24034 800 24064
rect 1209 24034 1275 24037
rect 0 24032 1275 24034
rect 0 23976 1214 24032
rect 1270 23976 1275 24032
rect 0 23974 1275 23976
rect 0 23944 800 23974
rect 1209 23971 1275 23974
rect 6494 23972 6500 24036
rect 6564 24034 6570 24036
rect 6913 24034 6979 24037
rect 8201 24036 8267 24037
rect 6564 24032 6979 24034
rect 6564 23976 6918 24032
rect 6974 23976 6979 24032
rect 6564 23974 6979 23976
rect 6564 23972 6570 23974
rect 6913 23971 6979 23974
rect 8150 23972 8156 24036
rect 8220 24034 8267 24036
rect 9029 24034 9095 24037
rect 9765 24034 9831 24037
rect 17861 24034 17927 24037
rect 19057 24034 19123 24037
rect 8220 24032 8312 24034
rect 8262 23976 8312 24032
rect 8220 23974 8312 23976
rect 9029 24032 19123 24034
rect 9029 23976 9034 24032
rect 9090 23976 9770 24032
rect 9826 23976 17866 24032
rect 17922 23976 19062 24032
rect 19118 23976 19123 24032
rect 9029 23974 19123 23976
rect 8220 23972 8267 23974
rect 8201 23971 8267 23972
rect 9029 23971 9095 23974
rect 9765 23971 9831 23974
rect 17861 23971 17927 23974
rect 19057 23971 19123 23974
rect 19190 23972 19196 24036
rect 19260 24034 19266 24036
rect 19333 24034 19399 24037
rect 19260 24032 19399 24034
rect 19260 23976 19338 24032
rect 19394 23976 19399 24032
rect 19260 23974 19399 23976
rect 19260 23972 19266 23974
rect 19333 23971 19399 23974
rect 19977 24034 20043 24037
rect 21081 24034 21147 24037
rect 19977 24032 21147 24034
rect 19977 23976 19982 24032
rect 20038 23976 21086 24032
rect 21142 23976 21147 24032
rect 19977 23974 21147 23976
rect 22050 24034 22110 24110
rect 22553 24034 22619 24037
rect 22694 24036 22754 24518
rect 22829 24515 22895 24518
rect 23565 24578 23631 24581
rect 28165 24578 28231 24581
rect 23565 24576 28231 24578
rect 23565 24520 23570 24576
rect 23626 24520 28170 24576
rect 28226 24520 28231 24576
rect 23565 24518 28231 24520
rect 23565 24515 23631 24518
rect 28165 24515 28231 24518
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 25773 24170 25839 24173
rect 26877 24170 26943 24173
rect 25773 24168 26943 24170
rect 25773 24112 25778 24168
rect 25834 24112 26882 24168
rect 26938 24112 26943 24168
rect 25773 24110 26943 24112
rect 25773 24107 25839 24110
rect 26877 24107 26943 24110
rect 22050 24032 22619 24034
rect 22050 23976 22558 24032
rect 22614 23976 22619 24032
rect 22050 23974 22619 23976
rect 19977 23971 20043 23974
rect 21081 23971 21147 23974
rect 22553 23971 22619 23974
rect 22686 23972 22692 24036
rect 22756 23972 22762 24036
rect 22829 24034 22895 24037
rect 25957 24034 26023 24037
rect 22829 24032 26023 24034
rect 22829 23976 22834 24032
rect 22890 23976 25962 24032
rect 26018 23976 26023 24032
rect 22829 23974 26023 23976
rect 22829 23971 22895 23974
rect 25957 23971 26023 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4153 23898 4219 23901
rect 5073 23898 5139 23901
rect 4153 23896 5139 23898
rect 4153 23840 4158 23896
rect 4214 23840 5078 23896
rect 5134 23840 5139 23896
rect 4153 23838 5139 23840
rect 4153 23835 4219 23838
rect 5073 23835 5139 23838
rect 5257 23898 5323 23901
rect 5390 23898 5396 23900
rect 5257 23896 5396 23898
rect 5257 23840 5262 23896
rect 5318 23840 5396 23896
rect 5257 23838 5396 23840
rect 5257 23835 5323 23838
rect 5390 23836 5396 23838
rect 5460 23836 5466 23900
rect 6862 23836 6868 23900
rect 6932 23898 6938 23900
rect 7097 23898 7163 23901
rect 6932 23896 7163 23898
rect 6932 23840 7102 23896
rect 7158 23840 7163 23896
rect 6932 23838 7163 23840
rect 6932 23836 6938 23838
rect 7097 23835 7163 23838
rect 11053 23898 11119 23901
rect 12249 23898 12315 23901
rect 19425 23900 19491 23901
rect 19374 23898 19380 23900
rect 11053 23896 12315 23898
rect 11053 23840 11058 23896
rect 11114 23840 12254 23896
rect 12310 23840 12315 23896
rect 11053 23838 12315 23840
rect 19334 23838 19380 23898
rect 19444 23896 19491 23900
rect 21173 23900 21239 23901
rect 21173 23898 21220 23900
rect 19486 23840 19491 23896
rect 11053 23835 11119 23838
rect 12249 23835 12315 23838
rect 19374 23836 19380 23838
rect 19444 23836 19491 23840
rect 21128 23896 21220 23898
rect 21128 23840 21178 23896
rect 21128 23838 21220 23840
rect 19425 23835 19491 23836
rect 21173 23836 21220 23838
rect 21284 23836 21290 23900
rect 21909 23898 21975 23901
rect 25773 23898 25839 23901
rect 21909 23896 25839 23898
rect 21909 23840 21914 23896
rect 21970 23840 25778 23896
rect 25834 23840 25839 23896
rect 21909 23838 25839 23840
rect 21173 23835 21239 23836
rect 21909 23835 21975 23838
rect 25773 23835 25839 23838
rect 26141 23898 26207 23901
rect 26550 23898 26556 23900
rect 26141 23896 26556 23898
rect 26141 23840 26146 23896
rect 26202 23840 26556 23896
rect 26141 23838 26556 23840
rect 26141 23835 26207 23838
rect 26550 23836 26556 23838
rect 26620 23836 26626 23900
rect 3182 23700 3188 23764
rect 3252 23762 3258 23764
rect 12617 23762 12683 23765
rect 3252 23760 12683 23762
rect 3252 23704 12622 23760
rect 12678 23704 12683 23760
rect 3252 23702 12683 23704
rect 3252 23700 3258 23702
rect 12617 23699 12683 23702
rect 17309 23762 17375 23765
rect 19796 23762 20132 23796
rect 22001 23762 22067 23765
rect 17309 23760 22067 23762
rect 17309 23704 17314 23760
rect 17370 23736 22006 23760
rect 17370 23704 19856 23736
rect 17309 23702 19856 23704
rect 20072 23704 22006 23736
rect 22062 23704 22067 23760
rect 20072 23702 22067 23704
rect 17309 23699 17375 23702
rect 22001 23699 22067 23702
rect 24342 23700 24348 23764
rect 24412 23762 24418 23764
rect 28441 23762 28507 23765
rect 24412 23760 28507 23762
rect 24412 23704 28446 23760
rect 28502 23704 28507 23760
rect 24412 23702 28507 23704
rect 24412 23700 24418 23702
rect 28441 23699 28507 23702
rect 4521 23626 4587 23629
rect 5533 23626 5599 23629
rect 4521 23624 5599 23626
rect 4521 23568 4526 23624
rect 4582 23568 5538 23624
rect 5594 23568 5599 23624
rect 4521 23566 5599 23568
rect 4521 23563 4587 23566
rect 5533 23563 5599 23566
rect 6126 23564 6132 23628
rect 6196 23626 6202 23628
rect 6729 23626 6795 23629
rect 12065 23628 12131 23629
rect 6196 23624 6795 23626
rect 6196 23568 6734 23624
rect 6790 23568 6795 23624
rect 6196 23566 6795 23568
rect 6196 23564 6202 23566
rect 6729 23563 6795 23566
rect 12014 23564 12020 23628
rect 12084 23626 12131 23628
rect 31477 23626 31543 23629
rect 12084 23624 12176 23626
rect 12126 23568 12176 23624
rect 12084 23566 12176 23568
rect 17036 23624 31543 23626
rect 17036 23568 31482 23624
rect 31538 23568 31543 23624
rect 17036 23566 31543 23568
rect 12084 23564 12131 23566
rect 12065 23563 12131 23564
rect 5022 23428 5028 23492
rect 5092 23490 5098 23492
rect 5257 23490 5323 23493
rect 5092 23488 5323 23490
rect 5092 23432 5262 23488
rect 5318 23432 5323 23488
rect 5092 23430 5323 23432
rect 5092 23428 5098 23430
rect 5257 23427 5323 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 4705 23354 4771 23357
rect 5993 23354 6059 23357
rect 6126 23354 6132 23356
rect 4705 23352 6132 23354
rect 4705 23296 4710 23352
rect 4766 23296 5998 23352
rect 6054 23296 6132 23352
rect 4705 23294 6132 23296
rect 4705 23291 4771 23294
rect 5993 23291 6059 23294
rect 6126 23292 6132 23294
rect 6196 23354 6202 23356
rect 7005 23354 7071 23357
rect 6196 23352 7071 23354
rect 6196 23296 7010 23352
rect 7066 23296 7071 23352
rect 6196 23294 7071 23296
rect 6196 23292 6202 23294
rect 7005 23291 7071 23294
rect 7230 23292 7236 23356
rect 7300 23354 7306 23356
rect 7373 23354 7439 23357
rect 7300 23352 7439 23354
rect 7300 23296 7378 23352
rect 7434 23296 7439 23352
rect 7300 23294 7439 23296
rect 7300 23292 7306 23294
rect 7373 23291 7439 23294
rect 13629 23354 13695 23357
rect 16297 23354 16363 23357
rect 13629 23352 16363 23354
rect 13629 23296 13634 23352
rect 13690 23296 16302 23352
rect 16358 23296 16363 23352
rect 13629 23294 16363 23296
rect 13629 23291 13695 23294
rect 16297 23291 16363 23294
rect 17036 23221 17096 23566
rect 31477 23563 31543 23566
rect 17677 23492 17743 23493
rect 17677 23490 17724 23492
rect 17632 23488 17724 23490
rect 17632 23432 17682 23488
rect 17632 23430 17724 23432
rect 17677 23428 17724 23430
rect 17788 23428 17794 23492
rect 24301 23490 24367 23493
rect 26049 23490 26115 23493
rect 27153 23492 27219 23493
rect 19290 23430 21972 23490
rect 17677 23427 17743 23428
rect 18505 23354 18571 23357
rect 19290 23354 19350 23430
rect 21912 23357 21972 23430
rect 24301 23488 26115 23490
rect 24301 23432 24306 23488
rect 24362 23432 26054 23488
rect 26110 23432 26115 23488
rect 24301 23430 26115 23432
rect 24301 23427 24367 23430
rect 26049 23427 26115 23430
rect 27102 23428 27108 23492
rect 27172 23490 27219 23492
rect 27172 23488 27264 23490
rect 27214 23432 27264 23488
rect 27172 23430 27264 23432
rect 27172 23428 27219 23430
rect 27153 23427 27219 23428
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 18505 23352 19350 23354
rect 18505 23296 18510 23352
rect 18566 23296 19350 23352
rect 18505 23294 19350 23296
rect 19885 23354 19951 23357
rect 20662 23354 20668 23356
rect 19885 23352 20668 23354
rect 19885 23296 19890 23352
rect 19946 23296 20668 23352
rect 19885 23294 20668 23296
rect 18505 23291 18571 23294
rect 19885 23291 19951 23294
rect 20662 23292 20668 23294
rect 20732 23292 20738 23356
rect 21909 23352 21975 23357
rect 21909 23296 21914 23352
rect 21970 23296 21975 23352
rect 21909 23291 21975 23296
rect 22277 23354 22343 23357
rect 27889 23354 27955 23357
rect 22277 23352 27955 23354
rect 22277 23296 22282 23352
rect 22338 23296 27894 23352
rect 27950 23296 27955 23352
rect 22277 23294 27955 23296
rect 22277 23291 22343 23294
rect 27889 23291 27955 23294
rect 3325 23218 3391 23221
rect 5809 23218 5875 23221
rect 3325 23216 5875 23218
rect 3325 23160 3330 23216
rect 3386 23160 5814 23216
rect 5870 23160 5875 23216
rect 3325 23158 5875 23160
rect 3325 23155 3391 23158
rect 5809 23155 5875 23158
rect 10593 23218 10659 23221
rect 14917 23218 14983 23221
rect 10593 23216 14983 23218
rect 10593 23160 10598 23216
rect 10654 23160 14922 23216
rect 14978 23160 14983 23216
rect 10593 23158 14983 23160
rect 10593 23155 10659 23158
rect 14917 23155 14983 23158
rect 17033 23216 17099 23221
rect 17033 23160 17038 23216
rect 17094 23160 17099 23216
rect 17033 23155 17099 23160
rect 17217 23218 17283 23221
rect 17769 23218 17835 23221
rect 17217 23216 17835 23218
rect 17217 23160 17222 23216
rect 17278 23160 17774 23216
rect 17830 23160 17835 23216
rect 17217 23158 17835 23160
rect 17217 23155 17283 23158
rect 17769 23155 17835 23158
rect 18045 23218 18111 23221
rect 24577 23218 24643 23221
rect 18045 23216 24643 23218
rect 18045 23160 18050 23216
rect 18106 23160 24582 23216
rect 24638 23160 24643 23216
rect 18045 23158 24643 23160
rect 18045 23155 18111 23158
rect 24577 23155 24643 23158
rect 24853 23218 24919 23221
rect 26325 23218 26391 23221
rect 24853 23216 26391 23218
rect 24853 23160 24858 23216
rect 24914 23160 26330 23216
rect 26386 23160 26391 23216
rect 24853 23158 26391 23160
rect 24853 23155 24919 23158
rect 26325 23155 26391 23158
rect 3049 23082 3115 23085
rect 6361 23082 6427 23085
rect 6913 23084 6979 23085
rect 3049 23080 6427 23082
rect 3049 23024 3054 23080
rect 3110 23024 6366 23080
rect 6422 23024 6427 23080
rect 3049 23022 6427 23024
rect 3049 23019 3115 23022
rect 6361 23019 6427 23022
rect 6862 23020 6868 23084
rect 6932 23082 6979 23084
rect 6932 23080 7024 23082
rect 6974 23024 7024 23080
rect 6932 23022 7024 23024
rect 6932 23020 6979 23022
rect 9622 23020 9628 23084
rect 9692 23082 9698 23084
rect 11053 23082 11119 23085
rect 9692 23080 11119 23082
rect 9692 23024 11058 23080
rect 11114 23024 11119 23080
rect 9692 23022 11119 23024
rect 9692 23020 9698 23022
rect 6913 23019 6979 23020
rect 11053 23019 11119 23022
rect 11605 23082 11671 23085
rect 16430 23082 16436 23084
rect 11605 23080 16436 23082
rect 11605 23024 11610 23080
rect 11666 23024 16436 23080
rect 11605 23022 16436 23024
rect 11605 23019 11671 23022
rect 16430 23020 16436 23022
rect 16500 23020 16506 23084
rect 16982 23020 16988 23084
rect 17052 23082 17058 23084
rect 17309 23082 17375 23085
rect 17052 23080 17375 23082
rect 17052 23024 17314 23080
rect 17370 23024 17375 23080
rect 17052 23022 17375 23024
rect 17052 23020 17058 23022
rect 17309 23019 17375 23022
rect 18321 23082 18387 23085
rect 25405 23082 25471 23085
rect 28533 23084 28599 23085
rect 28533 23082 28580 23084
rect 18321 23080 25471 23082
rect 18321 23024 18326 23080
rect 18382 23024 25410 23080
rect 25466 23024 25471 23080
rect 18321 23022 25471 23024
rect 28488 23080 28580 23082
rect 28488 23024 28538 23080
rect 28488 23022 28580 23024
rect 18321 23019 18387 23022
rect 25405 23019 25471 23022
rect 28533 23020 28580 23022
rect 28644 23020 28650 23084
rect 28533 23019 28599 23020
rect 0 22946 800 22976
rect 1209 22946 1275 22949
rect 0 22944 1275 22946
rect 0 22888 1214 22944
rect 1270 22888 1275 22944
rect 0 22886 1275 22888
rect 0 22856 800 22886
rect 1209 22883 1275 22886
rect 2957 22946 3023 22949
rect 2957 22944 5136 22946
rect 2957 22888 2962 22944
rect 3018 22888 5136 22944
rect 2957 22886 5136 22888
rect 2957 22883 3023 22886
rect 3918 22748 3924 22812
rect 3988 22810 3994 22812
rect 4797 22810 4863 22813
rect 3988 22808 4863 22810
rect 3988 22752 4802 22808
rect 4858 22752 4863 22808
rect 3988 22750 4863 22752
rect 5076 22810 5136 22886
rect 5206 22884 5212 22948
rect 5276 22946 5282 22948
rect 6913 22946 6979 22949
rect 5276 22944 6979 22946
rect 5276 22888 6918 22944
rect 6974 22888 6979 22944
rect 5276 22886 6979 22888
rect 5276 22884 5282 22886
rect 6913 22883 6979 22886
rect 9581 22946 9647 22949
rect 10358 22946 10364 22948
rect 9581 22944 10364 22946
rect 9581 22888 9586 22944
rect 9642 22888 10364 22944
rect 9581 22886 10364 22888
rect 9581 22883 9647 22886
rect 10358 22884 10364 22886
rect 10428 22884 10434 22948
rect 10593 22946 10659 22949
rect 13353 22946 13419 22949
rect 10593 22944 13419 22946
rect 10593 22888 10598 22944
rect 10654 22888 13358 22944
rect 13414 22888 13419 22944
rect 10593 22886 13419 22888
rect 10593 22883 10659 22886
rect 13353 22883 13419 22886
rect 17309 22946 17375 22949
rect 18086 22946 18092 22948
rect 17309 22944 18092 22946
rect 17309 22888 17314 22944
rect 17370 22888 18092 22944
rect 17309 22886 18092 22888
rect 17309 22883 17375 22886
rect 18086 22884 18092 22886
rect 18156 22946 18162 22948
rect 18781 22946 18847 22949
rect 18156 22944 18847 22946
rect 18156 22888 18786 22944
rect 18842 22888 18847 22944
rect 18156 22886 18847 22888
rect 18156 22884 18162 22886
rect 18781 22883 18847 22886
rect 20253 22946 20319 22949
rect 22185 22946 22251 22949
rect 28257 22946 28323 22949
rect 20253 22944 28323 22946
rect 20253 22888 20258 22944
rect 20314 22888 22190 22944
rect 22246 22888 28262 22944
rect 28318 22888 28323 22944
rect 20253 22886 28323 22888
rect 20253 22883 20319 22886
rect 22185 22883 22251 22886
rect 28257 22883 28323 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 5349 22810 5415 22813
rect 5076 22808 5415 22810
rect 5076 22752 5354 22808
rect 5410 22752 5415 22808
rect 5076 22750 5415 22752
rect 3988 22748 3994 22750
rect 4797 22747 4863 22750
rect 5349 22747 5415 22750
rect 11237 22810 11303 22813
rect 11830 22810 11836 22812
rect 11237 22808 11836 22810
rect 11237 22752 11242 22808
rect 11298 22752 11836 22808
rect 11237 22750 11836 22752
rect 11237 22747 11303 22750
rect 11830 22748 11836 22750
rect 11900 22748 11906 22812
rect 18270 22748 18276 22812
rect 18340 22810 18346 22812
rect 18873 22810 18939 22813
rect 18340 22808 18939 22810
rect 18340 22752 18878 22808
rect 18934 22752 18939 22808
rect 18340 22750 18939 22752
rect 18340 22748 18346 22750
rect 18873 22747 18939 22750
rect 20621 22810 20687 22813
rect 23013 22810 23079 22813
rect 27889 22810 27955 22813
rect 20621 22808 21834 22810
rect 20621 22752 20626 22808
rect 20682 22752 21834 22808
rect 20621 22750 21834 22752
rect 20621 22747 20687 22750
rect 3049 22674 3115 22677
rect 9029 22674 9095 22677
rect 3049 22672 9095 22674
rect 3049 22616 3054 22672
rect 3110 22616 9034 22672
rect 9090 22616 9095 22672
rect 3049 22614 9095 22616
rect 3049 22611 3115 22614
rect 9029 22611 9095 22614
rect 10777 22674 10843 22677
rect 11973 22674 12039 22677
rect 10777 22672 12039 22674
rect 10777 22616 10782 22672
rect 10838 22616 11978 22672
rect 12034 22616 12039 22672
rect 10777 22614 12039 22616
rect 10777 22611 10843 22614
rect 11973 22611 12039 22614
rect 17217 22674 17283 22677
rect 17217 22672 18752 22674
rect 17217 22616 17222 22672
rect 17278 22616 18752 22672
rect 17217 22614 18752 22616
rect 17217 22611 17283 22614
rect 4245 22538 4311 22541
rect 5165 22538 5231 22541
rect 4245 22536 5231 22538
rect 4245 22480 4250 22536
rect 4306 22480 5170 22536
rect 5226 22480 5231 22536
rect 4245 22478 5231 22480
rect 4245 22475 4311 22478
rect 5165 22475 5231 22478
rect 5349 22538 5415 22541
rect 6085 22538 6151 22541
rect 5349 22536 6151 22538
rect 5349 22480 5354 22536
rect 5410 22480 6090 22536
rect 6146 22480 6151 22536
rect 5349 22478 6151 22480
rect 5349 22475 5415 22478
rect 6085 22475 6151 22478
rect 6310 22476 6316 22540
rect 6380 22538 6386 22540
rect 6545 22538 6611 22541
rect 6380 22536 6611 22538
rect 6380 22480 6550 22536
rect 6606 22480 6611 22536
rect 6380 22478 6611 22480
rect 6380 22476 6386 22478
rect 6545 22475 6611 22478
rect 7414 22476 7420 22540
rect 7484 22538 7490 22540
rect 7557 22538 7623 22541
rect 7484 22536 7623 22538
rect 7484 22480 7562 22536
rect 7618 22480 7623 22536
rect 7484 22478 7623 22480
rect 7484 22476 7490 22478
rect 7557 22475 7623 22478
rect 9254 22476 9260 22540
rect 9324 22538 9330 22540
rect 9489 22538 9555 22541
rect 9324 22536 9555 22538
rect 9324 22480 9494 22536
rect 9550 22480 9555 22536
rect 9324 22478 9555 22480
rect 9324 22476 9330 22478
rect 9489 22475 9555 22478
rect 10869 22538 10935 22541
rect 11605 22538 11671 22541
rect 10869 22536 11671 22538
rect 10869 22480 10874 22536
rect 10930 22480 11610 22536
rect 11666 22480 11671 22536
rect 10869 22478 11671 22480
rect 10869 22475 10935 22478
rect 11605 22475 11671 22478
rect 12525 22540 12591 22541
rect 12525 22536 12572 22540
rect 12636 22538 12642 22540
rect 15929 22538 15995 22541
rect 17401 22538 17467 22541
rect 12525 22480 12530 22536
rect 12525 22476 12572 22480
rect 12636 22478 12682 22538
rect 15929 22536 17467 22538
rect 15929 22480 15934 22536
rect 15990 22480 17406 22536
rect 17462 22480 17467 22536
rect 15929 22478 17467 22480
rect 18692 22538 18752 22614
rect 19374 22612 19380 22676
rect 19444 22674 19450 22676
rect 19609 22674 19675 22677
rect 19444 22672 19675 22674
rect 19444 22616 19614 22672
rect 19670 22616 19675 22672
rect 19444 22614 19675 22616
rect 19444 22612 19450 22614
rect 19609 22611 19675 22614
rect 19793 22674 19859 22677
rect 21633 22674 21699 22677
rect 19793 22672 21699 22674
rect 19793 22616 19798 22672
rect 19854 22616 21638 22672
rect 21694 22616 21699 22672
rect 19793 22614 21699 22616
rect 21774 22674 21834 22750
rect 23013 22808 27955 22810
rect 23013 22752 23018 22808
rect 23074 22752 27894 22808
rect 27950 22752 27955 22808
rect 23013 22750 27955 22752
rect 23013 22747 23079 22750
rect 27889 22747 27955 22750
rect 24393 22674 24459 22677
rect 21774 22672 24459 22674
rect 21774 22616 24398 22672
rect 24454 22616 24459 22672
rect 21774 22614 24459 22616
rect 19793 22611 19859 22614
rect 21633 22611 21699 22614
rect 24393 22611 24459 22614
rect 19241 22538 19307 22541
rect 25865 22538 25931 22541
rect 18692 22536 25931 22538
rect 18692 22480 19246 22536
rect 19302 22480 25870 22536
rect 25926 22480 25931 22536
rect 18692 22478 25931 22480
rect 12636 22476 12642 22478
rect 12525 22475 12591 22476
rect 15929 22475 15995 22478
rect 17401 22475 17467 22478
rect 19241 22475 19307 22478
rect 25865 22475 25931 22478
rect 27838 22476 27844 22540
rect 27908 22538 27914 22540
rect 28349 22538 28415 22541
rect 27908 22536 28415 22538
rect 27908 22480 28354 22536
rect 28410 22480 28415 22536
rect 27908 22478 28415 22480
rect 27908 22476 27914 22478
rect 28349 22475 28415 22478
rect 5073 22402 5139 22405
rect 5901 22404 5967 22405
rect 5390 22402 5396 22404
rect 5073 22400 5396 22402
rect 5073 22344 5078 22400
rect 5134 22344 5396 22400
rect 5073 22342 5396 22344
rect 5073 22339 5139 22342
rect 5390 22340 5396 22342
rect 5460 22340 5466 22404
rect 5901 22400 5948 22404
rect 6012 22402 6018 22404
rect 6269 22402 6335 22405
rect 8385 22402 8451 22405
rect 5901 22344 5906 22400
rect 5901 22340 5948 22344
rect 6012 22342 6058 22402
rect 6269 22400 8451 22402
rect 6269 22344 6274 22400
rect 6330 22344 8390 22400
rect 8446 22344 8451 22400
rect 6269 22342 8451 22344
rect 6012 22340 6018 22342
rect 5901 22339 5967 22340
rect 6269 22339 6335 22342
rect 8385 22339 8451 22342
rect 10409 22402 10475 22405
rect 10777 22402 10843 22405
rect 11421 22402 11487 22405
rect 10409 22400 11487 22402
rect 10409 22344 10414 22400
rect 10470 22344 10782 22400
rect 10838 22344 11426 22400
rect 11482 22344 11487 22400
rect 10409 22342 11487 22344
rect 10409 22339 10475 22342
rect 10777 22339 10843 22342
rect 11421 22339 11487 22342
rect 15009 22402 15075 22405
rect 15142 22402 15148 22404
rect 15009 22400 15148 22402
rect 15009 22344 15014 22400
rect 15070 22344 15148 22400
rect 15009 22342 15148 22344
rect 15009 22339 15075 22342
rect 15142 22340 15148 22342
rect 15212 22340 15218 22404
rect 17585 22402 17651 22405
rect 18638 22402 18644 22404
rect 17585 22400 18644 22402
rect 17585 22344 17590 22400
rect 17646 22344 18644 22400
rect 17585 22342 18644 22344
rect 17585 22339 17651 22342
rect 18638 22340 18644 22342
rect 18708 22402 18714 22404
rect 18965 22402 19031 22405
rect 20069 22404 20135 22405
rect 20069 22402 20116 22404
rect 18708 22400 19031 22402
rect 18708 22344 18970 22400
rect 19026 22344 19031 22400
rect 18708 22342 19031 22344
rect 20024 22400 20116 22402
rect 20024 22344 20074 22400
rect 20024 22342 20116 22344
rect 18708 22340 18714 22342
rect 18965 22339 19031 22342
rect 20069 22340 20116 22342
rect 20180 22340 20186 22404
rect 20529 22400 20595 22405
rect 21541 22404 21607 22405
rect 21541 22402 21588 22404
rect 20529 22344 20534 22400
rect 20590 22344 20595 22400
rect 20069 22339 20135 22340
rect 20529 22339 20595 22344
rect 21496 22400 21588 22402
rect 21496 22344 21546 22400
rect 21496 22342 21588 22344
rect 21541 22340 21588 22342
rect 21652 22340 21658 22404
rect 21817 22402 21883 22405
rect 28533 22402 28599 22405
rect 21817 22400 28599 22402
rect 21817 22344 21822 22400
rect 21878 22344 28538 22400
rect 28594 22344 28599 22400
rect 21817 22342 28599 22344
rect 21541 22339 21607 22340
rect 21817 22339 21883 22342
rect 28533 22339 28599 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 7557 22266 7623 22269
rect 4662 22264 7623 22266
rect 4662 22208 7562 22264
rect 7618 22208 7623 22264
rect 4662 22206 7623 22208
rect 2037 22130 2103 22133
rect 4662 22130 4722 22206
rect 7557 22203 7623 22206
rect 8293 22268 8359 22269
rect 8293 22264 8340 22268
rect 8404 22266 8410 22268
rect 11881 22266 11947 22269
rect 8293 22208 8298 22264
rect 8293 22204 8340 22208
rect 8404 22206 8450 22266
rect 9630 22264 11947 22266
rect 9630 22208 11886 22264
rect 11942 22208 11947 22264
rect 9630 22206 11947 22208
rect 8404 22204 8410 22206
rect 8293 22203 8359 22204
rect 4981 22130 5047 22133
rect 2037 22128 4722 22130
rect 2037 22072 2042 22128
rect 2098 22072 4722 22128
rect 2037 22070 4722 22072
rect 4846 22128 5047 22130
rect 4846 22072 4986 22128
rect 5042 22072 5047 22128
rect 4846 22070 5047 22072
rect 2037 22067 2103 22070
rect 3601 21994 3667 21997
rect 4245 21994 4311 21997
rect 4846 21994 4906 22070
rect 4981 22067 5047 22070
rect 5349 22130 5415 22133
rect 5574 22130 5580 22132
rect 5349 22128 5580 22130
rect 5349 22072 5354 22128
rect 5410 22072 5580 22128
rect 5349 22070 5580 22072
rect 5349 22067 5415 22070
rect 5574 22068 5580 22070
rect 5644 22068 5650 22132
rect 5901 22130 5967 22133
rect 6913 22130 6979 22133
rect 5901 22128 6979 22130
rect 5901 22072 5906 22128
rect 5962 22072 6918 22128
rect 6974 22072 6979 22128
rect 5901 22070 6979 22072
rect 5901 22067 5967 22070
rect 6913 22067 6979 22070
rect 9397 22130 9463 22133
rect 9630 22130 9690 22206
rect 11881 22203 11947 22206
rect 18321 22266 18387 22269
rect 18505 22266 18571 22269
rect 18321 22264 18571 22266
rect 18321 22208 18326 22264
rect 18382 22208 18510 22264
rect 18566 22208 18571 22264
rect 18321 22206 18571 22208
rect 18321 22203 18387 22206
rect 18505 22203 18571 22206
rect 18965 22266 19031 22269
rect 20345 22266 20411 22269
rect 18965 22264 20411 22266
rect 18965 22208 18970 22264
rect 19026 22208 20350 22264
rect 20406 22208 20411 22264
rect 18965 22206 20411 22208
rect 20532 22266 20592 22339
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 25957 22266 26023 22269
rect 20532 22264 26023 22266
rect 20532 22208 25962 22264
rect 26018 22208 26023 22264
rect 20532 22206 26023 22208
rect 18965 22203 19031 22206
rect 20345 22203 20411 22206
rect 25957 22203 26023 22206
rect 9397 22128 9690 22130
rect 9397 22072 9402 22128
rect 9458 22072 9690 22128
rect 9397 22070 9690 22072
rect 9397 22067 9463 22070
rect 9990 22068 9996 22132
rect 10060 22130 10066 22132
rect 10133 22130 10199 22133
rect 10060 22128 10199 22130
rect 10060 22072 10138 22128
rect 10194 22072 10199 22128
rect 10060 22070 10199 22072
rect 10060 22068 10066 22070
rect 10133 22067 10199 22070
rect 16481 22130 16547 22133
rect 16941 22130 17007 22133
rect 20161 22130 20227 22133
rect 16481 22128 20227 22130
rect 16481 22072 16486 22128
rect 16542 22072 16946 22128
rect 17002 22072 20166 22128
rect 20222 22072 20227 22128
rect 16481 22070 20227 22072
rect 16481 22067 16547 22070
rect 16941 22067 17007 22070
rect 20161 22067 20227 22070
rect 20294 22068 20300 22132
rect 20364 22130 20370 22132
rect 20529 22130 20595 22133
rect 20364 22128 20595 22130
rect 20364 22072 20534 22128
rect 20590 22072 20595 22128
rect 20364 22070 20595 22072
rect 20364 22068 20370 22070
rect 20529 22067 20595 22070
rect 21173 22130 21239 22133
rect 23381 22132 23447 22133
rect 21173 22128 23306 22130
rect 21173 22072 21178 22128
rect 21234 22072 23306 22128
rect 21173 22070 23306 22072
rect 21173 22067 21239 22070
rect 3601 21992 4906 21994
rect 3601 21936 3606 21992
rect 3662 21936 4250 21992
rect 4306 21936 4906 21992
rect 3601 21934 4906 21936
rect 4981 21996 5047 21997
rect 4981 21992 5028 21996
rect 5092 21994 5098 21996
rect 7281 21994 7347 21997
rect 10501 21994 10567 21997
rect 5092 21992 7347 21994
rect 4981 21936 4986 21992
rect 5092 21936 7286 21992
rect 7342 21936 7347 21992
rect 3601 21931 3667 21934
rect 4245 21931 4311 21934
rect 4981 21932 5028 21936
rect 5092 21934 7347 21936
rect 5092 21932 5098 21934
rect 4981 21931 5047 21932
rect 7281 21931 7347 21934
rect 8250 21992 10567 21994
rect 8250 21936 10506 21992
rect 10562 21936 10567 21992
rect 8250 21934 10567 21936
rect 0 21858 800 21888
rect 1209 21858 1275 21861
rect 0 21856 1275 21858
rect 0 21800 1214 21856
rect 1270 21800 1275 21856
rect 0 21798 1275 21800
rect 0 21768 800 21798
rect 1209 21795 1275 21798
rect 4153 21858 4219 21861
rect 4153 21856 4722 21858
rect 4153 21800 4158 21856
rect 4214 21800 4722 21856
rect 4153 21798 4722 21800
rect 4153 21795 4219 21798
rect 3877 21722 3943 21725
rect 4521 21722 4587 21725
rect 3877 21720 4587 21722
rect 3877 21664 3882 21720
rect 3938 21664 4526 21720
rect 4582 21664 4587 21720
rect 3877 21662 4587 21664
rect 4662 21722 4722 21798
rect 5206 21796 5212 21860
rect 5276 21858 5282 21860
rect 5349 21858 5415 21861
rect 5276 21856 5415 21858
rect 5276 21800 5354 21856
rect 5410 21800 5415 21856
rect 5276 21798 5415 21800
rect 5276 21796 5282 21798
rect 5349 21795 5415 21798
rect 6545 21858 6611 21861
rect 8250 21858 8310 21934
rect 10501 21931 10567 21934
rect 13905 21994 13971 21997
rect 14590 21994 14596 21996
rect 13905 21992 14596 21994
rect 13905 21936 13910 21992
rect 13966 21936 14596 21992
rect 13905 21934 14596 21936
rect 13905 21931 13971 21934
rect 14590 21932 14596 21934
rect 14660 21932 14666 21996
rect 15009 21994 15075 21997
rect 20437 21994 20503 21997
rect 15009 21992 20503 21994
rect 15009 21936 15014 21992
rect 15070 21936 20442 21992
rect 20498 21936 20503 21992
rect 15009 21934 20503 21936
rect 15009 21931 15075 21934
rect 20437 21931 20503 21934
rect 21398 21932 21404 21996
rect 21468 21932 21474 21996
rect 23246 21994 23306 22070
rect 23381 22128 23428 22132
rect 23492 22130 23498 22132
rect 24761 22130 24827 22133
rect 25589 22130 25655 22133
rect 23381 22072 23386 22128
rect 23381 22068 23428 22072
rect 23492 22070 23538 22130
rect 24761 22128 25655 22130
rect 24761 22072 24766 22128
rect 24822 22072 25594 22128
rect 25650 22072 25655 22128
rect 24761 22070 25655 22072
rect 23492 22068 23498 22070
rect 23381 22067 23447 22068
rect 24761 22067 24827 22070
rect 25589 22067 25655 22070
rect 24025 21994 24091 21997
rect 23246 21992 24091 21994
rect 23246 21936 24030 21992
rect 24086 21936 24091 21992
rect 23246 21934 24091 21936
rect 6545 21856 8310 21858
rect 6545 21800 6550 21856
rect 6606 21800 8310 21856
rect 6545 21798 8310 21800
rect 8385 21858 8451 21861
rect 9305 21858 9371 21861
rect 8385 21856 9371 21858
rect 8385 21800 8390 21856
rect 8446 21800 9310 21856
rect 9366 21800 9371 21856
rect 8385 21798 9371 21800
rect 6545 21795 6611 21798
rect 8385 21795 8451 21798
rect 9305 21795 9371 21798
rect 10133 21858 10199 21861
rect 11421 21858 11487 21861
rect 10133 21856 11487 21858
rect 10133 21800 10138 21856
rect 10194 21800 11426 21856
rect 11482 21800 11487 21856
rect 10133 21798 11487 21800
rect 10133 21795 10199 21798
rect 11421 21795 11487 21798
rect 17493 21858 17559 21861
rect 17861 21858 17927 21861
rect 18965 21858 19031 21861
rect 17493 21856 17927 21858
rect 17493 21800 17498 21856
rect 17554 21800 17866 21856
rect 17922 21800 17927 21856
rect 17493 21798 17927 21800
rect 17493 21795 17559 21798
rect 17861 21795 17927 21798
rect 18508 21856 19031 21858
rect 18508 21800 18970 21856
rect 19026 21800 19031 21856
rect 18508 21798 19031 21800
rect 18508 21725 18568 21798
rect 18965 21795 19031 21798
rect 19149 21860 19215 21861
rect 19149 21856 19196 21860
rect 19260 21858 19266 21860
rect 20345 21858 20411 21861
rect 21406 21858 21466 21932
rect 24025 21931 24091 21934
rect 25589 21994 25655 21997
rect 26233 21994 26299 21997
rect 25589 21992 26299 21994
rect 25589 21936 25594 21992
rect 25650 21936 26238 21992
rect 26294 21936 26299 21992
rect 25589 21934 26299 21936
rect 25589 21931 25655 21934
rect 26233 21931 26299 21934
rect 19149 21800 19154 21856
rect 19149 21796 19196 21800
rect 19260 21798 19306 21858
rect 20345 21856 21466 21858
rect 20345 21800 20350 21856
rect 20406 21800 21466 21856
rect 20345 21798 21466 21800
rect 22553 21858 22619 21861
rect 22921 21858 22987 21861
rect 22553 21856 22987 21858
rect 22553 21800 22558 21856
rect 22614 21800 22926 21856
rect 22982 21800 22987 21856
rect 22553 21798 22987 21800
rect 19260 21796 19266 21798
rect 19149 21795 19215 21796
rect 20345 21795 20411 21798
rect 22553 21795 22619 21798
rect 22921 21795 22987 21798
rect 23105 21858 23171 21861
rect 24669 21858 24735 21861
rect 23105 21856 24735 21858
rect 23105 21800 23110 21856
rect 23166 21800 24674 21856
rect 24730 21800 24735 21856
rect 23105 21798 24735 21800
rect 23105 21795 23171 21798
rect 24669 21795 24735 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 5533 21722 5599 21725
rect 4662 21720 5599 21722
rect 4662 21664 5538 21720
rect 5594 21664 5599 21720
rect 4662 21662 5599 21664
rect 3877 21659 3943 21662
rect 4521 21659 4587 21662
rect 5533 21659 5599 21662
rect 7925 21722 7991 21725
rect 8569 21722 8635 21725
rect 8937 21722 9003 21725
rect 7925 21720 8172 21722
rect 7925 21664 7930 21720
rect 7986 21664 8172 21720
rect 7925 21662 8172 21664
rect 7925 21659 7991 21662
rect 1945 21586 2011 21589
rect 5625 21586 5691 21589
rect 1945 21584 5691 21586
rect 1945 21528 1950 21584
rect 2006 21528 5630 21584
rect 5686 21528 5691 21584
rect 1945 21526 5691 21528
rect 1945 21523 2011 21526
rect 5625 21523 5691 21526
rect 7005 21586 7071 21589
rect 7925 21586 7991 21589
rect 7005 21584 7991 21586
rect 7005 21528 7010 21584
rect 7066 21528 7930 21584
rect 7986 21528 7991 21584
rect 7005 21526 7991 21528
rect 8112 21586 8172 21662
rect 8569 21720 9003 21722
rect 8569 21664 8574 21720
rect 8630 21664 8942 21720
rect 8998 21664 9003 21720
rect 8569 21662 9003 21664
rect 8569 21659 8635 21662
rect 8937 21659 9003 21662
rect 9765 21722 9831 21725
rect 13629 21722 13695 21725
rect 9765 21720 13695 21722
rect 9765 21664 9770 21720
rect 9826 21664 13634 21720
rect 13690 21664 13695 21720
rect 9765 21662 13695 21664
rect 9765 21659 9831 21662
rect 13629 21659 13695 21662
rect 14917 21722 14983 21725
rect 18505 21722 18571 21725
rect 18965 21724 19031 21725
rect 18965 21722 19012 21724
rect 14917 21720 18571 21722
rect 14917 21664 14922 21720
rect 14978 21664 18510 21720
rect 18566 21664 18571 21720
rect 14917 21662 18571 21664
rect 18920 21720 19012 21722
rect 18920 21664 18970 21720
rect 18920 21662 19012 21664
rect 14917 21659 14983 21662
rect 18505 21659 18571 21662
rect 18965 21660 19012 21662
rect 19076 21660 19082 21724
rect 20253 21722 20319 21725
rect 21633 21722 21699 21725
rect 30189 21722 30255 21725
rect 20253 21720 21699 21722
rect 20253 21664 20258 21720
rect 20314 21664 21638 21720
rect 21694 21664 21699 21720
rect 20253 21662 21699 21664
rect 18965 21659 19074 21660
rect 20253 21659 20319 21662
rect 21633 21659 21699 21662
rect 21774 21720 30255 21722
rect 21774 21664 30194 21720
rect 30250 21664 30255 21720
rect 21774 21662 30255 21664
rect 8937 21586 9003 21589
rect 11513 21586 11579 21589
rect 8112 21584 11579 21586
rect 8112 21528 8942 21584
rect 8998 21528 11518 21584
rect 11574 21528 11579 21584
rect 8112 21526 11579 21528
rect 7005 21523 7071 21526
rect 7925 21523 7991 21526
rect 8937 21523 9003 21526
rect 11513 21523 11579 21526
rect 14958 21524 14964 21588
rect 15028 21586 15034 21588
rect 16573 21586 16639 21589
rect 15028 21584 16639 21586
rect 15028 21528 16578 21584
rect 16634 21528 16639 21584
rect 15028 21526 16639 21528
rect 19014 21586 19074 21659
rect 20294 21586 20300 21588
rect 19014 21526 20300 21586
rect 15028 21524 15034 21526
rect 16573 21523 16639 21526
rect 20294 21524 20300 21526
rect 20364 21524 20370 21588
rect 21081 21586 21147 21589
rect 21214 21586 21220 21588
rect 21081 21584 21220 21586
rect 21081 21528 21086 21584
rect 21142 21528 21220 21584
rect 21081 21526 21220 21528
rect 21081 21523 21147 21526
rect 21214 21524 21220 21526
rect 21284 21586 21290 21588
rect 21774 21586 21834 21662
rect 30189 21659 30255 21662
rect 21284 21526 21834 21586
rect 21909 21586 21975 21589
rect 23933 21586 23999 21589
rect 21909 21584 23999 21586
rect 21909 21528 21914 21584
rect 21970 21528 23938 21584
rect 23994 21528 23999 21584
rect 21909 21526 23999 21528
rect 21284 21524 21290 21526
rect 21909 21523 21975 21526
rect 23933 21523 23999 21526
rect 25313 21586 25379 21589
rect 25773 21586 25839 21589
rect 28533 21586 28599 21589
rect 25313 21584 28599 21586
rect 25313 21528 25318 21584
rect 25374 21528 25778 21584
rect 25834 21528 28538 21584
rect 28594 21528 28599 21584
rect 25313 21526 28599 21528
rect 25313 21523 25379 21526
rect 25773 21523 25839 21526
rect 28533 21523 28599 21526
rect 4245 21450 4311 21453
rect 6545 21450 6611 21453
rect 9397 21450 9463 21453
rect 11053 21450 11119 21453
rect 4245 21448 6611 21450
rect 4245 21392 4250 21448
rect 4306 21392 6550 21448
rect 6606 21392 6611 21448
rect 4245 21390 6611 21392
rect 4245 21387 4311 21390
rect 6545 21387 6611 21390
rect 6686 21448 11119 21450
rect 6686 21392 9402 21448
rect 9458 21392 11058 21448
rect 11114 21392 11119 21448
rect 6686 21390 11119 21392
rect 4889 21314 4955 21317
rect 6269 21314 6335 21317
rect 4889 21312 6335 21314
rect 4889 21256 4894 21312
rect 4950 21256 6274 21312
rect 6330 21256 6335 21312
rect 4889 21254 6335 21256
rect 4889 21251 4955 21254
rect 6269 21251 6335 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 5257 21178 5323 21181
rect 5809 21178 5875 21181
rect 5257 21176 5875 21178
rect 5257 21120 5262 21176
rect 5318 21120 5814 21176
rect 5870 21120 5875 21176
rect 5257 21118 5875 21120
rect 5257 21115 5323 21118
rect 5809 21115 5875 21118
rect 6361 21178 6427 21181
rect 6686 21178 6746 21390
rect 9397 21387 9463 21390
rect 11053 21387 11119 21390
rect 12893 21450 12959 21453
rect 15101 21450 15167 21453
rect 12893 21448 15167 21450
rect 12893 21392 12898 21448
rect 12954 21392 15106 21448
rect 15162 21392 15167 21448
rect 12893 21390 15167 21392
rect 12893 21387 12959 21390
rect 15101 21387 15167 21390
rect 16430 21388 16436 21452
rect 16500 21450 16506 21452
rect 16757 21450 16823 21453
rect 16500 21448 16823 21450
rect 16500 21392 16762 21448
rect 16818 21392 16823 21448
rect 16500 21390 16823 21392
rect 16500 21388 16506 21390
rect 16757 21387 16823 21390
rect 17125 21452 17191 21453
rect 17125 21448 17172 21452
rect 17236 21450 17242 21452
rect 17493 21450 17559 21453
rect 22645 21452 22711 21453
rect 22645 21450 22692 21452
rect 17125 21392 17130 21448
rect 17125 21388 17172 21392
rect 17236 21390 17282 21450
rect 17493 21448 22524 21450
rect 17493 21392 17498 21448
rect 17554 21392 22524 21448
rect 17493 21390 22524 21392
rect 22600 21448 22692 21450
rect 22600 21392 22650 21448
rect 22600 21390 22692 21392
rect 17236 21388 17242 21390
rect 17125 21387 17191 21388
rect 17493 21387 17559 21390
rect 7373 21314 7439 21317
rect 11329 21314 11395 21317
rect 7373 21312 11395 21314
rect 7373 21256 7378 21312
rect 7434 21256 11334 21312
rect 11390 21256 11395 21312
rect 7373 21254 11395 21256
rect 7373 21251 7439 21254
rect 11329 21251 11395 21254
rect 13997 21314 14063 21317
rect 14825 21314 14891 21317
rect 13997 21312 14891 21314
rect 13997 21256 14002 21312
rect 14058 21256 14830 21312
rect 14886 21256 14891 21312
rect 13997 21254 14891 21256
rect 13997 21251 14063 21254
rect 14825 21251 14891 21254
rect 16481 21314 16547 21317
rect 19793 21314 19859 21317
rect 21449 21314 21515 21317
rect 21909 21314 21975 21317
rect 16481 21312 21975 21314
rect 16481 21256 16486 21312
rect 16542 21256 19798 21312
rect 19854 21256 21454 21312
rect 21510 21256 21914 21312
rect 21970 21256 21975 21312
rect 16481 21254 21975 21256
rect 22464 21314 22524 21390
rect 22645 21388 22692 21390
rect 22756 21388 22762 21452
rect 22645 21387 22711 21388
rect 22829 21314 22895 21317
rect 22464 21312 22895 21314
rect 22464 21256 22834 21312
rect 22890 21256 22895 21312
rect 22464 21254 22895 21256
rect 16481 21251 16547 21254
rect 19793 21251 19859 21254
rect 21449 21251 21515 21254
rect 21909 21251 21975 21254
rect 22829 21251 22895 21254
rect 23289 21312 23355 21317
rect 23289 21256 23294 21312
rect 23350 21256 23355 21312
rect 23289 21251 23355 21256
rect 6361 21176 6746 21178
rect 6361 21120 6366 21176
rect 6422 21120 6746 21176
rect 6361 21118 6746 21120
rect 6913 21178 6979 21181
rect 7046 21178 7052 21180
rect 6913 21176 7052 21178
rect 6913 21120 6918 21176
rect 6974 21120 7052 21176
rect 6913 21118 7052 21120
rect 6361 21115 6427 21118
rect 6913 21115 6979 21118
rect 7046 21116 7052 21118
rect 7116 21116 7122 21180
rect 7782 21116 7788 21180
rect 7852 21178 7858 21180
rect 8109 21178 8175 21181
rect 7852 21176 8175 21178
rect 7852 21120 8114 21176
rect 8170 21120 8175 21176
rect 7852 21118 8175 21120
rect 7852 21116 7858 21118
rect 8109 21115 8175 21118
rect 11145 21178 11211 21181
rect 13353 21178 13419 21181
rect 11145 21176 13419 21178
rect 11145 21120 11150 21176
rect 11206 21120 13358 21176
rect 13414 21120 13419 21176
rect 11145 21118 13419 21120
rect 11145 21115 11211 21118
rect 13353 21115 13419 21118
rect 15653 21178 15719 21181
rect 19241 21178 19307 21181
rect 22737 21178 22803 21181
rect 15653 21176 18476 21178
rect 15653 21120 15658 21176
rect 15714 21120 18476 21176
rect 15653 21118 18476 21120
rect 15653 21115 15719 21118
rect 2497 21042 2563 21045
rect 4889 21042 4955 21045
rect 2497 21040 4955 21042
rect 2497 20984 2502 21040
rect 2558 20984 4894 21040
rect 4950 20984 4955 21040
rect 2497 20982 4955 20984
rect 2497 20979 2563 20982
rect 4889 20979 4955 20982
rect 7189 21042 7255 21045
rect 9397 21042 9463 21045
rect 7189 21040 9463 21042
rect 7189 20984 7194 21040
rect 7250 20984 9402 21040
rect 9458 20984 9463 21040
rect 7189 20982 9463 20984
rect 7189 20979 7255 20982
rect 9397 20979 9463 20982
rect 12065 21042 12131 21045
rect 12433 21042 12499 21045
rect 12065 21040 12499 21042
rect 12065 20984 12070 21040
rect 12126 20984 12438 21040
rect 12494 20984 12499 21040
rect 12065 20982 12499 20984
rect 12065 20979 12131 20982
rect 12433 20979 12499 20982
rect 18045 21042 18111 21045
rect 18270 21042 18276 21044
rect 18045 21040 18276 21042
rect 18045 20984 18050 21040
rect 18106 20984 18276 21040
rect 18045 20982 18276 20984
rect 18045 20979 18111 20982
rect 18270 20980 18276 20982
rect 18340 20980 18346 21044
rect 18416 21042 18476 21118
rect 19241 21176 22803 21178
rect 19241 21120 19246 21176
rect 19302 21120 22742 21176
rect 22798 21120 22803 21176
rect 19241 21118 22803 21120
rect 19241 21115 19307 21118
rect 22737 21115 22803 21118
rect 22870 21116 22876 21180
rect 22940 21178 22946 21180
rect 23292 21178 23352 21251
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 22940 21118 23352 21178
rect 22940 21116 22946 21118
rect 19977 21042 20043 21045
rect 20110 21042 20116 21044
rect 18416 21040 20116 21042
rect 18416 20984 19982 21040
rect 20038 20984 20116 21040
rect 18416 20982 20116 20984
rect 3693 20906 3759 20909
rect 7373 20906 7439 20909
rect 8017 20908 8083 20909
rect 3693 20904 7439 20906
rect 3693 20848 3698 20904
rect 3754 20848 7378 20904
rect 7434 20848 7439 20904
rect 3693 20846 7439 20848
rect 3693 20843 3759 20846
rect 7373 20843 7439 20846
rect 7966 20844 7972 20908
rect 8036 20906 8083 20908
rect 8201 20906 8267 20909
rect 8702 20906 8708 20908
rect 8036 20904 8128 20906
rect 8078 20848 8128 20904
rect 8036 20846 8128 20848
rect 8201 20904 8708 20906
rect 8201 20848 8206 20904
rect 8262 20848 8708 20904
rect 8201 20846 8708 20848
rect 8036 20844 8083 20846
rect 7974 20843 8083 20844
rect 8201 20843 8267 20846
rect 8702 20844 8708 20846
rect 8772 20844 8778 20908
rect 10041 20906 10107 20909
rect 15745 20906 15811 20909
rect 10041 20904 15811 20906
rect 10041 20848 10046 20904
rect 10102 20848 15750 20904
rect 15806 20848 15811 20904
rect 10041 20846 15811 20848
rect 10041 20843 10107 20846
rect 15745 20843 15811 20846
rect 16573 20906 16639 20909
rect 17902 20906 17908 20908
rect 16573 20904 17908 20906
rect 16573 20848 16578 20904
rect 16634 20848 17908 20904
rect 16573 20846 17908 20848
rect 16573 20843 16639 20846
rect 17902 20844 17908 20846
rect 17972 20844 17978 20908
rect 18278 20906 18338 20980
rect 19977 20979 20043 20982
rect 20110 20980 20116 20982
rect 20180 20980 20186 21044
rect 20253 21042 20319 21045
rect 20846 21042 20852 21044
rect 20253 21040 20852 21042
rect 20253 20984 20258 21040
rect 20314 20984 20852 21040
rect 20253 20982 20852 20984
rect 20253 20979 20319 20982
rect 20846 20980 20852 20982
rect 20916 21042 20922 21044
rect 21817 21042 21883 21045
rect 20916 21040 21883 21042
rect 20916 20984 21822 21040
rect 21878 20984 21883 21040
rect 20916 20982 21883 20984
rect 20916 20980 20922 20982
rect 21817 20979 21883 20982
rect 23657 21042 23723 21045
rect 25037 21042 25103 21045
rect 26417 21042 26483 21045
rect 23657 21040 26483 21042
rect 23657 20984 23662 21040
rect 23718 20984 25042 21040
rect 25098 20984 26422 21040
rect 26478 20984 26483 21040
rect 23657 20982 26483 20984
rect 23657 20979 23723 20982
rect 25037 20979 25103 20982
rect 26417 20979 26483 20982
rect 18689 20906 18755 20909
rect 19885 20906 19951 20909
rect 22829 20906 22895 20909
rect 23054 20906 23060 20908
rect 18278 20904 18755 20906
rect 18278 20848 18694 20904
rect 18750 20848 18755 20904
rect 18278 20846 18755 20848
rect 18689 20843 18755 20846
rect 19290 20904 21972 20906
rect 19290 20848 19890 20904
rect 19946 20848 21972 20904
rect 19290 20846 21972 20848
rect 0 20770 800 20800
rect 1209 20770 1275 20773
rect 0 20768 1275 20770
rect 0 20712 1214 20768
rect 1270 20712 1275 20768
rect 0 20710 1275 20712
rect 0 20680 800 20710
rect 1209 20707 1275 20710
rect 2497 20770 2563 20773
rect 4705 20770 4771 20773
rect 5574 20770 5580 20772
rect 2497 20768 5580 20770
rect 2497 20712 2502 20768
rect 2558 20712 4710 20768
rect 4766 20712 5580 20768
rect 2497 20710 5580 20712
rect 2497 20707 2563 20710
rect 4705 20707 4771 20710
rect 5574 20708 5580 20710
rect 5644 20708 5650 20772
rect 5758 20708 5764 20772
rect 5828 20770 5834 20772
rect 6177 20770 6243 20773
rect 5828 20768 6243 20770
rect 5828 20712 6182 20768
rect 6238 20712 6243 20768
rect 5828 20710 6243 20712
rect 5828 20708 5834 20710
rect 6177 20707 6243 20710
rect 6821 20770 6887 20773
rect 7189 20770 7255 20773
rect 6821 20768 7255 20770
rect 6821 20712 6826 20768
rect 6882 20712 7194 20768
rect 7250 20712 7255 20768
rect 6821 20710 7255 20712
rect 6821 20707 6887 20710
rect 7189 20707 7255 20710
rect 7557 20772 7623 20773
rect 7557 20768 7604 20772
rect 7668 20770 7674 20772
rect 7557 20712 7562 20768
rect 7557 20708 7604 20712
rect 7668 20710 7714 20770
rect 7668 20708 7674 20710
rect 7557 20707 7623 20708
rect 4153 20634 4219 20637
rect 6545 20634 6611 20637
rect 6678 20634 6684 20636
rect 4153 20632 6684 20634
rect 4153 20576 4158 20632
rect 4214 20576 6550 20632
rect 6606 20576 6684 20632
rect 4153 20574 6684 20576
rect 4153 20571 4219 20574
rect 6545 20571 6611 20574
rect 6678 20572 6684 20574
rect 6748 20572 6754 20636
rect 6821 20634 6887 20637
rect 7974 20634 8034 20843
rect 10777 20770 10843 20773
rect 11053 20772 11119 20773
rect 10910 20770 10916 20772
rect 10777 20768 10916 20770
rect 10777 20712 10782 20768
rect 10838 20712 10916 20768
rect 10777 20710 10916 20712
rect 10777 20707 10843 20710
rect 10910 20708 10916 20710
rect 10980 20708 10986 20772
rect 11053 20768 11100 20772
rect 11164 20770 11170 20772
rect 11053 20712 11058 20768
rect 11053 20708 11100 20712
rect 11164 20710 11210 20770
rect 11164 20708 11170 20710
rect 12750 20708 12756 20772
rect 12820 20770 12826 20772
rect 12893 20770 12959 20773
rect 12820 20768 12959 20770
rect 12820 20712 12898 20768
rect 12954 20712 12959 20768
rect 12820 20710 12959 20712
rect 12820 20708 12826 20710
rect 11053 20707 11119 20708
rect 12893 20707 12959 20710
rect 16573 20770 16639 20773
rect 19290 20770 19350 20846
rect 19885 20843 19951 20846
rect 16573 20768 19350 20770
rect 16573 20712 16578 20768
rect 16634 20712 19350 20768
rect 16573 20710 19350 20712
rect 20161 20770 20227 20773
rect 20662 20770 20668 20772
rect 20161 20768 20668 20770
rect 20161 20712 20166 20768
rect 20222 20712 20668 20768
rect 20161 20710 20668 20712
rect 16573 20707 16639 20710
rect 20161 20707 20227 20710
rect 20662 20708 20668 20710
rect 20732 20708 20738 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 6821 20632 8034 20634
rect 6821 20576 6826 20632
rect 6882 20576 8034 20632
rect 6821 20574 8034 20576
rect 8293 20634 8359 20637
rect 8518 20634 8524 20636
rect 8293 20632 8524 20634
rect 8293 20576 8298 20632
rect 8354 20576 8524 20632
rect 8293 20574 8524 20576
rect 6821 20571 6887 20574
rect 8293 20571 8359 20574
rect 8518 20572 8524 20574
rect 8588 20572 8594 20636
rect 17309 20632 17375 20637
rect 17309 20576 17314 20632
rect 17370 20576 17375 20632
rect 17309 20571 17375 20576
rect 18413 20636 18479 20637
rect 18413 20632 18460 20636
rect 18524 20634 18530 20636
rect 19425 20634 19491 20637
rect 18413 20576 18418 20632
rect 18413 20572 18460 20576
rect 18524 20574 18570 20634
rect 18646 20632 19491 20634
rect 18646 20576 19430 20632
rect 19486 20576 19491 20632
rect 18646 20574 19491 20576
rect 18524 20572 18530 20574
rect 18413 20571 18479 20572
rect 3417 20498 3483 20501
rect 4521 20498 4587 20501
rect 5165 20498 5231 20501
rect 6913 20498 6979 20501
rect 3417 20496 6979 20498
rect 3417 20440 3422 20496
rect 3478 20440 4526 20496
rect 4582 20440 5170 20496
rect 5226 20440 6918 20496
rect 6974 20440 6979 20496
rect 3417 20438 6979 20440
rect 3417 20435 3483 20438
rect 4521 20435 4587 20438
rect 5165 20435 5231 20438
rect 6913 20435 6979 20438
rect 7373 20498 7439 20501
rect 7925 20498 7991 20501
rect 7373 20496 7991 20498
rect 7373 20440 7378 20496
rect 7434 20440 7930 20496
rect 7986 20440 7991 20496
rect 7373 20438 7991 20440
rect 7373 20435 7439 20438
rect 7925 20435 7991 20438
rect 8385 20498 8451 20501
rect 9397 20498 9463 20501
rect 8385 20496 9463 20498
rect 8385 20440 8390 20496
rect 8446 20440 9402 20496
rect 9458 20440 9463 20496
rect 8385 20438 9463 20440
rect 8385 20435 8451 20438
rect 9397 20435 9463 20438
rect 9765 20498 9831 20501
rect 10317 20498 10383 20501
rect 9765 20496 10383 20498
rect 9765 20440 9770 20496
rect 9826 20440 10322 20496
rect 10378 20440 10383 20496
rect 9765 20438 10383 20440
rect 9765 20435 9831 20438
rect 10317 20435 10383 20438
rect 12157 20498 12223 20501
rect 13077 20498 13143 20501
rect 12157 20496 13143 20498
rect 12157 20440 12162 20496
rect 12218 20440 13082 20496
rect 13138 20440 13143 20496
rect 12157 20438 13143 20440
rect 17312 20498 17372 20571
rect 18646 20498 18706 20574
rect 19425 20571 19491 20574
rect 20345 20634 20411 20637
rect 20805 20634 20871 20637
rect 20345 20632 20871 20634
rect 20345 20576 20350 20632
rect 20406 20576 20810 20632
rect 20866 20576 20871 20632
rect 20345 20574 20871 20576
rect 21912 20634 21972 20846
rect 22829 20904 23060 20906
rect 22829 20848 22834 20904
rect 22890 20848 23060 20904
rect 22829 20846 23060 20848
rect 22829 20843 22895 20846
rect 23054 20844 23060 20846
rect 23124 20844 23130 20908
rect 23657 20906 23723 20909
rect 26509 20906 26575 20909
rect 27654 20906 27660 20908
rect 23657 20904 24594 20906
rect 23657 20848 23662 20904
rect 23718 20848 24594 20904
rect 23657 20846 24594 20848
rect 23657 20843 23723 20846
rect 22737 20770 22803 20773
rect 23841 20770 23907 20773
rect 22737 20768 23907 20770
rect 22737 20712 22742 20768
rect 22798 20712 23846 20768
rect 23902 20712 23907 20768
rect 22737 20710 23907 20712
rect 22737 20707 22803 20710
rect 23841 20707 23907 20710
rect 24025 20770 24091 20773
rect 24158 20770 24164 20772
rect 24025 20768 24164 20770
rect 24025 20712 24030 20768
rect 24086 20712 24164 20768
rect 24025 20710 24164 20712
rect 24025 20707 24091 20710
rect 24158 20708 24164 20710
rect 24228 20708 24234 20772
rect 24534 20770 24594 20846
rect 26509 20904 27660 20906
rect 26509 20848 26514 20904
rect 26570 20848 27660 20904
rect 26509 20846 27660 20848
rect 26509 20843 26575 20846
rect 27654 20844 27660 20846
rect 27724 20844 27730 20908
rect 26877 20770 26943 20773
rect 24534 20768 26943 20770
rect 24534 20712 26882 20768
rect 26938 20712 26943 20768
rect 24534 20710 26943 20712
rect 26877 20707 26943 20710
rect 21912 20574 23352 20634
rect 20345 20571 20411 20574
rect 20805 20571 20871 20574
rect 17312 20438 18706 20498
rect 18781 20498 18847 20501
rect 23013 20498 23079 20501
rect 18781 20496 23079 20498
rect 18781 20440 18786 20496
rect 18842 20440 23018 20496
rect 23074 20440 23079 20496
rect 18781 20438 23079 20440
rect 12157 20435 12223 20438
rect 13077 20435 13143 20438
rect 18781 20435 18847 20438
rect 23013 20435 23079 20438
rect 3049 20362 3115 20365
rect 8477 20362 8543 20365
rect 3049 20360 8543 20362
rect 3049 20304 3054 20360
rect 3110 20304 8482 20360
rect 8538 20304 8543 20360
rect 3049 20302 8543 20304
rect 3049 20299 3115 20302
rect 8477 20299 8543 20302
rect 10869 20362 10935 20365
rect 13169 20362 13235 20365
rect 14825 20362 14891 20365
rect 10869 20360 14891 20362
rect 10869 20304 10874 20360
rect 10930 20304 13174 20360
rect 13230 20304 14830 20360
rect 14886 20304 14891 20360
rect 10869 20302 14891 20304
rect 10869 20299 10935 20302
rect 13169 20299 13235 20302
rect 14825 20299 14891 20302
rect 17718 20300 17724 20364
rect 17788 20362 17794 20364
rect 19977 20362 20043 20365
rect 23292 20362 23352 20574
rect 23422 20572 23428 20636
rect 23492 20634 23498 20636
rect 23933 20634 23999 20637
rect 23492 20632 23999 20634
rect 23492 20576 23938 20632
rect 23994 20576 23999 20632
rect 23492 20574 23999 20576
rect 23492 20572 23498 20574
rect 23933 20571 23999 20574
rect 26366 20572 26372 20636
rect 26436 20634 26442 20636
rect 26601 20634 26667 20637
rect 26436 20632 26667 20634
rect 26436 20576 26606 20632
rect 26662 20576 26667 20632
rect 26436 20574 26667 20576
rect 26436 20572 26442 20574
rect 26601 20571 26667 20574
rect 24025 20498 24091 20501
rect 24342 20498 24348 20500
rect 24025 20496 24348 20498
rect 24025 20440 24030 20496
rect 24086 20440 24348 20496
rect 24025 20438 24348 20440
rect 24025 20435 24091 20438
rect 24342 20436 24348 20438
rect 24412 20436 24418 20500
rect 27153 20498 27219 20501
rect 28257 20498 28323 20501
rect 27153 20496 28323 20498
rect 27153 20440 27158 20496
rect 27214 20440 28262 20496
rect 28318 20440 28323 20496
rect 27153 20438 28323 20440
rect 27153 20435 27219 20438
rect 28257 20435 28323 20438
rect 24209 20362 24275 20365
rect 17788 20360 20043 20362
rect 17788 20304 19982 20360
rect 20038 20304 20043 20360
rect 17788 20302 20043 20304
rect 17788 20300 17794 20302
rect 19977 20299 20043 20302
rect 20118 20302 22110 20362
rect 23292 20360 24275 20362
rect 23292 20304 24214 20360
rect 24270 20304 24275 20360
rect 23292 20302 24275 20304
rect 4889 20226 4955 20229
rect 8702 20226 8708 20228
rect 4889 20224 8708 20226
rect 4889 20168 4894 20224
rect 4950 20168 8708 20224
rect 4889 20166 8708 20168
rect 4889 20163 4955 20166
rect 8702 20164 8708 20166
rect 8772 20164 8778 20228
rect 9305 20226 9371 20229
rect 10685 20226 10751 20229
rect 11145 20226 11211 20229
rect 9305 20224 11211 20226
rect 9305 20168 9310 20224
rect 9366 20168 10690 20224
rect 10746 20168 11150 20224
rect 11206 20168 11211 20224
rect 9305 20166 11211 20168
rect 9305 20163 9371 20166
rect 10685 20163 10751 20166
rect 11145 20163 11211 20166
rect 11881 20226 11947 20229
rect 12985 20226 13051 20229
rect 11881 20224 13051 20226
rect 11881 20168 11886 20224
rect 11942 20168 12990 20224
rect 13046 20168 13051 20224
rect 11881 20166 13051 20168
rect 11881 20163 11947 20166
rect 12985 20163 13051 20166
rect 19241 20226 19307 20229
rect 20118 20226 20178 20302
rect 19241 20224 20178 20226
rect 19241 20168 19246 20224
rect 19302 20168 20178 20224
rect 19241 20166 20178 20168
rect 19241 20163 19307 20166
rect 20294 20164 20300 20228
rect 20364 20226 20370 20228
rect 21081 20226 21147 20229
rect 20364 20224 21147 20226
rect 20364 20168 21086 20224
rect 21142 20168 21147 20224
rect 20364 20166 21147 20168
rect 22050 20226 22110 20302
rect 24209 20299 24275 20302
rect 26233 20362 26299 20365
rect 26233 20360 28136 20362
rect 26233 20304 26238 20360
rect 26294 20304 28136 20360
rect 26233 20302 28136 20304
rect 26233 20299 26299 20302
rect 28076 20229 28136 20302
rect 25129 20226 25195 20229
rect 27838 20226 27844 20228
rect 22050 20224 27844 20226
rect 22050 20168 25134 20224
rect 25190 20168 27844 20224
rect 22050 20166 27844 20168
rect 20364 20164 20370 20166
rect 21081 20163 21147 20166
rect 25129 20163 25195 20166
rect 27838 20164 27844 20166
rect 27908 20164 27914 20228
rect 28073 20224 28139 20229
rect 28073 20168 28078 20224
rect 28134 20168 28139 20224
rect 28073 20163 28139 20168
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 5022 20028 5028 20092
rect 5092 20028 5098 20092
rect 5257 20090 5323 20093
rect 7649 20090 7715 20093
rect 8201 20092 8267 20093
rect 8150 20090 8156 20092
rect 5257 20088 7715 20090
rect 5257 20032 5262 20088
rect 5318 20032 7654 20088
rect 7710 20032 7715 20088
rect 5257 20030 7715 20032
rect 8110 20030 8156 20090
rect 8220 20088 8267 20092
rect 8262 20032 8267 20088
rect 5030 19957 5090 20028
rect 5257 20027 5323 20030
rect 7649 20027 7715 20030
rect 8150 20028 8156 20030
rect 8220 20028 8267 20032
rect 8201 20027 8267 20028
rect 10409 20090 10475 20093
rect 10869 20090 10935 20093
rect 12341 20090 12407 20093
rect 10409 20088 12407 20090
rect 10409 20032 10414 20088
rect 10470 20032 10874 20088
rect 10930 20032 12346 20088
rect 12402 20032 12407 20088
rect 10409 20030 12407 20032
rect 10409 20027 10475 20030
rect 10869 20027 10935 20030
rect 12341 20027 12407 20030
rect 14457 20090 14523 20093
rect 22461 20090 22527 20093
rect 14457 20088 22527 20090
rect 14457 20032 14462 20088
rect 14518 20032 22466 20088
rect 22522 20032 22527 20088
rect 14457 20030 22527 20032
rect 14457 20027 14523 20030
rect 22461 20027 22527 20030
rect 23289 20090 23355 20093
rect 27337 20090 27403 20093
rect 23289 20088 27403 20090
rect 23289 20032 23294 20088
rect 23350 20032 27342 20088
rect 27398 20032 27403 20088
rect 23289 20030 27403 20032
rect 23289 20027 23355 20030
rect 27337 20027 27403 20030
rect 4981 19952 5090 19957
rect 4981 19896 4986 19952
rect 5042 19896 5090 19952
rect 4981 19894 5090 19896
rect 5257 19954 5323 19957
rect 5901 19954 5967 19957
rect 5257 19952 5967 19954
rect 5257 19896 5262 19952
rect 5318 19896 5906 19952
rect 5962 19896 5967 19952
rect 5257 19894 5967 19896
rect 4981 19891 5047 19894
rect 5257 19891 5323 19894
rect 5901 19891 5967 19894
rect 6177 19954 6243 19957
rect 7741 19954 7807 19957
rect 6177 19952 7807 19954
rect 6177 19896 6182 19952
rect 6238 19896 7746 19952
rect 7802 19896 7807 19952
rect 6177 19894 7807 19896
rect 6177 19891 6243 19894
rect 7741 19891 7807 19894
rect 11329 19954 11395 19957
rect 14089 19954 14155 19957
rect 11329 19952 14155 19954
rect 11329 19896 11334 19952
rect 11390 19896 14094 19952
rect 14150 19896 14155 19952
rect 11329 19894 14155 19896
rect 11329 19891 11395 19894
rect 14089 19891 14155 19894
rect 16389 19954 16455 19957
rect 18321 19954 18387 19957
rect 22870 19954 22876 19956
rect 16389 19952 22876 19954
rect 16389 19896 16394 19952
rect 16450 19896 18326 19952
rect 18382 19896 22876 19952
rect 16389 19894 22876 19896
rect 16389 19891 16455 19894
rect 18321 19891 18387 19894
rect 22870 19892 22876 19894
rect 22940 19954 22946 19956
rect 24577 19954 24643 19957
rect 22940 19952 24643 19954
rect 22940 19896 24582 19952
rect 24638 19896 24643 19952
rect 22940 19894 24643 19896
rect 22940 19892 22946 19894
rect 24577 19891 24643 19894
rect 4245 19818 4311 19821
rect 4613 19818 4679 19821
rect 5257 19818 5323 19821
rect 6361 19820 6427 19821
rect 4245 19816 5323 19818
rect 4245 19760 4250 19816
rect 4306 19760 4618 19816
rect 4674 19760 5262 19816
rect 5318 19760 5323 19816
rect 4245 19758 5323 19760
rect 4245 19755 4311 19758
rect 4613 19755 4679 19758
rect 5257 19755 5323 19758
rect 6310 19756 6316 19820
rect 6380 19818 6427 19820
rect 7465 19818 7531 19821
rect 7598 19818 7604 19820
rect 6380 19816 6472 19818
rect 6422 19760 6472 19816
rect 6380 19758 6472 19760
rect 7465 19816 7604 19818
rect 7465 19760 7470 19816
rect 7526 19760 7604 19816
rect 7465 19758 7604 19760
rect 6380 19756 6427 19758
rect 6361 19755 6427 19756
rect 7465 19755 7531 19758
rect 7598 19756 7604 19758
rect 7668 19756 7674 19820
rect 7741 19818 7807 19821
rect 8753 19818 8819 19821
rect 7741 19816 8819 19818
rect 7741 19760 7746 19816
rect 7802 19760 8758 19816
rect 8814 19760 8819 19816
rect 7741 19758 8819 19760
rect 7741 19755 7807 19758
rect 8753 19755 8819 19758
rect 13302 19756 13308 19820
rect 13372 19818 13378 19820
rect 13537 19818 13603 19821
rect 13372 19816 13603 19818
rect 13372 19760 13542 19816
rect 13598 19760 13603 19816
rect 13372 19758 13603 19760
rect 13372 19756 13378 19758
rect 13537 19755 13603 19758
rect 15510 19756 15516 19820
rect 15580 19818 15586 19820
rect 15653 19818 15719 19821
rect 15580 19816 15719 19818
rect 15580 19760 15658 19816
rect 15714 19760 15719 19816
rect 15580 19758 15719 19760
rect 15580 19756 15586 19758
rect 15653 19755 15719 19758
rect 17902 19756 17908 19820
rect 17972 19818 17978 19820
rect 18965 19818 19031 19821
rect 19701 19818 19767 19821
rect 17972 19816 19031 19818
rect 17972 19760 18970 19816
rect 19026 19760 19031 19816
rect 17972 19758 19031 19760
rect 17972 19756 17978 19758
rect 18965 19755 19031 19758
rect 19382 19816 19767 19818
rect 19382 19760 19706 19816
rect 19762 19760 19767 19816
rect 19382 19758 19767 19760
rect 0 19682 800 19712
rect 1209 19682 1275 19685
rect 0 19680 1275 19682
rect 0 19624 1214 19680
rect 1270 19624 1275 19680
rect 0 19622 1275 19624
rect 0 19592 800 19622
rect 1209 19619 1275 19622
rect 3918 19620 3924 19684
rect 3988 19620 3994 19684
rect 4061 19682 4127 19685
rect 9581 19682 9647 19685
rect 12065 19682 12131 19685
rect 4061 19680 9647 19682
rect 4061 19624 4066 19680
rect 4122 19624 9586 19680
rect 9642 19624 9647 19680
rect 4061 19622 9647 19624
rect 3926 19546 3986 19620
rect 4061 19619 4127 19622
rect 9581 19619 9647 19622
rect 9998 19680 12131 19682
rect 9998 19624 12070 19680
rect 12126 19624 12131 19680
rect 9998 19622 12131 19624
rect 4521 19546 4587 19549
rect 3926 19544 4587 19546
rect 3926 19488 4526 19544
rect 4582 19488 4587 19544
rect 3926 19486 4587 19488
rect 4521 19483 4587 19486
rect 5165 19546 5231 19549
rect 7281 19546 7347 19549
rect 5165 19544 7347 19546
rect 5165 19488 5170 19544
rect 5226 19488 7286 19544
rect 7342 19488 7347 19544
rect 5165 19486 7347 19488
rect 5165 19483 5231 19486
rect 7281 19483 7347 19486
rect 7782 19484 7788 19548
rect 7852 19546 7858 19548
rect 8109 19546 8175 19549
rect 9998 19548 10058 19622
rect 12065 19619 12131 19622
rect 18597 19682 18663 19685
rect 19382 19682 19442 19758
rect 19701 19755 19767 19758
rect 23105 19818 23171 19821
rect 23565 19818 23631 19821
rect 23105 19816 23631 19818
rect 23105 19760 23110 19816
rect 23166 19760 23570 19816
rect 23626 19760 23631 19816
rect 23105 19758 23631 19760
rect 23105 19755 23171 19758
rect 23565 19755 23631 19758
rect 27337 19818 27403 19821
rect 29637 19818 29703 19821
rect 27337 19816 29703 19818
rect 27337 19760 27342 19816
rect 27398 19760 29642 19816
rect 29698 19760 29703 19816
rect 27337 19758 29703 19760
rect 27337 19755 27403 19758
rect 29637 19755 29703 19758
rect 18597 19680 19442 19682
rect 18597 19624 18602 19680
rect 18658 19624 19442 19680
rect 18597 19622 19442 19624
rect 21449 19682 21515 19685
rect 22001 19682 22067 19685
rect 21449 19680 22067 19682
rect 21449 19624 21454 19680
rect 21510 19624 22006 19680
rect 22062 19624 22067 19680
rect 21449 19622 22067 19624
rect 18597 19619 18663 19622
rect 21449 19619 21515 19622
rect 22001 19619 22067 19622
rect 22921 19682 22987 19685
rect 25957 19682 26023 19685
rect 22921 19680 26023 19682
rect 22921 19624 22926 19680
rect 22982 19624 25962 19680
rect 26018 19624 26023 19680
rect 22921 19622 26023 19624
rect 22921 19619 22987 19622
rect 25957 19619 26023 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 9990 19546 9996 19548
rect 7852 19544 8175 19546
rect 7852 19488 8114 19544
rect 8170 19488 8175 19544
rect 7852 19486 8175 19488
rect 7852 19484 7858 19486
rect 8109 19483 8175 19486
rect 9630 19486 9996 19546
rect 4981 19410 5047 19413
rect 6862 19410 6868 19412
rect 4981 19408 6868 19410
rect 4981 19352 4986 19408
rect 5042 19352 6868 19408
rect 4981 19350 6868 19352
rect 4981 19347 5047 19350
rect 6862 19348 6868 19350
rect 6932 19410 6938 19412
rect 7373 19410 7439 19413
rect 6932 19408 7439 19410
rect 6932 19352 7378 19408
rect 7434 19352 7439 19408
rect 6932 19350 7439 19352
rect 6932 19348 6938 19350
rect 7373 19347 7439 19350
rect 3049 19274 3115 19277
rect 9630 19274 9690 19486
rect 9990 19484 9996 19486
rect 10060 19484 10066 19548
rect 14181 19546 14247 19549
rect 11976 19544 14247 19546
rect 11976 19488 14186 19544
rect 14242 19488 14247 19544
rect 11976 19486 14247 19488
rect 11976 19413 12036 19486
rect 14181 19483 14247 19486
rect 11830 19348 11836 19412
rect 11900 19410 11906 19412
rect 11973 19410 12039 19413
rect 11900 19408 12039 19410
rect 11900 19352 11978 19408
rect 12034 19352 12039 19408
rect 11900 19350 12039 19352
rect 11900 19348 11906 19350
rect 11973 19347 12039 19350
rect 15142 19348 15148 19412
rect 15212 19410 15218 19412
rect 19885 19410 19951 19413
rect 20478 19410 20484 19412
rect 15212 19408 20484 19410
rect 15212 19352 19890 19408
rect 19946 19352 20484 19408
rect 15212 19350 20484 19352
rect 15212 19348 15218 19350
rect 19885 19347 19951 19350
rect 20478 19348 20484 19350
rect 20548 19348 20554 19412
rect 21582 19410 21588 19412
rect 20670 19350 21588 19410
rect 3049 19272 9690 19274
rect 3049 19216 3054 19272
rect 3110 19216 9690 19272
rect 3049 19214 9690 19216
rect 15377 19274 15443 19277
rect 17309 19276 17375 19277
rect 17585 19276 17651 19277
rect 16982 19274 16988 19276
rect 15377 19272 16988 19274
rect 15377 19216 15382 19272
rect 15438 19216 16988 19272
rect 15377 19214 16988 19216
rect 3049 19211 3115 19214
rect 15377 19211 15443 19214
rect 16982 19212 16988 19214
rect 17052 19212 17058 19276
rect 17309 19274 17356 19276
rect 17264 19272 17356 19274
rect 17264 19216 17314 19272
rect 17264 19214 17356 19216
rect 17309 19212 17356 19214
rect 17420 19212 17426 19276
rect 17534 19212 17540 19276
rect 17604 19274 17651 19276
rect 18045 19274 18111 19277
rect 20345 19274 20411 19277
rect 17604 19272 17696 19274
rect 17646 19216 17696 19272
rect 17604 19214 17696 19216
rect 18045 19272 20411 19274
rect 18045 19216 18050 19272
rect 18106 19216 20350 19272
rect 20406 19216 20411 19272
rect 18045 19214 20411 19216
rect 17604 19212 17651 19214
rect 17309 19211 17375 19212
rect 17585 19211 17651 19212
rect 18045 19211 18111 19214
rect 20345 19211 20411 19214
rect 6085 19138 6151 19141
rect 6913 19138 6979 19141
rect 6085 19136 6979 19138
rect 6085 19080 6090 19136
rect 6146 19080 6918 19136
rect 6974 19080 6979 19136
rect 6085 19078 6979 19080
rect 6085 19075 6151 19078
rect 6913 19075 6979 19078
rect 7189 19138 7255 19141
rect 11053 19138 11119 19141
rect 7189 19136 11119 19138
rect 7189 19080 7194 19136
rect 7250 19080 11058 19136
rect 11114 19080 11119 19136
rect 7189 19078 11119 19080
rect 7189 19075 7255 19078
rect 11053 19075 11119 19078
rect 15101 19138 15167 19141
rect 20670 19138 20730 19350
rect 21582 19348 21588 19350
rect 21652 19410 21658 19412
rect 21909 19410 21975 19413
rect 21652 19408 21975 19410
rect 21652 19352 21914 19408
rect 21970 19352 21975 19408
rect 21652 19350 21975 19352
rect 21652 19348 21658 19350
rect 21909 19347 21975 19350
rect 23289 19276 23355 19277
rect 23238 19212 23244 19276
rect 23308 19274 23355 19276
rect 23308 19272 23400 19274
rect 23350 19216 23400 19272
rect 23308 19214 23400 19216
rect 23308 19212 23355 19214
rect 23289 19211 23355 19212
rect 15101 19136 20730 19138
rect 15101 19080 15106 19136
rect 15162 19080 20730 19136
rect 15101 19078 20730 19080
rect 21449 19138 21515 19141
rect 26233 19138 26299 19141
rect 21449 19136 26299 19138
rect 21449 19080 21454 19136
rect 21510 19080 26238 19136
rect 26294 19080 26299 19136
rect 21449 19078 26299 19080
rect 15101 19075 15167 19078
rect 21449 19075 21515 19078
rect 26233 19075 26299 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 8385 19002 8451 19005
rect 10869 19002 10935 19005
rect 8385 19000 10935 19002
rect 8385 18944 8390 19000
rect 8446 18944 10874 19000
rect 10930 18944 10935 19000
rect 8385 18942 10935 18944
rect 8385 18939 8451 18942
rect 10869 18939 10935 18942
rect 13721 19002 13787 19005
rect 16113 19002 16179 19005
rect 13721 19000 16179 19002
rect 13721 18944 13726 19000
rect 13782 18944 16118 19000
rect 16174 18944 16179 19000
rect 13721 18942 16179 18944
rect 13721 18939 13787 18942
rect 16113 18939 16179 18942
rect 18413 19002 18479 19005
rect 20805 19002 20871 19005
rect 21357 19002 21423 19005
rect 22277 19002 22343 19005
rect 18413 19000 21423 19002
rect 18413 18944 18418 19000
rect 18474 18944 20810 19000
rect 20866 18944 21362 19000
rect 21418 18944 21423 19000
rect 18413 18942 21423 18944
rect 18413 18939 18479 18942
rect 20805 18939 20871 18942
rect 21357 18939 21423 18942
rect 21590 19000 22343 19002
rect 21590 18944 22282 19000
rect 22338 18944 22343 19000
rect 21590 18942 22343 18944
rect 3509 18866 3575 18869
rect 9857 18866 9923 18869
rect 3509 18864 9923 18866
rect 3509 18808 3514 18864
rect 3570 18808 9862 18864
rect 9918 18808 9923 18864
rect 3509 18806 9923 18808
rect 3509 18803 3575 18806
rect 9857 18803 9923 18806
rect 10777 18866 10843 18869
rect 14273 18866 14339 18869
rect 10777 18864 14339 18866
rect 10777 18808 10782 18864
rect 10838 18808 14278 18864
rect 14334 18808 14339 18864
rect 10777 18806 14339 18808
rect 10777 18803 10843 18806
rect 14273 18803 14339 18806
rect 16113 18866 16179 18869
rect 16757 18866 16823 18869
rect 16113 18864 16823 18866
rect 16113 18808 16118 18864
rect 16174 18808 16762 18864
rect 16818 18808 16823 18864
rect 16113 18806 16823 18808
rect 16113 18803 16179 18806
rect 16757 18803 16823 18806
rect 19701 18866 19767 18869
rect 21590 18866 21650 18942
rect 22277 18939 22343 18942
rect 24393 19002 24459 19005
rect 25957 19002 26023 19005
rect 29085 19002 29151 19005
rect 24393 19000 29151 19002
rect 24393 18944 24398 19000
rect 24454 18944 25962 19000
rect 26018 18944 29090 19000
rect 29146 18944 29151 19000
rect 24393 18942 29151 18944
rect 24393 18939 24459 18942
rect 25957 18939 26023 18942
rect 29085 18939 29151 18942
rect 19701 18864 21650 18866
rect 19701 18808 19706 18864
rect 19762 18808 21650 18864
rect 19701 18806 21650 18808
rect 21725 18866 21791 18869
rect 25129 18866 25195 18869
rect 21725 18864 25195 18866
rect 21725 18808 21730 18864
rect 21786 18808 25134 18864
rect 25190 18808 25195 18864
rect 21725 18806 25195 18808
rect 19701 18803 19767 18806
rect 21725 18803 21791 18806
rect 25129 18803 25195 18806
rect 6126 18668 6132 18732
rect 6196 18730 6202 18732
rect 6269 18730 6335 18733
rect 6196 18728 6335 18730
rect 6196 18672 6274 18728
rect 6330 18672 6335 18728
rect 6196 18670 6335 18672
rect 6196 18668 6202 18670
rect 6269 18667 6335 18670
rect 10501 18730 10567 18733
rect 12617 18730 12683 18733
rect 21357 18730 21423 18733
rect 22093 18730 22159 18733
rect 25497 18730 25563 18733
rect 27102 18730 27108 18732
rect 10501 18728 12683 18730
rect 10501 18672 10506 18728
rect 10562 18672 12622 18728
rect 12678 18672 12683 18728
rect 10501 18670 12683 18672
rect 10501 18667 10567 18670
rect 12617 18667 12683 18670
rect 18416 18670 20362 18730
rect 0 18594 800 18624
rect 18416 18597 18476 18670
rect 1209 18594 1275 18597
rect 0 18592 1275 18594
rect 0 18536 1214 18592
rect 1270 18536 1275 18592
rect 0 18534 1275 18536
rect 0 18504 800 18534
rect 1209 18531 1275 18534
rect 8385 18594 8451 18597
rect 9121 18594 9187 18597
rect 8385 18592 9187 18594
rect 8385 18536 8390 18592
rect 8446 18536 9126 18592
rect 9182 18536 9187 18592
rect 8385 18534 9187 18536
rect 8385 18531 8451 18534
rect 9121 18531 9187 18534
rect 18413 18592 18479 18597
rect 18413 18536 18418 18592
rect 18474 18536 18479 18592
rect 18413 18531 18479 18536
rect 20302 18594 20362 18670
rect 21357 18728 22159 18730
rect 21357 18672 21362 18728
rect 21418 18672 22098 18728
rect 22154 18672 22159 18728
rect 21357 18670 22159 18672
rect 21357 18667 21423 18670
rect 22093 18667 22159 18670
rect 24902 18728 27108 18730
rect 24902 18672 25502 18728
rect 25558 18672 27108 18728
rect 24902 18670 27108 18672
rect 21030 18594 21036 18596
rect 20302 18534 21036 18594
rect 21030 18532 21036 18534
rect 21100 18594 21106 18596
rect 22185 18594 22251 18597
rect 23289 18594 23355 18597
rect 21100 18534 22110 18594
rect 21100 18532 21106 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 3601 18458 3667 18461
rect 11094 18458 11100 18460
rect 3601 18456 11100 18458
rect 3601 18400 3606 18456
rect 3662 18400 11100 18456
rect 3601 18398 11100 18400
rect 3601 18395 3667 18398
rect 11094 18396 11100 18398
rect 11164 18396 11170 18460
rect 14549 18458 14615 18461
rect 16021 18458 16087 18461
rect 14549 18456 16087 18458
rect 14549 18400 14554 18456
rect 14610 18400 16026 18456
rect 16082 18400 16087 18456
rect 14549 18398 16087 18400
rect 14549 18395 14615 18398
rect 16021 18395 16087 18398
rect 16481 18458 16547 18461
rect 18781 18458 18847 18461
rect 16481 18456 18847 18458
rect 16481 18400 16486 18456
rect 16542 18400 18786 18456
rect 18842 18400 18847 18456
rect 16481 18398 18847 18400
rect 22050 18458 22110 18534
rect 22185 18592 23355 18594
rect 22185 18536 22190 18592
rect 22246 18536 23294 18592
rect 23350 18536 23355 18592
rect 22185 18534 23355 18536
rect 22185 18531 22251 18534
rect 23289 18531 23355 18534
rect 24902 18458 24962 18670
rect 25497 18667 25563 18670
rect 27102 18668 27108 18670
rect 27172 18668 27178 18732
rect 22050 18398 24962 18458
rect 16481 18395 16547 18398
rect 18781 18395 18847 18398
rect 6545 18322 6611 18325
rect 7281 18322 7347 18325
rect 13813 18322 13879 18325
rect 14273 18322 14339 18325
rect 6545 18320 7666 18322
rect 6545 18264 6550 18320
rect 6606 18264 7286 18320
rect 7342 18264 7666 18320
rect 6545 18262 7666 18264
rect 6545 18259 6611 18262
rect 7281 18259 7347 18262
rect 7606 18186 7666 18262
rect 13813 18320 14339 18322
rect 13813 18264 13818 18320
rect 13874 18264 14278 18320
rect 14334 18264 14339 18320
rect 13813 18262 14339 18264
rect 13813 18259 13879 18262
rect 14273 18259 14339 18262
rect 15285 18322 15351 18325
rect 17585 18322 17651 18325
rect 24117 18322 24183 18325
rect 24761 18322 24827 18325
rect 15285 18320 15394 18322
rect 15285 18264 15290 18320
rect 15346 18264 15394 18320
rect 15285 18259 15394 18264
rect 17585 18320 24827 18322
rect 17585 18264 17590 18320
rect 17646 18264 24122 18320
rect 24178 18264 24766 18320
rect 24822 18264 24827 18320
rect 17585 18262 24827 18264
rect 17585 18259 17651 18262
rect 24117 18259 24183 18262
rect 24761 18259 24827 18262
rect 9581 18186 9647 18189
rect 7606 18184 9647 18186
rect 7606 18128 9586 18184
rect 9642 18128 9647 18184
rect 7606 18126 9647 18128
rect 9581 18123 9647 18126
rect 13445 18186 13511 18189
rect 14641 18186 14707 18189
rect 15193 18188 15259 18189
rect 15142 18186 15148 18188
rect 13445 18184 14707 18186
rect 13445 18128 13450 18184
rect 13506 18128 14646 18184
rect 14702 18128 14707 18184
rect 13445 18126 14707 18128
rect 15102 18126 15148 18186
rect 15212 18184 15259 18188
rect 15254 18128 15259 18184
rect 13445 18123 13511 18126
rect 14641 18123 14707 18126
rect 15142 18124 15148 18126
rect 15212 18124 15259 18128
rect 15334 18186 15394 18259
rect 16389 18186 16455 18189
rect 22829 18186 22895 18189
rect 15334 18184 22895 18186
rect 15334 18128 16394 18184
rect 16450 18128 22834 18184
rect 22890 18128 22895 18184
rect 15334 18126 22895 18128
rect 15193 18123 15259 18124
rect 16389 18123 16455 18126
rect 22829 18123 22895 18126
rect 7097 18050 7163 18053
rect 7741 18050 7807 18053
rect 7097 18048 7807 18050
rect 7097 17992 7102 18048
rect 7158 17992 7746 18048
rect 7802 17992 7807 18048
rect 7097 17990 7807 17992
rect 7097 17987 7163 17990
rect 7741 17987 7807 17990
rect 8385 18050 8451 18053
rect 9121 18050 9187 18053
rect 8385 18048 9187 18050
rect 8385 17992 8390 18048
rect 8446 17992 9126 18048
rect 9182 17992 9187 18048
rect 8385 17990 9187 17992
rect 8385 17987 8451 17990
rect 9121 17987 9187 17990
rect 13670 17988 13676 18052
rect 13740 18050 13746 18052
rect 17401 18050 17467 18053
rect 13740 18048 17467 18050
rect 13740 17992 17406 18048
rect 17462 17992 17467 18048
rect 13740 17990 17467 17992
rect 13740 17988 13746 17990
rect 17401 17987 17467 17990
rect 22001 18050 22067 18053
rect 23841 18050 23907 18053
rect 22001 18048 23907 18050
rect 22001 17992 22006 18048
rect 22062 17992 23846 18048
rect 23902 17992 23907 18048
rect 22001 17990 23907 17992
rect 22001 17987 22067 17990
rect 23841 17987 23907 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 7189 17916 7255 17917
rect 7189 17914 7236 17916
rect 7144 17912 7236 17914
rect 7144 17856 7194 17912
rect 7144 17854 7236 17856
rect 7189 17852 7236 17854
rect 7300 17852 7306 17916
rect 8201 17914 8267 17917
rect 8334 17914 8340 17916
rect 8201 17912 8340 17914
rect 8201 17856 8206 17912
rect 8262 17856 8340 17912
rect 8201 17854 8340 17856
rect 7189 17851 7255 17852
rect 8201 17851 8267 17854
rect 8334 17852 8340 17854
rect 8404 17852 8410 17916
rect 10961 17914 11027 17917
rect 12750 17914 12756 17916
rect 10961 17912 12756 17914
rect 10961 17856 10966 17912
rect 11022 17856 12756 17912
rect 10961 17854 12756 17856
rect 10961 17851 11027 17854
rect 12750 17852 12756 17854
rect 12820 17852 12826 17916
rect 13169 17914 13235 17917
rect 16297 17914 16363 17917
rect 13169 17912 16363 17914
rect 13169 17856 13174 17912
rect 13230 17856 16302 17912
rect 16358 17856 16363 17912
rect 13169 17854 16363 17856
rect 13169 17851 13235 17854
rect 16297 17851 16363 17854
rect 19517 17914 19583 17917
rect 20529 17914 20595 17917
rect 21817 17914 21883 17917
rect 19517 17912 21883 17914
rect 19517 17856 19522 17912
rect 19578 17856 20534 17912
rect 20590 17856 21822 17912
rect 21878 17856 21883 17912
rect 19517 17854 21883 17856
rect 19517 17851 19583 17854
rect 20529 17851 20595 17854
rect 21817 17851 21883 17854
rect 22185 17914 22251 17917
rect 24158 17914 24164 17916
rect 22185 17912 24164 17914
rect 22185 17856 22190 17912
rect 22246 17856 24164 17912
rect 22185 17854 24164 17856
rect 22185 17851 22251 17854
rect 24158 17852 24164 17854
rect 24228 17914 24234 17916
rect 25681 17914 25747 17917
rect 24228 17912 25747 17914
rect 24228 17856 25686 17912
rect 25742 17856 25747 17912
rect 24228 17854 25747 17856
rect 24228 17852 24234 17854
rect 25681 17851 25747 17854
rect 4061 17778 4127 17781
rect 9622 17778 9628 17780
rect 4061 17776 9628 17778
rect 4061 17720 4066 17776
rect 4122 17720 9628 17776
rect 4061 17718 9628 17720
rect 4061 17715 4127 17718
rect 9622 17716 9628 17718
rect 9692 17716 9698 17780
rect 12617 17778 12683 17781
rect 14825 17778 14891 17781
rect 12617 17776 14891 17778
rect 12617 17720 12622 17776
rect 12678 17720 14830 17776
rect 14886 17720 14891 17776
rect 12617 17718 14891 17720
rect 12617 17715 12683 17718
rect 14825 17715 14891 17718
rect 15285 17778 15351 17781
rect 17585 17778 17651 17781
rect 15285 17776 17651 17778
rect 15285 17720 15290 17776
rect 15346 17720 17590 17776
rect 17646 17720 17651 17776
rect 15285 17718 17651 17720
rect 15285 17715 15351 17718
rect 17585 17715 17651 17718
rect 21081 17778 21147 17781
rect 26693 17778 26759 17781
rect 21081 17776 26759 17778
rect 21081 17720 21086 17776
rect 21142 17720 26698 17776
rect 26754 17720 26759 17776
rect 21081 17718 26759 17720
rect 21081 17715 21147 17718
rect 26693 17715 26759 17718
rect 5717 17642 5783 17645
rect 7005 17642 7071 17645
rect 5717 17640 7071 17642
rect 5717 17584 5722 17640
rect 5778 17584 7010 17640
rect 7066 17584 7071 17640
rect 5717 17582 7071 17584
rect 5717 17579 5783 17582
rect 7005 17579 7071 17582
rect 13629 17642 13695 17645
rect 16205 17642 16271 17645
rect 16849 17642 16915 17645
rect 13629 17640 16915 17642
rect 13629 17584 13634 17640
rect 13690 17584 16210 17640
rect 16266 17584 16854 17640
rect 16910 17584 16915 17640
rect 13629 17582 16915 17584
rect 13629 17579 13695 17582
rect 16205 17579 16271 17582
rect 16849 17579 16915 17582
rect 18413 17642 18479 17645
rect 20161 17642 20227 17645
rect 20897 17642 20963 17645
rect 18413 17640 20963 17642
rect 18413 17584 18418 17640
rect 18474 17584 20166 17640
rect 20222 17584 20902 17640
rect 20958 17584 20963 17640
rect 18413 17582 20963 17584
rect 18413 17579 18479 17582
rect 20161 17579 20227 17582
rect 20897 17579 20963 17582
rect 21357 17642 21423 17645
rect 23657 17642 23723 17645
rect 21357 17640 23723 17642
rect 21357 17584 21362 17640
rect 21418 17584 23662 17640
rect 23718 17584 23723 17640
rect 21357 17582 23723 17584
rect 21357 17579 21423 17582
rect 23657 17579 23723 17582
rect 0 17506 800 17536
rect 1209 17506 1275 17509
rect 0 17504 1275 17506
rect 0 17448 1214 17504
rect 1270 17448 1275 17504
rect 0 17446 1275 17448
rect 0 17416 800 17446
rect 1209 17443 1275 17446
rect 7046 17444 7052 17508
rect 7116 17506 7122 17508
rect 7281 17506 7347 17509
rect 7116 17504 7347 17506
rect 7116 17448 7286 17504
rect 7342 17448 7347 17504
rect 7116 17446 7347 17448
rect 7116 17444 7122 17446
rect 7281 17443 7347 17446
rect 21449 17506 21515 17509
rect 25589 17506 25655 17509
rect 21449 17504 25655 17506
rect 21449 17448 21454 17504
rect 21510 17448 25594 17504
rect 25650 17448 25655 17504
rect 21449 17446 25655 17448
rect 21449 17443 21515 17446
rect 25589 17443 25655 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 13445 17370 13511 17373
rect 17309 17370 17375 17373
rect 13445 17368 17375 17370
rect 13445 17312 13450 17368
rect 13506 17312 17314 17368
rect 17370 17312 17375 17368
rect 13445 17310 17375 17312
rect 13445 17307 13511 17310
rect 17309 17307 17375 17310
rect 13629 17234 13695 17237
rect 13997 17234 14063 17237
rect 15101 17234 15167 17237
rect 13629 17232 15167 17234
rect 13629 17176 13634 17232
rect 13690 17176 14002 17232
rect 14058 17176 15106 17232
rect 15162 17176 15167 17232
rect 13629 17174 15167 17176
rect 13629 17171 13695 17174
rect 13997 17171 14063 17174
rect 15101 17171 15167 17174
rect 19885 17234 19951 17237
rect 21357 17234 21423 17237
rect 19885 17232 21423 17234
rect 19885 17176 19890 17232
rect 19946 17176 21362 17232
rect 21418 17176 21423 17232
rect 19885 17174 21423 17176
rect 19885 17171 19951 17174
rect 21357 17171 21423 17174
rect 21633 17234 21699 17237
rect 23565 17234 23631 17237
rect 21633 17232 23631 17234
rect 21633 17176 21638 17232
rect 21694 17176 23570 17232
rect 23626 17176 23631 17232
rect 21633 17174 23631 17176
rect 21633 17171 21699 17174
rect 23565 17171 23631 17174
rect 5758 17036 5764 17100
rect 5828 17098 5834 17100
rect 5993 17098 6059 17101
rect 5828 17096 6059 17098
rect 5828 17040 5998 17096
rect 6054 17040 6059 17096
rect 5828 17038 6059 17040
rect 5828 17036 5834 17038
rect 5993 17035 6059 17038
rect 13537 17098 13603 17101
rect 15745 17098 15811 17101
rect 13537 17096 15811 17098
rect 13537 17040 13542 17096
rect 13598 17040 15750 17096
rect 15806 17040 15811 17096
rect 13537 17038 15811 17040
rect 13537 17035 13603 17038
rect 15745 17035 15811 17038
rect 5901 16964 5967 16965
rect 5901 16962 5948 16964
rect 5856 16960 5948 16962
rect 5856 16904 5906 16960
rect 5856 16902 5948 16904
rect 5901 16900 5948 16902
rect 6012 16900 6018 16964
rect 15009 16962 15075 16965
rect 16573 16962 16639 16965
rect 15009 16960 16639 16962
rect 15009 16904 15014 16960
rect 15070 16904 16578 16960
rect 16634 16904 16639 16960
rect 15009 16902 16639 16904
rect 5901 16899 5967 16900
rect 15009 16899 15075 16902
rect 16573 16899 16639 16902
rect 43161 16962 43227 16965
rect 44200 16962 45000 16992
rect 43161 16960 45000 16962
rect 43161 16904 43166 16960
rect 43222 16904 45000 16960
rect 43161 16902 45000 16904
rect 43161 16899 43227 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 44200 16872 45000 16902
rect 34930 16831 35246 16832
rect 7649 16690 7715 16693
rect 11697 16690 11763 16693
rect 7649 16688 11763 16690
rect 7649 16632 7654 16688
rect 7710 16632 11702 16688
rect 11758 16632 11763 16688
rect 7649 16630 11763 16632
rect 7649 16627 7715 16630
rect 11697 16627 11763 16630
rect 12065 16690 12131 16693
rect 14181 16690 14247 16693
rect 12065 16688 14247 16690
rect 12065 16632 12070 16688
rect 12126 16632 14186 16688
rect 14242 16632 14247 16688
rect 12065 16630 14247 16632
rect 12065 16627 12131 16630
rect 14181 16627 14247 16630
rect 7373 16556 7439 16557
rect 7373 16554 7420 16556
rect 7328 16552 7420 16554
rect 7328 16496 7378 16552
rect 7328 16494 7420 16496
rect 7373 16492 7420 16494
rect 7484 16492 7490 16556
rect 12157 16554 12223 16557
rect 13813 16556 13879 16557
rect 12566 16554 12572 16556
rect 12157 16552 12572 16554
rect 12157 16496 12162 16552
rect 12218 16496 12572 16552
rect 12157 16494 12572 16496
rect 7373 16491 7439 16492
rect 12157 16491 12223 16494
rect 12566 16492 12572 16494
rect 12636 16492 12642 16556
rect 13813 16554 13860 16556
rect 13768 16552 13860 16554
rect 13768 16496 13818 16552
rect 13768 16494 13860 16496
rect 13813 16492 13860 16494
rect 13924 16492 13930 16556
rect 14406 16492 14412 16556
rect 14476 16554 14482 16556
rect 15377 16554 15443 16557
rect 14476 16552 15443 16554
rect 14476 16496 15382 16552
rect 15438 16496 15443 16552
rect 14476 16494 15443 16496
rect 14476 16492 14482 16494
rect 13813 16491 13879 16492
rect 15377 16491 15443 16494
rect 18505 16554 18571 16557
rect 18638 16554 18644 16556
rect 18505 16552 18644 16554
rect 18505 16496 18510 16552
rect 18566 16496 18644 16552
rect 18505 16494 18644 16496
rect 18505 16491 18571 16494
rect 18638 16492 18644 16494
rect 18708 16492 18714 16556
rect 20662 16492 20668 16556
rect 20732 16554 20738 16556
rect 22553 16554 22619 16557
rect 20732 16552 22619 16554
rect 20732 16496 22558 16552
rect 22614 16496 22619 16552
rect 20732 16494 22619 16496
rect 20732 16492 20738 16494
rect 22553 16491 22619 16494
rect 0 16418 800 16448
rect 1209 16418 1275 16421
rect 0 16416 1275 16418
rect 0 16360 1214 16416
rect 1270 16360 1275 16416
rect 0 16358 1275 16360
rect 0 16328 800 16358
rect 1209 16355 1275 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4061 16146 4127 16149
rect 6453 16146 6519 16149
rect 13302 16146 13308 16148
rect 4061 16144 13308 16146
rect 4061 16088 4066 16144
rect 4122 16088 6458 16144
rect 6514 16088 13308 16144
rect 4061 16086 13308 16088
rect 4061 16083 4127 16086
rect 6453 16083 6519 16086
rect 13302 16084 13308 16086
rect 13372 16084 13378 16148
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 13169 15602 13235 15605
rect 15009 15602 15075 15605
rect 13169 15600 15075 15602
rect 13169 15544 13174 15600
rect 13230 15544 15014 15600
rect 15070 15544 15075 15600
rect 13169 15542 15075 15544
rect 13169 15539 13235 15542
rect 15009 15539 15075 15542
rect 0 15330 800 15360
rect 1209 15330 1275 15333
rect 0 15328 1275 15330
rect 0 15272 1214 15328
rect 1270 15272 1275 15328
rect 0 15270 1275 15272
rect 0 15240 800 15270
rect 1209 15267 1275 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 7833 15194 7899 15197
rect 8518 15194 8524 15196
rect 7833 15192 8524 15194
rect 7833 15136 7838 15192
rect 7894 15136 8524 15192
rect 7833 15134 8524 15136
rect 7833 15131 7899 15134
rect 8518 15132 8524 15134
rect 8588 15132 8594 15196
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14242 800 14272
rect 1209 14242 1275 14245
rect 0 14240 1275 14242
rect 0 14184 1214 14240
rect 1270 14184 1275 14240
rect 0 14182 1275 14184
rect 0 14152 800 14182
rect 1209 14179 1275 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13154 800 13184
rect 1209 13154 1275 13157
rect 0 13152 1275 13154
rect 0 13096 1214 13152
rect 1270 13096 1275 13152
rect 0 13094 1275 13096
rect 0 13064 800 13094
rect 1209 13091 1275 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12066 800 12096
rect 1209 12066 1275 12069
rect 0 12064 1275 12066
rect 0 12008 1214 12064
rect 1270 12008 1275 12064
rect 0 12006 1275 12008
rect 0 11976 800 12006
rect 1209 12003 1275 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 9890 800 9920
rect 1209 9890 1275 9893
rect 0 9888 1275 9890
rect 0 9832 1214 9888
rect 1270 9832 1275 9888
rect 0 9830 1275 9832
rect 0 9800 800 9830
rect 1209 9827 1275 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 3141 8938 3207 8941
rect 12014 8938 12020 8940
rect 3141 8936 12020 8938
rect 3141 8880 3146 8936
rect 3202 8880 12020 8936
rect 3141 8878 12020 8880
rect 3141 8875 3207 8878
rect 12014 8876 12020 8878
rect 12084 8876 12090 8940
rect 0 8802 800 8832
rect 1209 8802 1275 8805
rect 0 8800 1275 8802
rect 0 8744 1214 8800
rect 1270 8744 1275 8800
rect 0 8742 1275 8744
rect 0 8712 800 8742
rect 1209 8739 1275 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 0 7714 800 7744
rect 1209 7714 1275 7717
rect 0 7712 1275 7714
rect 0 7656 1214 7712
rect 1270 7656 1275 7712
rect 0 7654 1275 7656
rect 0 7624 800 7654
rect 1209 7651 1275 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6626 800 6656
rect 1209 6626 1275 6629
rect 0 6624 1275 6626
rect 0 6568 1214 6624
rect 1270 6568 1275 6624
rect 0 6566 1275 6568
rect 0 6536 800 6566
rect 1209 6563 1275 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 40677 5810 40743 5813
rect 44200 5810 45000 5840
rect 40677 5808 45000 5810
rect 40677 5752 40682 5808
rect 40738 5752 45000 5808
rect 40677 5750 45000 5752
rect 40677 5747 40743 5750
rect 44200 5720 45000 5750
rect 0 5538 800 5568
rect 1853 5538 1919 5541
rect 0 5536 1919 5538
rect 0 5480 1858 5536
rect 1914 5480 1919 5536
rect 0 5478 1919 5480
rect 0 5448 800 5478
rect 1853 5475 1919 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 0 4450 800 4480
rect 1209 4450 1275 4453
rect 0 4448 1275 4450
rect 0 4392 1214 4448
rect 1270 4392 1275 4448
rect 0 4390 1275 4392
rect 0 4360 800 4390
rect 1209 4387 1275 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 3141 4044 3207 4045
rect 3141 4042 3188 4044
rect 3096 4040 3188 4042
rect 3096 3984 3146 4040
rect 3096 3982 3188 3984
rect 3141 3980 3188 3982
rect 3252 3980 3258 4044
rect 3141 3979 3207 3980
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3362 800 3392
rect 1209 3362 1275 3365
rect 0 3360 1275 3362
rect 0 3304 1214 3360
rect 1270 3304 1275 3360
rect 0 3302 1275 3304
rect 0 3272 800 3302
rect 1209 3299 1275 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 24669 2682 24735 2685
rect 24894 2682 24900 2684
rect 24669 2680 24900 2682
rect 24669 2624 24674 2680
rect 24730 2624 24900 2680
rect 24669 2622 24900 2624
rect 24669 2619 24735 2622
rect 24894 2620 24900 2622
rect 24964 2620 24970 2684
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 10364 38388 10428 38452
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 8340 35940 8404 36004
rect 25636 35940 25700 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 9444 35124 9508 35188
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 8156 34716 8220 34780
rect 11468 34580 11532 34644
rect 11836 34444 11900 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 25452 34172 25516 34236
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 26372 33492 26436 33556
rect 24900 33416 24964 33420
rect 24900 33360 24950 33416
rect 24950 33360 24964 33416
rect 24900 33356 24964 33360
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 27660 33084 27724 33148
rect 18460 32736 18524 32740
rect 18460 32680 18510 32736
rect 18510 32680 18524 32736
rect 18460 32676 18524 32680
rect 28580 32676 28644 32740
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 6132 31996 6196 32060
rect 25820 31996 25884 32060
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 25268 31452 25332 31516
rect 18092 31316 18156 31380
rect 25452 31044 25516 31108
rect 25820 31044 25884 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 26188 30908 26252 30972
rect 21036 30772 21100 30836
rect 9628 30500 9692 30564
rect 16436 30500 16500 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 26556 30500 26620 30564
rect 5212 30424 5276 30428
rect 5212 30368 5226 30424
rect 5226 30368 5276 30424
rect 5212 30364 5276 30368
rect 10916 30364 10980 30428
rect 14596 30364 14660 30428
rect 14964 30364 15028 30428
rect 26372 30364 26436 30428
rect 25268 30092 25332 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 17908 29140 17972 29204
rect 23244 29004 23308 29068
rect 9260 28868 9324 28932
rect 9628 28868 9692 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 8156 28732 8220 28796
rect 16252 28732 16316 28796
rect 26556 28868 26620 28932
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 24900 28732 24964 28796
rect 27660 28384 27724 28388
rect 27660 28328 27710 28384
rect 27710 28328 27724 28384
rect 27660 28324 27724 28328
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 7052 28052 7116 28116
rect 5580 27916 5644 27980
rect 16620 27916 16684 27980
rect 7604 27780 7668 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 17908 27508 17972 27572
rect 13860 27236 13924 27300
rect 14596 27236 14660 27300
rect 25636 27508 25700 27572
rect 26188 27236 26252 27300
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 8340 27160 8404 27164
rect 8340 27104 8354 27160
rect 8354 27104 8404 27160
rect 8340 27100 8404 27104
rect 26924 27100 26988 27164
rect 6500 26828 6564 26892
rect 13676 26692 13740 26756
rect 20668 26692 20732 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 16436 26616 16500 26620
rect 16436 26560 16450 26616
rect 16450 26560 16500 26616
rect 16436 26556 16500 26560
rect 17356 26344 17420 26348
rect 17356 26288 17370 26344
rect 17370 26288 17420 26344
rect 17356 26284 17420 26288
rect 20300 26148 20364 26212
rect 27660 26284 27724 26348
rect 25268 26148 25332 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 9444 26012 9508 26076
rect 16436 26012 16500 26076
rect 24164 26012 24228 26076
rect 7972 25876 8036 25940
rect 26372 25740 26436 25804
rect 6868 25604 6932 25668
rect 7236 25604 7300 25668
rect 11836 25664 11900 25668
rect 11836 25608 11886 25664
rect 11886 25608 11900 25664
rect 11836 25604 11900 25608
rect 26556 25604 26620 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 9260 25332 9324 25396
rect 11468 25392 11532 25396
rect 11468 25336 11518 25392
rect 11518 25336 11532 25392
rect 11468 25332 11532 25336
rect 16620 25332 16684 25396
rect 20300 25332 20364 25396
rect 26924 25468 26988 25532
rect 7236 25120 7300 25124
rect 7236 25064 7250 25120
rect 7250 25064 7300 25120
rect 7236 25060 7300 25064
rect 16252 25196 16316 25260
rect 17540 25256 17604 25260
rect 17540 25200 17554 25256
rect 17554 25200 17604 25256
rect 17540 25196 17604 25200
rect 23060 25196 23124 25260
rect 15516 25060 15580 25124
rect 20116 25120 20180 25124
rect 20116 25064 20166 25120
rect 20166 25064 20180 25120
rect 20116 25060 20180 25064
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 6684 24924 6748 24988
rect 14412 24924 14476 24988
rect 17172 24984 17236 24988
rect 17172 24928 17222 24984
rect 17222 24928 17236 24984
rect 17172 24924 17236 24928
rect 20300 24924 20364 24988
rect 20484 24984 20548 24988
rect 20484 24928 20498 24984
rect 20498 24928 20548 24984
rect 20484 24924 20548 24928
rect 21404 24924 21468 24988
rect 5580 24788 5644 24852
rect 7052 24788 7116 24852
rect 7604 24712 7668 24716
rect 7604 24656 7654 24712
rect 7654 24656 7668 24712
rect 7604 24652 7668 24656
rect 19012 24712 19076 24716
rect 19012 24656 19026 24712
rect 19026 24656 19076 24712
rect 19012 24652 19076 24656
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 5580 24168 5644 24172
rect 5580 24112 5594 24168
rect 5594 24112 5644 24168
rect 5580 24108 5644 24112
rect 20852 24108 20916 24172
rect 6500 23972 6564 24036
rect 8156 24032 8220 24036
rect 8156 23976 8206 24032
rect 8206 23976 8220 24032
rect 8156 23972 8220 23976
rect 19196 23972 19260 24036
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 22692 23972 22756 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 5396 23836 5460 23900
rect 6868 23836 6932 23900
rect 19380 23896 19444 23900
rect 19380 23840 19430 23896
rect 19430 23840 19444 23896
rect 19380 23836 19444 23840
rect 21220 23896 21284 23900
rect 21220 23840 21234 23896
rect 21234 23840 21284 23896
rect 21220 23836 21284 23840
rect 26556 23836 26620 23900
rect 3188 23700 3252 23764
rect 24348 23700 24412 23764
rect 6132 23564 6196 23628
rect 12020 23624 12084 23628
rect 12020 23568 12070 23624
rect 12070 23568 12084 23624
rect 12020 23564 12084 23568
rect 5028 23428 5092 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 6132 23292 6196 23356
rect 7236 23292 7300 23356
rect 17724 23488 17788 23492
rect 17724 23432 17738 23488
rect 17738 23432 17788 23488
rect 17724 23428 17788 23432
rect 27108 23488 27172 23492
rect 27108 23432 27158 23488
rect 27158 23432 27172 23488
rect 27108 23428 27172 23432
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 20668 23292 20732 23356
rect 6868 23080 6932 23084
rect 6868 23024 6918 23080
rect 6918 23024 6932 23080
rect 6868 23020 6932 23024
rect 9628 23020 9692 23084
rect 16436 23020 16500 23084
rect 16988 23020 17052 23084
rect 28580 23080 28644 23084
rect 28580 23024 28594 23080
rect 28594 23024 28644 23080
rect 28580 23020 28644 23024
rect 3924 22748 3988 22812
rect 5212 22884 5276 22948
rect 10364 22884 10428 22948
rect 18092 22884 18156 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 11836 22748 11900 22812
rect 18276 22748 18340 22812
rect 6316 22476 6380 22540
rect 7420 22476 7484 22540
rect 9260 22476 9324 22540
rect 12572 22536 12636 22540
rect 12572 22480 12586 22536
rect 12586 22480 12636 22536
rect 12572 22476 12636 22480
rect 19380 22612 19444 22676
rect 27844 22476 27908 22540
rect 5396 22340 5460 22404
rect 5948 22400 6012 22404
rect 5948 22344 5962 22400
rect 5962 22344 6012 22400
rect 5948 22340 6012 22344
rect 15148 22340 15212 22404
rect 18644 22340 18708 22404
rect 20116 22400 20180 22404
rect 20116 22344 20130 22400
rect 20130 22344 20180 22400
rect 20116 22340 20180 22344
rect 21588 22400 21652 22404
rect 21588 22344 21602 22400
rect 21602 22344 21652 22400
rect 21588 22340 21652 22344
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 8340 22264 8404 22268
rect 8340 22208 8354 22264
rect 8354 22208 8404 22264
rect 8340 22204 8404 22208
rect 5580 22068 5644 22132
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 9996 22068 10060 22132
rect 20300 22068 20364 22132
rect 5028 21992 5092 21996
rect 5028 21936 5042 21992
rect 5042 21936 5092 21992
rect 5028 21932 5092 21936
rect 5212 21796 5276 21860
rect 14596 21932 14660 21996
rect 21404 21932 21468 21996
rect 23428 22128 23492 22132
rect 23428 22072 23442 22128
rect 23442 22072 23492 22128
rect 23428 22068 23492 22072
rect 19196 21856 19260 21860
rect 19196 21800 19210 21856
rect 19210 21800 19260 21856
rect 19196 21796 19260 21800
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 19012 21720 19076 21724
rect 19012 21664 19026 21720
rect 19026 21664 19076 21720
rect 19012 21660 19076 21664
rect 14964 21524 15028 21588
rect 20300 21524 20364 21588
rect 21220 21524 21284 21588
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 16436 21388 16500 21452
rect 17172 21448 17236 21452
rect 17172 21392 17186 21448
rect 17186 21392 17236 21448
rect 17172 21388 17236 21392
rect 22692 21448 22756 21452
rect 22692 21392 22706 21448
rect 22706 21392 22756 21448
rect 22692 21388 22756 21392
rect 7052 21116 7116 21180
rect 7788 21116 7852 21180
rect 18276 20980 18340 21044
rect 22876 21116 22940 21180
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 7972 20904 8036 20908
rect 7972 20848 8022 20904
rect 8022 20848 8036 20904
rect 7972 20844 8036 20848
rect 8708 20844 8772 20908
rect 17908 20844 17972 20908
rect 20116 20980 20180 21044
rect 20852 20980 20916 21044
rect 5580 20708 5644 20772
rect 5764 20708 5828 20772
rect 7604 20768 7668 20772
rect 7604 20712 7618 20768
rect 7618 20712 7668 20768
rect 7604 20708 7668 20712
rect 6684 20572 6748 20636
rect 10916 20708 10980 20772
rect 11100 20768 11164 20772
rect 11100 20712 11114 20768
rect 11114 20712 11164 20768
rect 11100 20708 11164 20712
rect 12756 20708 12820 20772
rect 20668 20708 20732 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 8524 20572 8588 20636
rect 18460 20632 18524 20636
rect 18460 20576 18474 20632
rect 18474 20576 18524 20632
rect 18460 20572 18524 20576
rect 23060 20844 23124 20908
rect 24164 20708 24228 20772
rect 27660 20844 27724 20908
rect 17724 20300 17788 20364
rect 23428 20572 23492 20636
rect 26372 20572 26436 20636
rect 24348 20436 24412 20500
rect 8708 20164 8772 20228
rect 20300 20164 20364 20228
rect 27844 20164 27908 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 5028 20028 5092 20092
rect 8156 20088 8220 20092
rect 8156 20032 8206 20088
rect 8206 20032 8220 20088
rect 8156 20028 8220 20032
rect 22876 19892 22940 19956
rect 6316 19816 6380 19820
rect 6316 19760 6366 19816
rect 6366 19760 6380 19816
rect 6316 19756 6380 19760
rect 7604 19756 7668 19820
rect 13308 19756 13372 19820
rect 15516 19756 15580 19820
rect 17908 19756 17972 19820
rect 3924 19620 3988 19684
rect 7788 19484 7852 19548
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 6868 19348 6932 19412
rect 9996 19484 10060 19548
rect 11836 19348 11900 19412
rect 15148 19348 15212 19412
rect 20484 19348 20548 19412
rect 16988 19212 17052 19276
rect 17356 19272 17420 19276
rect 17356 19216 17370 19272
rect 17370 19216 17420 19272
rect 17356 19212 17420 19216
rect 17540 19272 17604 19276
rect 17540 19216 17590 19272
rect 17590 19216 17604 19272
rect 17540 19212 17604 19216
rect 21588 19348 21652 19412
rect 23244 19272 23308 19276
rect 23244 19216 23294 19272
rect 23294 19216 23308 19272
rect 23244 19212 23308 19216
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 6132 18668 6196 18732
rect 21036 18532 21100 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 11100 18396 11164 18460
rect 27108 18668 27172 18732
rect 15148 18184 15212 18188
rect 15148 18128 15198 18184
rect 15198 18128 15212 18184
rect 15148 18124 15212 18128
rect 13676 17988 13740 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 7236 17912 7300 17916
rect 7236 17856 7250 17912
rect 7250 17856 7300 17912
rect 7236 17852 7300 17856
rect 8340 17852 8404 17916
rect 12756 17852 12820 17916
rect 24164 17852 24228 17916
rect 9628 17716 9692 17780
rect 7052 17444 7116 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 5764 17036 5828 17100
rect 5948 16960 6012 16964
rect 5948 16904 5962 16960
rect 5962 16904 6012 16960
rect 5948 16900 6012 16904
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 7420 16552 7484 16556
rect 7420 16496 7434 16552
rect 7434 16496 7484 16552
rect 7420 16492 7484 16496
rect 12572 16492 12636 16556
rect 13860 16552 13924 16556
rect 13860 16496 13874 16552
rect 13874 16496 13924 16552
rect 13860 16492 13924 16496
rect 14412 16492 14476 16556
rect 18644 16492 18708 16556
rect 20668 16492 20732 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 13308 16084 13372 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 8524 15132 8588 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 12020 8876 12084 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 3188 4040 3252 4044
rect 3188 3984 3202 4040
rect 3202 3984 3252 4040
rect 3188 3980 3252 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 24900 2620 24964 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 41920 4528 42480
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 19568 42464 19888 42480
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 10363 38452 10429 38453
rect 10363 38388 10364 38452
rect 10428 38388 10429 38452
rect 10363 38387 10429 38388
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 8339 36004 8405 36005
rect 8339 35940 8340 36004
rect 8404 35940 8405 36004
rect 8339 35939 8405 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 8155 34780 8221 34781
rect 8155 34716 8156 34780
rect 8220 34716 8221 34780
rect 8155 34715 8221 34716
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 6131 32060 6197 32061
rect 6131 31996 6132 32060
rect 6196 31996 6197 32060
rect 6131 31995 6197 31996
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 5211 30428 5277 30429
rect 5211 30364 5212 30428
rect 5276 30364 5277 30428
rect 5211 30363 5277 30364
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3187 23764 3253 23765
rect 3187 23700 3188 23764
rect 3252 23700 3253 23764
rect 3187 23699 3253 23700
rect 3190 4045 3250 23699
rect 4208 23424 4528 24448
rect 5027 23492 5093 23493
rect 5027 23428 5028 23492
rect 5092 23428 5093 23492
rect 5027 23427 5093 23428
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 3923 22812 3989 22813
rect 3923 22748 3924 22812
rect 3988 22748 3989 22812
rect 3923 22747 3989 22748
rect 3926 19685 3986 22747
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 5030 21997 5090 23427
rect 5214 22949 5274 30363
rect 5579 27980 5645 27981
rect 5579 27916 5580 27980
rect 5644 27916 5645 27980
rect 5579 27915 5645 27916
rect 5582 24853 5642 27915
rect 5579 24852 5645 24853
rect 5579 24788 5580 24852
rect 5644 24788 5645 24852
rect 5579 24787 5645 24788
rect 5579 24172 5645 24173
rect 5579 24108 5580 24172
rect 5644 24108 5645 24172
rect 5579 24107 5645 24108
rect 5395 23900 5461 23901
rect 5395 23836 5396 23900
rect 5460 23836 5461 23900
rect 5395 23835 5461 23836
rect 5211 22948 5277 22949
rect 5211 22884 5212 22948
rect 5276 22884 5277 22948
rect 5211 22883 5277 22884
rect 5027 21996 5093 21997
rect 5027 21932 5028 21996
rect 5092 21932 5093 21996
rect 5027 21931 5093 21932
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3923 19684 3989 19685
rect 3923 19620 3924 19684
rect 3988 19620 3989 19684
rect 3923 19619 3989 19620
rect 4208 19072 4528 20096
rect 5030 20093 5090 21931
rect 5214 21861 5274 22883
rect 5398 22405 5458 23835
rect 5395 22404 5461 22405
rect 5395 22340 5396 22404
rect 5460 22340 5461 22404
rect 5395 22339 5461 22340
rect 5582 22133 5642 24107
rect 6134 23629 6194 31995
rect 8158 28797 8218 34715
rect 8155 28796 8221 28797
rect 8155 28732 8156 28796
rect 8220 28732 8221 28796
rect 8155 28731 8221 28732
rect 7051 28116 7117 28117
rect 7051 28052 7052 28116
rect 7116 28052 7117 28116
rect 7051 28051 7117 28052
rect 6499 26892 6565 26893
rect 6499 26828 6500 26892
rect 6564 26828 6565 26892
rect 6499 26827 6565 26828
rect 6502 24037 6562 26827
rect 6867 25668 6933 25669
rect 6867 25604 6868 25668
rect 6932 25604 6933 25668
rect 6867 25603 6933 25604
rect 6683 24988 6749 24989
rect 6683 24924 6684 24988
rect 6748 24924 6749 24988
rect 6683 24923 6749 24924
rect 6499 24036 6565 24037
rect 6499 23972 6500 24036
rect 6564 23972 6565 24036
rect 6499 23971 6565 23972
rect 6131 23628 6197 23629
rect 6131 23564 6132 23628
rect 6196 23564 6197 23628
rect 6131 23563 6197 23564
rect 6131 23356 6197 23357
rect 6131 23292 6132 23356
rect 6196 23292 6197 23356
rect 6131 23291 6197 23292
rect 5947 22404 6013 22405
rect 5947 22340 5948 22404
rect 6012 22340 6013 22404
rect 5947 22339 6013 22340
rect 5579 22132 5645 22133
rect 5579 22068 5580 22132
rect 5644 22068 5645 22132
rect 5579 22067 5645 22068
rect 5211 21860 5277 21861
rect 5211 21796 5212 21860
rect 5276 21796 5277 21860
rect 5211 21795 5277 21796
rect 5582 20773 5642 22067
rect 5579 20772 5645 20773
rect 5579 20708 5580 20772
rect 5644 20708 5645 20772
rect 5579 20707 5645 20708
rect 5763 20772 5829 20773
rect 5763 20708 5764 20772
rect 5828 20708 5829 20772
rect 5763 20707 5829 20708
rect 5027 20092 5093 20093
rect 5027 20028 5028 20092
rect 5092 20028 5093 20092
rect 5027 20027 5093 20028
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 5766 17101 5826 20707
rect 5763 17100 5829 17101
rect 5763 17036 5764 17100
rect 5828 17036 5829 17100
rect 5763 17035 5829 17036
rect 5950 16965 6010 22339
rect 6134 18733 6194 23291
rect 6315 22540 6381 22541
rect 6315 22476 6316 22540
rect 6380 22476 6381 22540
rect 6315 22475 6381 22476
rect 6318 19821 6378 22475
rect 6686 20637 6746 24923
rect 6870 23901 6930 25603
rect 7054 24853 7114 28051
rect 7603 27844 7669 27845
rect 7603 27780 7604 27844
rect 7668 27780 7669 27844
rect 7603 27779 7669 27780
rect 7235 25668 7301 25669
rect 7235 25604 7236 25668
rect 7300 25604 7301 25668
rect 7235 25603 7301 25604
rect 7238 25125 7298 25603
rect 7235 25124 7301 25125
rect 7235 25060 7236 25124
rect 7300 25060 7301 25124
rect 7235 25059 7301 25060
rect 7051 24852 7117 24853
rect 7051 24788 7052 24852
rect 7116 24788 7117 24852
rect 7051 24787 7117 24788
rect 7606 24717 7666 27779
rect 8342 27165 8402 35939
rect 9443 35188 9509 35189
rect 9443 35124 9444 35188
rect 9508 35124 9509 35188
rect 9443 35123 9509 35124
rect 9259 28932 9325 28933
rect 9259 28868 9260 28932
rect 9324 28868 9325 28932
rect 9259 28867 9325 28868
rect 8339 27164 8405 27165
rect 8339 27100 8340 27164
rect 8404 27100 8405 27164
rect 8339 27099 8405 27100
rect 7971 25940 8037 25941
rect 7971 25876 7972 25940
rect 8036 25876 8037 25940
rect 7971 25875 8037 25876
rect 7603 24716 7669 24717
rect 7603 24652 7604 24716
rect 7668 24652 7669 24716
rect 7603 24651 7669 24652
rect 6867 23900 6933 23901
rect 6867 23836 6868 23900
rect 6932 23836 6933 23900
rect 6867 23835 6933 23836
rect 7235 23356 7301 23357
rect 7235 23292 7236 23356
rect 7300 23292 7301 23356
rect 7235 23291 7301 23292
rect 6867 23084 6933 23085
rect 6867 23020 6868 23084
rect 6932 23020 6933 23084
rect 6867 23019 6933 23020
rect 6683 20636 6749 20637
rect 6683 20572 6684 20636
rect 6748 20572 6749 20636
rect 6683 20571 6749 20572
rect 6315 19820 6381 19821
rect 6315 19756 6316 19820
rect 6380 19756 6381 19820
rect 6315 19755 6381 19756
rect 6870 19413 6930 23019
rect 7051 21180 7117 21181
rect 7051 21116 7052 21180
rect 7116 21116 7117 21180
rect 7051 21115 7117 21116
rect 6867 19412 6933 19413
rect 6867 19348 6868 19412
rect 6932 19348 6933 19412
rect 6867 19347 6933 19348
rect 6131 18732 6197 18733
rect 6131 18668 6132 18732
rect 6196 18668 6197 18732
rect 6131 18667 6197 18668
rect 7054 17509 7114 21115
rect 7238 17917 7298 23291
rect 7419 22540 7485 22541
rect 7419 22476 7420 22540
rect 7484 22476 7485 22540
rect 7419 22475 7485 22476
rect 7235 17916 7301 17917
rect 7235 17852 7236 17916
rect 7300 17852 7301 17916
rect 7235 17851 7301 17852
rect 7051 17508 7117 17509
rect 7051 17444 7052 17508
rect 7116 17444 7117 17508
rect 7051 17443 7117 17444
rect 5947 16964 6013 16965
rect 5947 16900 5948 16964
rect 6012 16900 6013 16964
rect 5947 16899 6013 16900
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 7422 16557 7482 22475
rect 7787 21180 7853 21181
rect 7787 21116 7788 21180
rect 7852 21116 7853 21180
rect 7787 21115 7853 21116
rect 7603 20772 7669 20773
rect 7603 20708 7604 20772
rect 7668 20708 7669 20772
rect 7603 20707 7669 20708
rect 7606 19821 7666 20707
rect 7603 19820 7669 19821
rect 7603 19756 7604 19820
rect 7668 19756 7669 19820
rect 7603 19755 7669 19756
rect 7790 19549 7850 21115
rect 7974 20909 8034 25875
rect 9262 25397 9322 28867
rect 9446 26077 9506 35123
rect 9627 30564 9693 30565
rect 9627 30500 9628 30564
rect 9692 30500 9693 30564
rect 9627 30499 9693 30500
rect 9630 28933 9690 30499
rect 9627 28932 9693 28933
rect 9627 28868 9628 28932
rect 9692 28868 9693 28932
rect 9627 28867 9693 28868
rect 9443 26076 9509 26077
rect 9443 26012 9444 26076
rect 9508 26012 9509 26076
rect 9443 26011 9509 26012
rect 9259 25396 9325 25397
rect 9259 25332 9260 25396
rect 9324 25332 9325 25396
rect 9259 25331 9325 25332
rect 8155 24036 8221 24037
rect 8155 23972 8156 24036
rect 8220 23972 8221 24036
rect 8155 23971 8221 23972
rect 7971 20908 8037 20909
rect 7971 20844 7972 20908
rect 8036 20844 8037 20908
rect 7971 20843 8037 20844
rect 8158 20093 8218 23971
rect 9262 22541 9322 25331
rect 9627 23084 9693 23085
rect 9627 23020 9628 23084
rect 9692 23020 9693 23084
rect 9627 23019 9693 23020
rect 9259 22540 9325 22541
rect 9259 22476 9260 22540
rect 9324 22476 9325 22540
rect 9259 22475 9325 22476
rect 8339 22268 8405 22269
rect 8339 22204 8340 22268
rect 8404 22204 8405 22268
rect 8339 22203 8405 22204
rect 8155 20092 8221 20093
rect 8155 20028 8156 20092
rect 8220 20028 8221 20092
rect 8155 20027 8221 20028
rect 7787 19548 7853 19549
rect 7787 19484 7788 19548
rect 7852 19484 7853 19548
rect 7787 19483 7853 19484
rect 8342 17917 8402 22203
rect 8707 20908 8773 20909
rect 8707 20844 8708 20908
rect 8772 20844 8773 20908
rect 8707 20843 8773 20844
rect 8523 20636 8589 20637
rect 8523 20572 8524 20636
rect 8588 20572 8589 20636
rect 8523 20571 8589 20572
rect 8339 17916 8405 17917
rect 8339 17852 8340 17916
rect 8404 17852 8405 17916
rect 8339 17851 8405 17852
rect 7419 16556 7485 16557
rect 7419 16492 7420 16556
rect 7484 16492 7485 16556
rect 7419 16491 7485 16492
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 8526 15197 8586 20571
rect 8710 20229 8770 20843
rect 8707 20228 8773 20229
rect 8707 20164 8708 20228
rect 8772 20164 8773 20228
rect 8707 20163 8773 20164
rect 9630 17781 9690 23019
rect 10366 22949 10426 38387
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 41920 35248 42480
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 25635 36004 25701 36005
rect 25635 35940 25636 36004
rect 25700 35940 25701 36004
rect 25635 35939 25701 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 11467 34644 11533 34645
rect 11467 34580 11468 34644
rect 11532 34580 11533 34644
rect 11467 34579 11533 34580
rect 10915 30428 10981 30429
rect 10915 30364 10916 30428
rect 10980 30364 10981 30428
rect 10915 30363 10981 30364
rect 10363 22948 10429 22949
rect 10363 22884 10364 22948
rect 10428 22884 10429 22948
rect 10363 22883 10429 22884
rect 9995 22132 10061 22133
rect 9995 22068 9996 22132
rect 10060 22068 10061 22132
rect 9995 22067 10061 22068
rect 9998 19549 10058 22067
rect 10918 20773 10978 30363
rect 11470 25397 11530 34579
rect 11835 34508 11901 34509
rect 11835 34444 11836 34508
rect 11900 34444 11901 34508
rect 11835 34443 11901 34444
rect 11838 25669 11898 34443
rect 19568 33760 19888 34784
rect 25451 34236 25517 34237
rect 25451 34172 25452 34236
rect 25516 34172 25517 34236
rect 25451 34171 25517 34172
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 18459 32740 18525 32741
rect 18459 32676 18460 32740
rect 18524 32676 18525 32740
rect 18459 32675 18525 32676
rect 18091 31380 18157 31381
rect 18091 31316 18092 31380
rect 18156 31316 18157 31380
rect 18091 31315 18157 31316
rect 16435 30564 16501 30565
rect 16435 30500 16436 30564
rect 16500 30500 16501 30564
rect 16435 30499 16501 30500
rect 14595 30428 14661 30429
rect 14595 30364 14596 30428
rect 14660 30364 14661 30428
rect 14595 30363 14661 30364
rect 14963 30428 15029 30429
rect 14963 30364 14964 30428
rect 15028 30364 15029 30428
rect 14963 30363 15029 30364
rect 14598 27301 14658 30363
rect 13859 27300 13925 27301
rect 13859 27236 13860 27300
rect 13924 27236 13925 27300
rect 13859 27235 13925 27236
rect 14595 27300 14661 27301
rect 14595 27236 14596 27300
rect 14660 27236 14661 27300
rect 14595 27235 14661 27236
rect 13675 26756 13741 26757
rect 13675 26692 13676 26756
rect 13740 26692 13741 26756
rect 13675 26691 13741 26692
rect 11835 25668 11901 25669
rect 11835 25604 11836 25668
rect 11900 25604 11901 25668
rect 11835 25603 11901 25604
rect 11467 25396 11533 25397
rect 11467 25332 11468 25396
rect 11532 25332 11533 25396
rect 11467 25331 11533 25332
rect 12019 23628 12085 23629
rect 12019 23564 12020 23628
rect 12084 23564 12085 23628
rect 12019 23563 12085 23564
rect 11835 22812 11901 22813
rect 11835 22748 11836 22812
rect 11900 22748 11901 22812
rect 11835 22747 11901 22748
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 9995 19548 10061 19549
rect 9995 19484 9996 19548
rect 10060 19484 10061 19548
rect 9995 19483 10061 19484
rect 11102 18461 11162 20707
rect 11838 19413 11898 22747
rect 11835 19412 11901 19413
rect 11835 19348 11836 19412
rect 11900 19348 11901 19412
rect 11835 19347 11901 19348
rect 11099 18460 11165 18461
rect 11099 18396 11100 18460
rect 11164 18396 11165 18460
rect 11099 18395 11165 18396
rect 9627 17780 9693 17781
rect 9627 17716 9628 17780
rect 9692 17716 9693 17780
rect 9627 17715 9693 17716
rect 8523 15196 8589 15197
rect 8523 15132 8524 15196
rect 8588 15132 8589 15196
rect 8523 15131 8589 15132
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 12022 8941 12082 23563
rect 12571 22540 12637 22541
rect 12571 22476 12572 22540
rect 12636 22476 12637 22540
rect 12571 22475 12637 22476
rect 12574 16557 12634 22475
rect 12755 20772 12821 20773
rect 12755 20708 12756 20772
rect 12820 20708 12821 20772
rect 12755 20707 12821 20708
rect 12758 17917 12818 20707
rect 13307 19820 13373 19821
rect 13307 19756 13308 19820
rect 13372 19756 13373 19820
rect 13307 19755 13373 19756
rect 12755 17916 12821 17917
rect 12755 17852 12756 17916
rect 12820 17852 12821 17916
rect 12755 17851 12821 17852
rect 12571 16556 12637 16557
rect 12571 16492 12572 16556
rect 12636 16492 12637 16556
rect 12571 16491 12637 16492
rect 13310 16149 13370 19755
rect 13678 18053 13738 26691
rect 13675 18052 13741 18053
rect 13675 17988 13676 18052
rect 13740 17988 13741 18052
rect 13675 17987 13741 17988
rect 13862 16557 13922 27235
rect 14411 24988 14477 24989
rect 14411 24924 14412 24988
rect 14476 24924 14477 24988
rect 14411 24923 14477 24924
rect 14414 16557 14474 24923
rect 14598 21997 14658 27235
rect 14595 21996 14661 21997
rect 14595 21932 14596 21996
rect 14660 21932 14661 21996
rect 14595 21931 14661 21932
rect 14966 21589 15026 30363
rect 16251 28796 16317 28797
rect 16251 28732 16252 28796
rect 16316 28732 16317 28796
rect 16251 28731 16317 28732
rect 16254 25261 16314 28731
rect 16438 26621 16498 30499
rect 17907 29204 17973 29205
rect 17907 29140 17908 29204
rect 17972 29140 17973 29204
rect 17907 29139 17973 29140
rect 16619 27980 16685 27981
rect 16619 27916 16620 27980
rect 16684 27916 16685 27980
rect 16619 27915 16685 27916
rect 16435 26620 16501 26621
rect 16435 26556 16436 26620
rect 16500 26556 16501 26620
rect 16435 26555 16501 26556
rect 16435 26076 16501 26077
rect 16435 26012 16436 26076
rect 16500 26012 16501 26076
rect 16435 26011 16501 26012
rect 16251 25260 16317 25261
rect 16251 25196 16252 25260
rect 16316 25196 16317 25260
rect 16251 25195 16317 25196
rect 15515 25124 15581 25125
rect 15515 25060 15516 25124
rect 15580 25060 15581 25124
rect 15515 25059 15581 25060
rect 15147 22404 15213 22405
rect 15147 22340 15148 22404
rect 15212 22340 15213 22404
rect 15147 22339 15213 22340
rect 14963 21588 15029 21589
rect 14963 21524 14964 21588
rect 15028 21524 15029 21588
rect 14963 21523 15029 21524
rect 15150 19413 15210 22339
rect 15518 19821 15578 25059
rect 16438 23085 16498 26011
rect 16622 25397 16682 27915
rect 17910 27573 17970 29139
rect 17907 27572 17973 27573
rect 17907 27508 17908 27572
rect 17972 27508 17973 27572
rect 17907 27507 17973 27508
rect 17355 26348 17421 26349
rect 17355 26284 17356 26348
rect 17420 26284 17421 26348
rect 17355 26283 17421 26284
rect 16619 25396 16685 25397
rect 16619 25332 16620 25396
rect 16684 25332 16685 25396
rect 16619 25331 16685 25332
rect 17171 24988 17237 24989
rect 17171 24924 17172 24988
rect 17236 24924 17237 24988
rect 17171 24923 17237 24924
rect 16435 23084 16501 23085
rect 16435 23020 16436 23084
rect 16500 23020 16501 23084
rect 16435 23019 16501 23020
rect 16987 23084 17053 23085
rect 16987 23020 16988 23084
rect 17052 23020 17053 23084
rect 16987 23019 17053 23020
rect 16438 21453 16498 23019
rect 16435 21452 16501 21453
rect 16435 21388 16436 21452
rect 16500 21388 16501 21452
rect 16435 21387 16501 21388
rect 15515 19820 15581 19821
rect 15515 19756 15516 19820
rect 15580 19756 15581 19820
rect 15515 19755 15581 19756
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 15150 18189 15210 19347
rect 16990 19277 17050 23019
rect 17174 21453 17234 24923
rect 17171 21452 17237 21453
rect 17171 21388 17172 21452
rect 17236 21388 17237 21452
rect 17171 21387 17237 21388
rect 17358 19277 17418 26283
rect 17539 25260 17605 25261
rect 17539 25196 17540 25260
rect 17604 25196 17605 25260
rect 17539 25195 17605 25196
rect 17542 19277 17602 25195
rect 17723 23492 17789 23493
rect 17723 23428 17724 23492
rect 17788 23428 17789 23492
rect 17723 23427 17789 23428
rect 17726 20365 17786 23427
rect 18094 22949 18154 31315
rect 18091 22948 18157 22949
rect 18091 22884 18092 22948
rect 18156 22884 18157 22948
rect 18091 22883 18157 22884
rect 18275 22812 18341 22813
rect 18275 22748 18276 22812
rect 18340 22748 18341 22812
rect 18275 22747 18341 22748
rect 18278 21045 18338 22747
rect 18275 21044 18341 21045
rect 18275 20980 18276 21044
rect 18340 20980 18341 21044
rect 18275 20979 18341 20980
rect 17907 20908 17973 20909
rect 17907 20844 17908 20908
rect 17972 20844 17973 20908
rect 17907 20843 17973 20844
rect 17723 20364 17789 20365
rect 17723 20300 17724 20364
rect 17788 20300 17789 20364
rect 17723 20299 17789 20300
rect 17910 19821 17970 20843
rect 18462 20637 18522 32675
rect 19568 32672 19888 33696
rect 24899 33420 24965 33421
rect 24899 33356 24900 33420
rect 24964 33356 24965 33420
rect 24899 33355 24965 33356
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 21035 30836 21101 30837
rect 21035 30772 21036 30836
rect 21100 30772 21101 30836
rect 21035 30771 21101 30772
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 20667 26756 20733 26757
rect 20667 26692 20668 26756
rect 20732 26692 20733 26756
rect 20667 26691 20733 26692
rect 20299 26212 20365 26213
rect 20299 26148 20300 26212
rect 20364 26148 20365 26212
rect 20299 26147 20365 26148
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 20302 25397 20362 26147
rect 20299 25396 20365 25397
rect 20299 25332 20300 25396
rect 20364 25332 20365 25396
rect 20299 25331 20365 25332
rect 20115 25124 20181 25125
rect 20115 25060 20116 25124
rect 20180 25060 20181 25124
rect 20115 25059 20181 25060
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19011 24716 19077 24717
rect 19011 24652 19012 24716
rect 19076 24652 19077 24716
rect 19011 24651 19077 24652
rect 18643 22404 18709 22405
rect 18643 22340 18644 22404
rect 18708 22340 18709 22404
rect 18643 22339 18709 22340
rect 18459 20636 18525 20637
rect 18459 20572 18460 20636
rect 18524 20572 18525 20636
rect 18459 20571 18525 20572
rect 17907 19820 17973 19821
rect 17907 19756 17908 19820
rect 17972 19756 17973 19820
rect 17907 19755 17973 19756
rect 16987 19276 17053 19277
rect 16987 19212 16988 19276
rect 17052 19212 17053 19276
rect 16987 19211 17053 19212
rect 17355 19276 17421 19277
rect 17355 19212 17356 19276
rect 17420 19212 17421 19276
rect 17355 19211 17421 19212
rect 17539 19276 17605 19277
rect 17539 19212 17540 19276
rect 17604 19212 17605 19276
rect 17539 19211 17605 19212
rect 15147 18188 15213 18189
rect 15147 18124 15148 18188
rect 15212 18124 15213 18188
rect 15147 18123 15213 18124
rect 18646 16557 18706 22339
rect 19014 21725 19074 24651
rect 19195 24036 19261 24037
rect 19195 23972 19196 24036
rect 19260 23972 19261 24036
rect 19195 23971 19261 23972
rect 19198 21861 19258 23971
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19379 23900 19445 23901
rect 19379 23836 19380 23900
rect 19444 23836 19445 23900
rect 19379 23835 19445 23836
rect 19382 22677 19442 23835
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19379 22676 19445 22677
rect 19379 22612 19380 22676
rect 19444 22612 19445 22676
rect 19379 22611 19445 22612
rect 19195 21860 19261 21861
rect 19195 21796 19196 21860
rect 19260 21796 19261 21860
rect 19195 21795 19261 21796
rect 19568 21792 19888 22816
rect 20118 22405 20178 25059
rect 20299 24988 20365 24989
rect 20299 24924 20300 24988
rect 20364 24924 20365 24988
rect 20299 24923 20365 24924
rect 20483 24988 20549 24989
rect 20483 24924 20484 24988
rect 20548 24924 20549 24988
rect 20483 24923 20549 24924
rect 20115 22404 20181 22405
rect 20115 22340 20116 22404
rect 20180 22340 20181 22404
rect 20115 22339 20181 22340
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19011 21724 19077 21725
rect 19011 21660 19012 21724
rect 19076 21660 19077 21724
rect 19011 21659 19077 21660
rect 19568 20704 19888 21728
rect 20118 21045 20178 22339
rect 20302 22133 20362 24923
rect 20299 22132 20365 22133
rect 20299 22068 20300 22132
rect 20364 22068 20365 22132
rect 20299 22067 20365 22068
rect 20299 21588 20365 21589
rect 20299 21524 20300 21588
rect 20364 21524 20365 21588
rect 20299 21523 20365 21524
rect 20115 21044 20181 21045
rect 20115 20980 20116 21044
rect 20180 20980 20181 21044
rect 20115 20979 20181 20980
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 20302 20229 20362 21523
rect 20299 20228 20365 20229
rect 20299 20164 20300 20228
rect 20364 20164 20365 20228
rect 20299 20163 20365 20164
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20486 19413 20546 24923
rect 20670 23357 20730 26691
rect 20851 24172 20917 24173
rect 20851 24108 20852 24172
rect 20916 24108 20917 24172
rect 20851 24107 20917 24108
rect 20667 23356 20733 23357
rect 20667 23292 20668 23356
rect 20732 23292 20733 23356
rect 20667 23291 20733 23292
rect 20854 21045 20914 24107
rect 20851 21044 20917 21045
rect 20851 20980 20852 21044
rect 20916 20980 20917 21044
rect 20851 20979 20917 20980
rect 20667 20772 20733 20773
rect 20667 20708 20668 20772
rect 20732 20708 20733 20772
rect 20667 20707 20733 20708
rect 20483 19412 20549 19413
rect 20483 19348 20484 19412
rect 20548 19348 20549 19412
rect 20483 19347 20549 19348
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 13859 16556 13925 16557
rect 13859 16492 13860 16556
rect 13924 16492 13925 16556
rect 13859 16491 13925 16492
rect 14411 16556 14477 16557
rect 14411 16492 14412 16556
rect 14476 16492 14477 16556
rect 14411 16491 14477 16492
rect 18643 16556 18709 16557
rect 18643 16492 18644 16556
rect 18708 16492 18709 16556
rect 18643 16491 18709 16492
rect 19568 16352 19888 17376
rect 20670 16557 20730 20707
rect 21038 18597 21098 30771
rect 23243 29068 23309 29069
rect 23243 29004 23244 29068
rect 23308 29004 23309 29068
rect 23243 29003 23309 29004
rect 23059 25260 23125 25261
rect 23059 25196 23060 25260
rect 23124 25196 23125 25260
rect 23059 25195 23125 25196
rect 21403 24988 21469 24989
rect 21403 24924 21404 24988
rect 21468 24924 21469 24988
rect 21403 24923 21469 24924
rect 21219 23900 21285 23901
rect 21219 23836 21220 23900
rect 21284 23836 21285 23900
rect 21219 23835 21285 23836
rect 21222 21589 21282 23835
rect 21406 21997 21466 24923
rect 22691 24036 22757 24037
rect 22691 23972 22692 24036
rect 22756 23972 22757 24036
rect 22691 23971 22757 23972
rect 21587 22404 21653 22405
rect 21587 22340 21588 22404
rect 21652 22340 21653 22404
rect 21587 22339 21653 22340
rect 21403 21996 21469 21997
rect 21403 21932 21404 21996
rect 21468 21932 21469 21996
rect 21403 21931 21469 21932
rect 21219 21588 21285 21589
rect 21219 21524 21220 21588
rect 21284 21524 21285 21588
rect 21219 21523 21285 21524
rect 21590 19413 21650 22339
rect 22694 21453 22754 23971
rect 22691 21452 22757 21453
rect 22691 21388 22692 21452
rect 22756 21388 22757 21452
rect 22691 21387 22757 21388
rect 22875 21180 22941 21181
rect 22875 21116 22876 21180
rect 22940 21116 22941 21180
rect 22875 21115 22941 21116
rect 22878 19957 22938 21115
rect 23062 20909 23122 25195
rect 23059 20908 23125 20909
rect 23059 20844 23060 20908
rect 23124 20844 23125 20908
rect 23059 20843 23125 20844
rect 22875 19956 22941 19957
rect 22875 19892 22876 19956
rect 22940 19892 22941 19956
rect 22875 19891 22941 19892
rect 21587 19412 21653 19413
rect 21587 19348 21588 19412
rect 21652 19348 21653 19412
rect 21587 19347 21653 19348
rect 23246 19277 23306 29003
rect 24902 28797 24962 33355
rect 25267 31516 25333 31517
rect 25267 31452 25268 31516
rect 25332 31452 25333 31516
rect 25267 31451 25333 31452
rect 25270 30157 25330 31451
rect 25454 31109 25514 34171
rect 25451 31108 25517 31109
rect 25451 31044 25452 31108
rect 25516 31044 25517 31108
rect 25451 31043 25517 31044
rect 25267 30156 25333 30157
rect 25267 30092 25268 30156
rect 25332 30092 25333 30156
rect 25267 30091 25333 30092
rect 24899 28796 24965 28797
rect 24899 28732 24900 28796
rect 24964 28732 24965 28796
rect 24899 28731 24965 28732
rect 25638 27573 25698 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 26371 33556 26437 33557
rect 26371 33492 26372 33556
rect 26436 33492 26437 33556
rect 26371 33491 26437 33492
rect 25819 32060 25885 32061
rect 25819 31996 25820 32060
rect 25884 31996 25885 32060
rect 25819 31995 25885 31996
rect 25822 31109 25882 31995
rect 25819 31108 25885 31109
rect 25819 31044 25820 31108
rect 25884 31044 25885 31108
rect 25819 31043 25885 31044
rect 26187 30972 26253 30973
rect 26187 30908 26188 30972
rect 26252 30908 26253 30972
rect 26187 30907 26253 30908
rect 25635 27572 25701 27573
rect 25635 27508 25636 27572
rect 25700 27508 25701 27572
rect 25635 27507 25701 27508
rect 26190 27301 26250 30907
rect 26374 30429 26434 33491
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 27659 33148 27725 33149
rect 27659 33084 27660 33148
rect 27724 33084 27725 33148
rect 27659 33083 27725 33084
rect 26555 30564 26621 30565
rect 26555 30500 26556 30564
rect 26620 30500 26621 30564
rect 26555 30499 26621 30500
rect 26371 30428 26437 30429
rect 26371 30364 26372 30428
rect 26436 30364 26437 30428
rect 26371 30363 26437 30364
rect 26558 28933 26618 30499
rect 26555 28932 26621 28933
rect 26555 28868 26556 28932
rect 26620 28868 26621 28932
rect 26555 28867 26621 28868
rect 27662 28389 27722 33083
rect 28579 32740 28645 32741
rect 28579 32676 28580 32740
rect 28644 32676 28645 32740
rect 28579 32675 28645 32676
rect 27659 28388 27725 28389
rect 27659 28324 27660 28388
rect 27724 28324 27725 28388
rect 27659 28323 27725 28324
rect 26187 27300 26253 27301
rect 26187 27236 26188 27300
rect 26252 27236 26253 27300
rect 26187 27235 26253 27236
rect 26923 27164 26989 27165
rect 26923 27100 26924 27164
rect 26988 27100 26989 27164
rect 26923 27099 26989 27100
rect 25267 26212 25333 26213
rect 25267 26148 25268 26212
rect 25332 26148 25333 26212
rect 25267 26147 25333 26148
rect 24163 26076 24229 26077
rect 24163 26012 24164 26076
rect 24228 26012 24229 26076
rect 24163 26011 24229 26012
rect 23427 22132 23493 22133
rect 23427 22068 23428 22132
rect 23492 22068 23493 22132
rect 23427 22067 23493 22068
rect 23430 20637 23490 22067
rect 24166 20773 24226 26011
rect 24347 23764 24413 23765
rect 24347 23700 24348 23764
rect 24412 23700 24413 23764
rect 24347 23699 24413 23700
rect 24163 20772 24229 20773
rect 24163 20708 24164 20772
rect 24228 20708 24229 20772
rect 24163 20707 24229 20708
rect 23427 20636 23493 20637
rect 23427 20572 23428 20636
rect 23492 20572 23493 20636
rect 23427 20571 23493 20572
rect 23243 19276 23309 19277
rect 23243 19212 23244 19276
rect 23308 19212 23309 19276
rect 23243 19211 23309 19212
rect 21035 18596 21101 18597
rect 21035 18532 21036 18596
rect 21100 18532 21101 18596
rect 21035 18531 21101 18532
rect 24166 17917 24226 20707
rect 24350 20501 24410 23699
rect 25270 22110 25330 26147
rect 26371 25804 26437 25805
rect 26371 25740 26372 25804
rect 26436 25740 26437 25804
rect 26371 25739 26437 25740
rect 24902 22050 25330 22110
rect 24347 20500 24413 20501
rect 24347 20436 24348 20500
rect 24412 20436 24413 20500
rect 24347 20435 24413 20436
rect 24163 17916 24229 17917
rect 24163 17852 24164 17916
rect 24228 17852 24229 17916
rect 24163 17851 24229 17852
rect 20667 16556 20733 16557
rect 20667 16492 20668 16556
rect 20732 16492 20733 16556
rect 20667 16491 20733 16492
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 13307 16148 13373 16149
rect 13307 16084 13308 16148
rect 13372 16084 13373 16148
rect 13307 16083 13373 16084
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 12019 8940 12085 8941
rect 12019 8876 12020 8940
rect 12084 8876 12085 8940
rect 12019 8875 12085 8876
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 3187 4044 3253 4045
rect 3187 3980 3188 4044
rect 3252 3980 3253 4044
rect 3187 3979 3253 3980
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 24902 2685 24962 22050
rect 26374 20637 26434 25739
rect 26555 25668 26621 25669
rect 26555 25604 26556 25668
rect 26620 25604 26621 25668
rect 26555 25603 26621 25604
rect 26558 23901 26618 25603
rect 26926 25533 26986 27099
rect 27659 26348 27725 26349
rect 27659 26284 27660 26348
rect 27724 26284 27725 26348
rect 27659 26283 27725 26284
rect 26923 25532 26989 25533
rect 26923 25468 26924 25532
rect 26988 25468 26989 25532
rect 26923 25467 26989 25468
rect 26555 23900 26621 23901
rect 26555 23836 26556 23900
rect 26620 23836 26621 23900
rect 26555 23835 26621 23836
rect 27107 23492 27173 23493
rect 27107 23428 27108 23492
rect 27172 23428 27173 23492
rect 27107 23427 27173 23428
rect 26371 20636 26437 20637
rect 26371 20572 26372 20636
rect 26436 20572 26437 20636
rect 26371 20571 26437 20572
rect 27110 18733 27170 23427
rect 27662 20909 27722 26283
rect 28582 23085 28642 32675
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 28579 23084 28645 23085
rect 28579 23020 28580 23084
rect 28644 23020 28645 23084
rect 28579 23019 28645 23020
rect 27843 22540 27909 22541
rect 27843 22476 27844 22540
rect 27908 22476 27909 22540
rect 27843 22475 27909 22476
rect 27659 20908 27725 20909
rect 27659 20844 27660 20908
rect 27724 20844 27725 20908
rect 27659 20843 27725 20844
rect 27846 20229 27906 22475
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 27843 20228 27909 20229
rect 27843 20164 27844 20228
rect 27908 20164 27909 20228
rect 27843 20163 27909 20164
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 27107 18732 27173 18733
rect 27107 18668 27108 18732
rect 27172 18668 27173 18732
rect 27107 18667 27173 18668
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24899 2684 24965 2685
rect 24899 2620 24900 2684
rect 24964 2620 24965 2684
rect 24899 2619 24965 2620
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _1025_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1688980957
transform 1 0 20424 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1688980957
transform 1 0 19412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1688980957
transform 1 0 29716 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1688980957
transform 1 0 14904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1688980957
transform 1 0 22724 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1688980957
transform 1 0 25024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1688980957
transform 1 0 21804 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1688980957
transform 1 0 20792 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1040_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1041_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _1042_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1043_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1044_
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _1045_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _1046_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1047_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1048_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _1049_
timestamp 1688980957
transform 1 0 18308 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1050_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21528 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1051_
timestamp 1688980957
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1052_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1053_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1054_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _1055_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1056_
timestamp 1688980957
transform 1 0 19320 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _1057_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1058_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1059_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _1060_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1688980957
transform 1 0 20332 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1063_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_2  _1064_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1065_
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1066_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1067_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1068_
timestamp 1688980957
transform 1 0 19320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp 1688980957
transform 1 0 21344 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1070_
timestamp 1688980957
transform 1 0 19412 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1071_
timestamp 1688980957
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _1072_
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1073_
timestamp 1688980957
transform 1 0 17204 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1074_
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _1075_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _1076_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1077_
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1078_
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1079_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1080_
timestamp 1688980957
transform 1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_4  _1081_
timestamp 1688980957
transform 1 0 17848 0 -1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_2  _1082_
timestamp 1688980957
transform 1 0 19412 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_4  _1083_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1084_
timestamp 1688980957
transform 1 0 17756 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _1085_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__and4_2  _1086_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _1087_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_4  _1088_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 33728
box -38 -48 1326 592
use sky130_fd_sc_hd__nand4b_4  _1089_
timestamp 1688980957
transform 1 0 17664 0 -1 33728
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_1  _1090_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_4  _1091_
timestamp 1688980957
transform 1 0 18584 0 -1 34816
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _1092_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_8  _1093_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _1094_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1095_
timestamp 1688980957
transform 1 0 8280 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _1097_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_4  _1098_
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1099_
timestamp 1688980957
transform 1 0 15272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1688980957
transform 1 0 20424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_4  _1101_
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1103_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1104_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1105_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1106_
timestamp 1688980957
transform 1 0 16836 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _1107_
timestamp 1688980957
transform 1 0 19872 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1108_
timestamp 1688980957
transform 1 0 20424 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1109_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1110_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1111_
timestamp 1688980957
transform 1 0 19504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1112_
timestamp 1688980957
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1113_
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _1114_
timestamp 1688980957
transform 1 0 21712 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1115_
timestamp 1688980957
transform 1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1117_
timestamp 1688980957
transform 1 0 20792 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1118_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1688980957
transform 1 0 20148 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1120_
timestamp 1688980957
transform 1 0 19688 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1121_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _1123_
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1124_
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1125_
timestamp 1688980957
transform 1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1126_
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1127_
timestamp 1688980957
transform 1 0 17664 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1688980957
transform 1 0 19228 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1129_
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _1130_
timestamp 1688980957
transform 1 0 15088 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1131_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1133_
timestamp 1688980957
transform 1 0 20056 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1134_
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1135_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1136_
timestamp 1688980957
transform 1 0 21344 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1137_
timestamp 1688980957
transform 1 0 21252 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1688980957
transform 1 0 20884 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1139_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_8  _1140_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _1141_
timestamp 1688980957
transform 1 0 17664 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _1142_
timestamp 1688980957
transform 1 0 14076 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1144_
timestamp 1688980957
transform 1 0 17572 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1145_
timestamp 1688980957
transform 1 0 18032 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _1146_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1147_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1148_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _1149_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_2  _1150_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1151_
timestamp 1688980957
transform 1 0 13524 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1152_
timestamp 1688980957
transform 1 0 12420 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1153_
timestamp 1688980957
transform 1 0 14720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1154_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1156_
timestamp 1688980957
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1157_
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1158_
timestamp 1688980957
transform 1 0 6900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1159_
timestamp 1688980957
transform 1 0 5520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1160_
timestamp 1688980957
transform 1 0 6440 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1161_
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1162_
timestamp 1688980957
transform 1 0 6164 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1163_
timestamp 1688980957
transform 1 0 28888 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1164_
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1165_
timestamp 1688980957
transform 1 0 6900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1166_
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1167_
timestamp 1688980957
transform 1 0 7176 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 1688980957
transform 1 0 5428 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1169_
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1170_
timestamp 1688980957
transform 1 0 30728 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1171_
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1172_
timestamp 1688980957
transform 1 0 7636 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1173_
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1174_
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1175_
timestamp 1688980957
transform 1 0 15180 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1176_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1177_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1178_
timestamp 1688980957
transform 1 0 26956 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1180_
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1182_
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1183_
timestamp 1688980957
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1184_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211ai_1  _1185_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1186_
timestamp 1688980957
transform 1 0 11868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1187_
timestamp 1688980957
transform 1 0 29624 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1188_
timestamp 1688980957
transform 1 0 11316 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1189_
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1190_
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1191_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1192_
timestamp 1688980957
transform 1 0 11316 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1194_
timestamp 1688980957
transform 1 0 23276 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1195_
timestamp 1688980957
transform 1 0 12604 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1196_
timestamp 1688980957
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1197_
timestamp 1688980957
transform 1 0 11684 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1688980957
transform 1 0 19504 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1199_
timestamp 1688980957
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1200_
timestamp 1688980957
transform 1 0 17572 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211ai_2  _1201_
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1203_
timestamp 1688980957
transform 1 0 25852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1204_
timestamp 1688980957
transform 1 0 12696 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1205_
timestamp 1688980957
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1206_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1207_
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1209_
timestamp 1688980957
transform 1 0 4968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1210_
timestamp 1688980957
transform 1 0 4784 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1211_
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1212_
timestamp 1688980957
transform 1 0 4784 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1213_
timestamp 1688980957
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1214_
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1215_
timestamp 1688980957
transform 1 0 6716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1216_
timestamp 1688980957
transform 1 0 8096 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _1217_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1218_
timestamp 1688980957
transform 1 0 9752 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _1219_
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1220_
timestamp 1688980957
transform 1 0 9016 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _1221_
timestamp 1688980957
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1222_
timestamp 1688980957
transform 1 0 13340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1223_
timestamp 1688980957
transform 1 0 14904 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1224_
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1225_
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _1227_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1228_
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1229_
timestamp 1688980957
transform 1 0 21804 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1230_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _1231_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_2  _1232_
timestamp 1688980957
transform 1 0 42596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1233_
timestamp 1688980957
transform 1 0 42964 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1234_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42044 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1688980957
transform 1 0 15456 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _1236_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1237_
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1238_
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1688980957
transform 1 0 24196 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1240_
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1241_
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1242_
timestamp 1688980957
transform 1 0 23552 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1243_
timestamp 1688980957
transform 1 0 23000 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1244_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1245_
timestamp 1688980957
transform 1 0 22080 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1246_
timestamp 1688980957
transform 1 0 23000 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1247_
timestamp 1688980957
transform 1 0 15548 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1248_
timestamp 1688980957
transform 1 0 26036 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1249_
timestamp 1688980957
transform 1 0 25852 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1250_
timestamp 1688980957
transform 1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1251_
timestamp 1688980957
transform 1 0 28428 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1252_
timestamp 1688980957
transform 1 0 28428 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1253_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27784 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1254_
timestamp 1688980957
transform 1 0 26496 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1688980957
transform 1 0 25392 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1256_
timestamp 1688980957
transform 1 0 25208 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1688980957
transform 1 0 25392 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1258_
timestamp 1688980957
transform 1 0 25852 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1259_
timestamp 1688980957
transform 1 0 23276 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1260_
timestamp 1688980957
transform 1 0 24932 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1261_
timestamp 1688980957
transform 1 0 25852 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1262_
timestamp 1688980957
transform 1 0 26864 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1263_
timestamp 1688980957
transform 1 0 28704 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1264_
timestamp 1688980957
transform 1 0 27968 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1265_
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1266_
timestamp 1688980957
transform 1 0 28060 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1688980957
transform 1 0 27968 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1268_
timestamp 1688980957
transform 1 0 21896 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _1269_
timestamp 1688980957
transform 1 0 22172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1270_
timestamp 1688980957
transform 1 0 23460 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1271_
timestamp 1688980957
transform 1 0 28244 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1272_
timestamp 1688980957
transform 1 0 29532 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1273_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1274_
timestamp 1688980957
transform 1 0 25300 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1688980957
transform 1 0 27232 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1688980957
transform 1 0 28796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1688980957
transform 1 0 27324 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1278_
timestamp 1688980957
transform 1 0 27692 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1279_
timestamp 1688980957
transform 1 0 28612 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1280_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 1688980957
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1282_
timestamp 1688980957
transform 1 0 25852 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1283_
timestamp 1688980957
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1284_
timestamp 1688980957
transform 1 0 28428 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1688980957
transform 1 0 25944 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1286_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1287_
timestamp 1688980957
transform 1 0 26128 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1289_
timestamp 1688980957
transform 1 0 25208 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1290_
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1291_
timestamp 1688980957
transform 1 0 27140 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1292_
timestamp 1688980957
transform 1 0 26772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1293_
timestamp 1688980957
transform 1 0 27784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1688980957
transform 1 0 27324 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1688980957
transform 1 0 25024 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1296_
timestamp 1688980957
transform 1 0 25576 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1688980957
transform 1 0 26036 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1298_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26404 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1299_
timestamp 1688980957
transform 1 0 26404 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1300_
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1301_
timestamp 1688980957
transform 1 0 24840 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1302_
timestamp 1688980957
transform 1 0 27968 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1688980957
transform 1 0 27416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1304_
timestamp 1688980957
transform 1 0 27784 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1305_
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1688980957
transform 1 0 25392 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1307_
timestamp 1688980957
transform 1 0 27600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1308_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1688980957
transform 1 0 27784 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1310_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27692 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1311_
timestamp 1688980957
transform 1 0 28612 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1312_
timestamp 1688980957
transform 1 0 28336 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1313_
timestamp 1688980957
transform 1 0 28336 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1314_
timestamp 1688980957
transform 1 0 27600 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1315_
timestamp 1688980957
transform 1 0 23644 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1316_
timestamp 1688980957
transform 1 0 28704 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1317_
timestamp 1688980957
transform 1 0 25668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1318_
timestamp 1688980957
transform 1 0 26312 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1319_
timestamp 1688980957
transform 1 0 25760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1688980957
transform 1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1321_
timestamp 1688980957
transform 1 0 24840 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1322_
timestamp 1688980957
transform 1 0 23184 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1323_
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1324_
timestamp 1688980957
transform 1 0 24380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1325_
timestamp 1688980957
transform 1 0 22816 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1326_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1327_
timestamp 1688980957
transform 1 0 24564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1328_
timestamp 1688980957
transform 1 0 24380 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1329_
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1330_
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1331_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _1332_
timestamp 1688980957
transform 1 0 21068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1333_
timestamp 1688980957
transform 1 0 25300 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1334_
timestamp 1688980957
transform 1 0 25760 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 1688980957
transform 1 0 19780 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1336_
timestamp 1688980957
transform 1 0 27692 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1337_
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_8  _1338_
timestamp 1688980957
transform 1 0 19320 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1339_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1340_
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1341_
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1342_
timestamp 1688980957
transform 1 0 22448 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1343_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1346_
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1347_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1348_
timestamp 1688980957
transform 1 0 25852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1688980957
transform 1 0 26864 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1351_
timestamp 1688980957
transform 1 0 27600 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1352_
timestamp 1688980957
transform 1 0 27416 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1688980957
transform 1 0 28888 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1354_
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1688980957
transform 1 0 28060 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1356_
timestamp 1688980957
transform 1 0 28336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1358_
timestamp 1688980957
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1359_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1360_
timestamp 1688980957
transform 1 0 26220 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1361_
timestamp 1688980957
transform 1 0 26496 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _1362_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1363_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21528 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1688980957
transform 1 0 21896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1365_
timestamp 1688980957
transform 1 0 23828 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1366_
timestamp 1688980957
transform 1 0 22172 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1367_
timestamp 1688980957
transform 1 0 22356 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1368_
timestamp 1688980957
transform 1 0 28244 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1369_
timestamp 1688980957
transform 1 0 28244 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1370_
timestamp 1688980957
transform 1 0 23092 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1371_
timestamp 1688980957
transform 1 0 21988 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1372_
timestamp 1688980957
transform 1 0 25668 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _1373_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24932 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1374_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1375_
timestamp 1688980957
transform 1 0 27968 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1376_
timestamp 1688980957
transform 1 0 25852 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1377_
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1378_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1379_
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1380_
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1381_
timestamp 1688980957
transform 1 0 21804 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1382_
timestamp 1688980957
transform 1 0 24288 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1383_
timestamp 1688980957
transform 1 0 24104 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1385_
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1387_
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1388_
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1688980957
transform 1 0 25944 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1688980957
transform 1 0 27416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1391_
timestamp 1688980957
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1393_
timestamp 1688980957
transform 1 0 26680 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1394_
timestamp 1688980957
transform 1 0 26220 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1395_
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1688980957
transform 1 0 28244 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1397_
timestamp 1688980957
transform 1 0 25668 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1398_
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1688980957
transform 1 0 23184 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1688980957
transform 1 0 25852 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1401_
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1402_
timestamp 1688980957
transform 1 0 27692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1403_
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1688980957
transform 1 0 26404 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1405_
timestamp 1688980957
transform 1 0 25116 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1406_
timestamp 1688980957
transform 1 0 26312 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1407_
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1408_
timestamp 1688980957
transform 1 0 27784 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1409_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28336 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1410_
timestamp 1688980957
transform 1 0 25484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1411_
timestamp 1688980957
transform 1 0 26128 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1412_
timestamp 1688980957
transform 1 0 27232 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1413_
timestamp 1688980957
transform 1 0 27692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1414_
timestamp 1688980957
transform 1 0 23276 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1415_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1416_
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1417_
timestamp 1688980957
transform 1 0 24840 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1419_
timestamp 1688980957
transform 1 0 27140 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1420_
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1421_
timestamp 1688980957
transform 1 0 14444 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_4  _1422_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__a21o_2  _1423_
timestamp 1688980957
transform 1 0 14352 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1424_
timestamp 1688980957
transform 1 0 13064 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1425_
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1426_
timestamp 1688980957
transform 1 0 12696 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 1688980957
transform 1 0 11592 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1428_
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1429_
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 1688980957
transform 1 0 10120 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1432_
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1433_
timestamp 1688980957
transform 1 0 8740 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1434_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1435_
timestamp 1688980957
transform 1 0 9108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1436_
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1437_
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1438_
timestamp 1688980957
transform 1 0 6992 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1439_
timestamp 1688980957
transform 1 0 6992 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1440_
timestamp 1688980957
transform 1 0 6440 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1441_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1442_
timestamp 1688980957
transform 1 0 5704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1443_
timestamp 1688980957
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1445_
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1446_
timestamp 1688980957
transform 1 0 7176 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1447_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1448_
timestamp 1688980957
transform 1 0 14352 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1449_
timestamp 1688980957
transform 1 0 14720 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1450_
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_4  _1451_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__a221o_2  _1452_
timestamp 1688980957
transform 1 0 15364 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1453_
timestamp 1688980957
transform 1 0 14168 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1454_
timestamp 1688980957
transform 1 0 13432 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _1455_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1456_
timestamp 1688980957
transform 1 0 16192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1457_
timestamp 1688980957
transform 1 0 16836 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1458_
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1459_
timestamp 1688980957
transform 1 0 17112 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _1460_
timestamp 1688980957
transform 1 0 15824 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1461_
timestamp 1688980957
transform 1 0 4416 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _1462_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1463_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13892 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _1464_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1465_
timestamp 1688980957
transform 1 0 28244 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1466_
timestamp 1688980957
transform 1 0 21896 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1467_
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1468_
timestamp 1688980957
transform 1 0 12144 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1469_
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1470_
timestamp 1688980957
transform 1 0 3772 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _1471_
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1472_
timestamp 1688980957
transform 1 0 14536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1473_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1474_
timestamp 1688980957
transform 1 0 13432 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1475_
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1476_
timestamp 1688980957
transform 1 0 4784 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1477_
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1478_
timestamp 1688980957
transform 1 0 5520 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1479_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1480_
timestamp 1688980957
transform 1 0 23920 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1481_
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1482_
timestamp 1688980957
transform 1 0 30268 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1483_
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1484_
timestamp 1688980957
transform 1 0 20148 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1485_
timestamp 1688980957
transform 1 0 23368 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1486_
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1487_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1488_
timestamp 1688980957
transform 1 0 20056 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1489_
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1490_
timestamp 1688980957
transform 1 0 5336 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1491_
timestamp 1688980957
transform 1 0 2760 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1492_
timestamp 1688980957
transform 1 0 5060 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1493_
timestamp 1688980957
transform 1 0 4692 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1494_
timestamp 1688980957
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1688980957
transform 1 0 3496 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1496_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _1497_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1498_
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1500_
timestamp 1688980957
transform 1 0 14996 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1501_
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1688980957
transform 1 0 16100 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1688980957
transform 1 0 17112 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1688980957
transform 1 0 17572 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1505_
timestamp 1688980957
transform 1 0 10212 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1506_
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1688980957
transform 1 0 10672 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1508_
timestamp 1688980957
transform 1 0 11224 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1509_
timestamp 1688980957
transform 1 0 10580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1510_
timestamp 1688980957
transform 1 0 10948 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1511_
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1512_
timestamp 1688980957
transform 1 0 10396 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 1688980957
transform 1 0 13248 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1514_
timestamp 1688980957
transform 1 0 10948 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1515_
timestamp 1688980957
transform 1 0 12420 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1516_
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1517_
timestamp 1688980957
transform 1 0 12420 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1518_
timestamp 1688980957
transform 1 0 11776 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1519_
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1520_
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1521_
timestamp 1688980957
transform 1 0 11868 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1522_
timestamp 1688980957
transform 1 0 11776 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1523_
timestamp 1688980957
transform 1 0 12972 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1524_
timestamp 1688980957
transform 1 0 12420 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1525_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1527_
timestamp 1688980957
transform 1 0 9568 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1528_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1529_
timestamp 1688980957
transform 1 0 5060 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1530_
timestamp 1688980957
transform 1 0 8740 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1531_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1532_
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1533_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1688980957
transform 1 0 7544 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1535_
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1536_
timestamp 1688980957
transform 1 0 5060 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1537_
timestamp 1688980957
transform 1 0 8464 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1538_
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 1688980957
transform 1 0 9476 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1540_
timestamp 1688980957
transform 1 0 9660 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1541_
timestamp 1688980957
transform 1 0 10580 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1542_
timestamp 1688980957
transform 1 0 10948 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1544_
timestamp 1688980957
transform 1 0 8832 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1545_
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1546_
timestamp 1688980957
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1547_
timestamp 1688980957
transform 1 0 8188 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1548_
timestamp 1688980957
transform 1 0 10304 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1549_
timestamp 1688980957
transform 1 0 8832 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1550_
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1551_
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1552_
timestamp 1688980957
transform 1 0 23736 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1688980957
transform 1 0 27232 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1554_
timestamp 1688980957
transform 1 0 26772 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1555_
timestamp 1688980957
transform 1 0 28980 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1556_
timestamp 1688980957
transform 1 0 30820 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1557_
timestamp 1688980957
transform 1 0 31280 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1558_
timestamp 1688980957
transform 1 0 33580 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_4  _1559_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16376 0 1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1560_
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1688980957
transform 1 0 10396 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1562_
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 1688980957
transform 1 0 16744 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1565_
timestamp 1688980957
transform 1 0 5428 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 1688980957
transform 1 0 12604 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1568_
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1569_
timestamp 1688980957
transform 1 0 4600 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 1688980957
transform 1 0 4324 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1571_
timestamp 1688980957
transform 1 0 3864 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1688980957
transform 1 0 4968 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1573_
timestamp 1688980957
transform 1 0 5888 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1574_
timestamp 1688980957
transform 1 0 4784 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1575_
timestamp 1688980957
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1576_
timestamp 1688980957
transform 1 0 3956 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1577_
timestamp 1688980957
transform 1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1578_
timestamp 1688980957
transform 1 0 3496 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1579_
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1580_
timestamp 1688980957
transform 1 0 2208 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1688980957
transform 1 0 1840 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1582_
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1583_
timestamp 1688980957
transform 1 0 5060 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1584_
timestamp 1688980957
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 1688980957
transform 1 0 5060 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1586_
timestamp 1688980957
transform 1 0 5060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1587_
timestamp 1688980957
transform 1 0 4416 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1588_
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1589_
timestamp 1688980957
transform 1 0 4692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1590_
timestamp 1688980957
transform 1 0 3404 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1591_
timestamp 1688980957
transform 1 0 2852 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 1688980957
transform 1 0 2668 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1593_
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1594_
timestamp 1688980957
transform 1 0 6716 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1595_
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1596_
timestamp 1688980957
transform 1 0 8096 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1597_
timestamp 1688980957
transform 1 0 6716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1598_
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1599_
timestamp 1688980957
transform 1 0 7268 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1600_
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1601_
timestamp 1688980957
transform 1 0 6440 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1602_
timestamp 1688980957
transform 1 0 7268 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1603_
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1604_
timestamp 1688980957
transform 1 0 6624 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1605_
timestamp 1688980957
transform 1 0 6992 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1606_
timestamp 1688980957
transform 1 0 6532 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1607_
timestamp 1688980957
transform 1 0 6716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1608_
timestamp 1688980957
transform 1 0 12420 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1610_
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1611_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 1688980957
transform 1 0 10488 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1613_
timestamp 1688980957
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1614_
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1615_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1616_
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1617_
timestamp 1688980957
transform 1 0 10488 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1618_
timestamp 1688980957
transform 1 0 9752 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1619_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _1620_
timestamp 1688980957
transform 1 0 8464 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1621_
timestamp 1688980957
transform 1 0 8832 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1622_
timestamp 1688980957
transform 1 0 9200 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1688980957
transform 1 0 9476 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1624_
timestamp 1688980957
transform 1 0 9292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1625_
timestamp 1688980957
transform 1 0 10120 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1626_
timestamp 1688980957
transform 1 0 9568 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1627_
timestamp 1688980957
transform 1 0 8924 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1628_
timestamp 1688980957
transform 1 0 9292 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1688980957
transform 1 0 11684 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_4  _1631_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_1  _1632_
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1634_
timestamp 1688980957
transform 1 0 12696 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1635_
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 1688980957
transform 1 0 11316 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1637_
timestamp 1688980957
transform 1 0 10672 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1638_
timestamp 1688980957
transform 1 0 12052 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1639_
timestamp 1688980957
transform 1 0 10856 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1640_
timestamp 1688980957
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1642_
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1643_
timestamp 1688980957
transform 1 0 13524 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1644_
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1645_
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1646_
timestamp 1688980957
transform 1 0 12880 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1647_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1648_
timestamp 1688980957
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1649_
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1650_
timestamp 1688980957
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1651_
timestamp 1688980957
transform 1 0 11592 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1688980957
transform 1 0 12696 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1688980957
transform 1 0 12144 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1654_
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1655_
timestamp 1688980957
transform 1 0 11868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _1656_
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1657_
timestamp 1688980957
transform 1 0 11960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1658_
timestamp 1688980957
transform 1 0 9936 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1659_
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1660_
timestamp 1688980957
transform 1 0 10028 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1661_
timestamp 1688980957
transform 1 0 9200 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1662_
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1663_
timestamp 1688980957
transform 1 0 10304 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1665_
timestamp 1688980957
transform 1 0 8464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1666_
timestamp 1688980957
transform 1 0 9292 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1667_
timestamp 1688980957
transform 1 0 8740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1668_
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1669_
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1670_
timestamp 1688980957
transform 1 0 8372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1671_
timestamp 1688980957
transform 1 0 7820 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1672_
timestamp 1688980957
transform 1 0 7176 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1673_
timestamp 1688980957
transform 1 0 7820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1674_
timestamp 1688980957
transform 1 0 7728 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1675_
timestamp 1688980957
transform 1 0 6808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1688980957
transform 1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1677_
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1678_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1679_
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1680_
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1681_
timestamp 1688980957
transform 1 0 7360 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1682_
timestamp 1688980957
transform 1 0 1840 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1683_
timestamp 1688980957
transform 1 0 3680 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1684_
timestamp 1688980957
transform 1 0 5152 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1685_
timestamp 1688980957
transform 1 0 1472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1686_
timestamp 1688980957
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1687_
timestamp 1688980957
transform 1 0 2852 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1688_
timestamp 1688980957
transform 1 0 2944 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1689_
timestamp 1688980957
transform 1 0 5060 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1690_
timestamp 1688980957
transform 1 0 2392 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1691_
timestamp 1688980957
transform 1 0 5520 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1693_
timestamp 1688980957
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1694_
timestamp 1688980957
transform 1 0 5704 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1695_
timestamp 1688980957
transform 1 0 4600 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _1696_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1697_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1698_
timestamp 1688980957
transform 1 0 4508 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1699_
timestamp 1688980957
transform 1 0 3680 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1700_
timestamp 1688980957
transform 1 0 7912 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1701_
timestamp 1688980957
transform 1 0 12512 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1702_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1704_
timestamp 1688980957
transform 1 0 9660 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1705_
timestamp 1688980957
transform 1 0 7636 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1706_
timestamp 1688980957
transform 1 0 7912 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1707_
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1708_
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1709_
timestamp 1688980957
transform 1 0 6808 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1710_
timestamp 1688980957
transform 1 0 4784 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1712_
timestamp 1688980957
transform 1 0 2852 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1688980957
transform 1 0 2668 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1714_
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1715_
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1716_
timestamp 1688980957
transform 1 0 15272 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _1717_
timestamp 1688980957
transform 1 0 15088 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1718_
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1719_
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1720_
timestamp 1688980957
transform 1 0 13616 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1721_
timestamp 1688980957
transform 1 0 14536 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1722_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1723_
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1724_
timestamp 1688980957
transform 1 0 21160 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1725_
timestamp 1688980957
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1726_
timestamp 1688980957
transform 1 0 17204 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1727_
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1728_
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1729_
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1730_
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _1731_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1732_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1733_
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1734_
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1735_
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1736_
timestamp 1688980957
transform 1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1737_
timestamp 1688980957
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1738_
timestamp 1688980957
transform 1 0 15548 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1739_
timestamp 1688980957
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1740_
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1741_
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1742_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1743_
timestamp 1688980957
transform 1 0 11592 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _1744_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2_1  _1745_
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1746_
timestamp 1688980957
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1747_
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1748_
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1749_
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1750_
timestamp 1688980957
transform 1 0 9568 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1751_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1752_
timestamp 1688980957
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1688980957
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1754_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1755_
timestamp 1688980957
transform 1 0 8372 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1756_
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1757_
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1758_
timestamp 1688980957
transform 1 0 6992 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1759_
timestamp 1688980957
transform 1 0 7360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1760_
timestamp 1688980957
transform 1 0 7728 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1761_
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1762_
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1764_
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1765_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1766_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1767_
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1768_
timestamp 1688980957
transform 1 0 5152 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1769_
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1770_
timestamp 1688980957
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1771_
timestamp 1688980957
transform 1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1772_
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1773_
timestamp 1688980957
transform 1 0 4324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1774_
timestamp 1688980957
transform 1 0 13064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1775_
timestamp 1688980957
transform 1 0 14628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1776_
timestamp 1688980957
transform 1 0 11316 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1777_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1778_
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1779_
timestamp 1688980957
transform 1 0 12696 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1780_
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1781_
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1782_
timestamp 1688980957
transform 1 0 10948 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _1783_
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1784_
timestamp 1688980957
transform 1 0 8740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1785_
timestamp 1688980957
transform 1 0 10948 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1786_
timestamp 1688980957
transform 1 0 12236 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1787_
timestamp 1688980957
transform 1 0 10212 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1788_
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _1789_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1791_
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1792_
timestamp 1688980957
transform 1 0 10396 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1793_
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1794_
timestamp 1688980957
transform 1 0 9936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _1795_
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1796_
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1797_
timestamp 1688980957
transform 1 0 9292 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1798_
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1799_
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1800_
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _1801_
timestamp 1688980957
transform 1 0 6256 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1802_
timestamp 1688980957
transform 1 0 6440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1803_
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1804_
timestamp 1688980957
transform 1 0 7728 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1805_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1806_
timestamp 1688980957
transform 1 0 1472 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _1807_
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1808_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _1809_
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1810_
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1811_
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1812_
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _1813_
timestamp 1688980957
transform 1 0 4048 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1814_
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1815_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1816_
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1817_
timestamp 1688980957
transform 1 0 4416 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1818_
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1819_
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1820_
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1821_
timestamp 1688980957
transform 1 0 18952 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1822_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1823_
timestamp 1688980957
transform 1 0 20608 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1824_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1825_
timestamp 1688980957
transform 1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1826_
timestamp 1688980957
transform 1 0 18952 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1827_
timestamp 1688980957
transform 1 0 17940 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1828_
timestamp 1688980957
transform 1 0 18400 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1829_
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1830_
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_4  _1831_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1832_
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1833_
timestamp 1688980957
transform 1 0 1564 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1834_
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1835_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1836_
timestamp 1688980957
transform 1 0 3128 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1837_
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1838_
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1839_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1840_
timestamp 1688980957
transform 1 0 3220 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1841_
timestamp 1688980957
transform 1 0 5428 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1842_
timestamp 1688980957
transform 1 0 1472 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1843_
timestamp 1688980957
transform 1 0 4508 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1845_
timestamp 1688980957
transform 1 0 2852 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1847_
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1848_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1849_
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1850_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1851_
timestamp 1688980957
transform 1 0 10580 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1852_
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1853_
timestamp 1688980957
transform 1 0 10948 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1855_
timestamp 1688980957
transform 1 0 8096 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1856_
timestamp 1688980957
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1857_
timestamp 1688980957
transform 1 0 6808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1858_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1859_
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1860_
timestamp 1688980957
transform 1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1861_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1862_
timestamp 1688980957
transform 1 0 5704 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1863_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1864_
timestamp 1688980957
transform 1 0 21344 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1865_
timestamp 1688980957
transform 1 0 20884 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1866_
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1867_
timestamp 1688980957
transform 1 0 25116 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1868_
timestamp 1688980957
transform 1 0 31832 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1870_
timestamp 1688980957
transform 1 0 31280 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1871_
timestamp 1688980957
transform 1 0 20240 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1872_
timestamp 1688980957
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1873_
timestamp 1688980957
transform 1 0 30268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1874_
timestamp 1688980957
transform 1 0 23092 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1875_
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1876_
timestamp 1688980957
transform -1 0 25208 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1877_
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1878_
timestamp 1688980957
transform 1 0 23000 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1879_
timestamp 1688980957
transform 1 0 23828 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1880_
timestamp 1688980957
transform 1 0 28980 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1881_
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1882_
timestamp 1688980957
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1883_
timestamp 1688980957
transform 1 0 17204 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_2  _1884_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1885_
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1886_
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1887_
timestamp 1688980957
transform 1 0 15364 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1888_
timestamp 1688980957
transform 1 0 14536 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1889_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1890_
timestamp 1688980957
transform 1 0 15088 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1891_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1892_
timestamp 1688980957
transform 1 0 15272 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1893_
timestamp 1688980957
transform 1 0 17020 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1894_
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1895_
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1896_
timestamp 1688980957
transform 1 0 15088 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1897_
timestamp 1688980957
transform 1 0 15272 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1898_
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1899_
timestamp 1688980957
transform 1 0 21344 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1900_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1901_
timestamp 1688980957
transform 1 0 20516 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1902_
timestamp 1688980957
transform 1 0 20240 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1903_
timestamp 1688980957
transform 1 0 19596 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1904_
timestamp 1688980957
transform 1 0 19596 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1905_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1906_
timestamp 1688980957
transform 1 0 18584 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1688980957
transform 1 0 18032 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1908_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1909_
timestamp 1688980957
transform 1 0 17204 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1910_
timestamp 1688980957
transform 1 0 5612 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1911_
timestamp 1688980957
transform 1 0 14076 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1912_
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1913_
timestamp 1688980957
transform 1 0 14996 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1914_
timestamp 1688980957
transform 1 0 14076 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1915_
timestamp 1688980957
transform 1 0 17848 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1916_
timestamp 1688980957
transform 1 0 15088 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1917_
timestamp 1688980957
transform 1 0 15180 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1918_
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1919_
timestamp 1688980957
transform 1 0 27048 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1920_
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1921_
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1922_
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1923_
timestamp 1688980957
transform 1 0 23092 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1924_
timestamp 1688980957
transform 1 0 25484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1925_
timestamp 1688980957
transform 1 0 26404 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1926_
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1927_
timestamp 1688980957
transform 1 0 21804 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1928_
timestamp 1688980957
transform 1 0 24380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1929_
timestamp 1688980957
transform 1 0 28244 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1930_
timestamp 1688980957
transform 1 0 29072 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1931_
timestamp 1688980957
transform 1 0 24564 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1932_
timestamp 1688980957
transform 1 0 27692 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1688980957
transform 1 0 29992 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1934_
timestamp 1688980957
transform 1 0 30544 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1935_
timestamp 1688980957
transform 1 0 28520 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1936_
timestamp 1688980957
transform 1 0 29624 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1937_
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1938_
timestamp 1688980957
transform 1 0 30268 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1939_
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1940_
timestamp 1688980957
transform 1 0 24840 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1941_
timestamp 1688980957
transform 1 0 33396 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1942_
timestamp 1688980957
transform 1 0 14996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1943_
timestamp 1688980957
transform 1 0 28704 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1944_
timestamp 1688980957
transform 1 0 28888 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1945_
timestamp 1688980957
transform 1 0 28980 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1946_
timestamp 1688980957
transform 1 0 25944 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1947_
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1948_
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1949_
timestamp 1688980957
transform 1 0 24840 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1950_
timestamp 1688980957
transform 1 0 28060 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1951_
timestamp 1688980957
transform 1 0 25760 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1952_
timestamp 1688980957
transform 1 0 25668 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1953_
timestamp 1688980957
transform 1 0 26864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1954_
timestamp 1688980957
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1955_
timestamp 1688980957
transform 1 0 26036 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1956_
timestamp 1688980957
transform 1 0 28428 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1957_
timestamp 1688980957
transform 1 0 27324 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1958_
timestamp 1688980957
transform 1 0 25944 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1959_
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1960_
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1961_
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1962_
timestamp 1688980957
transform 1 0 27232 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1963_
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1964_
timestamp 1688980957
transform 1 0 26036 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1965_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1966_
timestamp 1688980957
transform 1 0 20700 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1967_
timestamp 1688980957
transform 1 0 25484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1968_
timestamp 1688980957
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1969_
timestamp 1688980957
transform 1 0 22264 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1970_
timestamp 1688980957
transform 1 0 23000 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1971_
timestamp 1688980957
transform 1 0 27600 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1972_
timestamp 1688980957
transform 1 0 28336 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1973_
timestamp 1688980957
transform 1 0 28060 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1974_
timestamp 1688980957
transform 1 0 27876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1975_
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1976_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1977_
timestamp 1688980957
transform 1 0 27692 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1978_
timestamp 1688980957
transform 1 0 25116 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1979_
timestamp 1688980957
transform 1 0 19412 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1980_
timestamp 1688980957
transform 1 0 27416 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1981_
timestamp 1688980957
transform 1 0 26680 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1982_
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1983_
timestamp 1688980957
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1984_
timestamp 1688980957
transform 1 0 24748 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1985_
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1986_
timestamp 1688980957
transform 1 0 28520 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1987_
timestamp 1688980957
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1988_
timestamp 1688980957
transform 1 0 29440 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1989_
timestamp 1688980957
transform 1 0 29624 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1990_
timestamp 1688980957
transform 1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1991_
timestamp 1688980957
transform 1 0 28796 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1992_
timestamp 1688980957
transform 1 0 29992 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1993_
timestamp 1688980957
transform 1 0 30544 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1994_
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1995_
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1996_
timestamp 1688980957
transform 1 0 21068 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1997_
timestamp 1688980957
transform 1 0 19412 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1998_
timestamp 1688980957
transform 1 0 19688 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1999_
timestamp 1688980957
transform 1 0 18400 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2000_
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2001_
timestamp 1688980957
transform 1 0 28612 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2002_
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2003_
timestamp 1688980957
transform 1 0 29348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2004_
timestamp 1688980957
transform 1 0 26496 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2005_
timestamp 1688980957
transform 1 0 25668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2006_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2007_
timestamp 1688980957
transform 1 0 22264 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2008_
timestamp 1688980957
transform 1 0 25024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2009_
timestamp 1688980957
transform 1 0 20332 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2010_
timestamp 1688980957
transform 1 0 20700 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2011_
timestamp 1688980957
transform 1 0 30084 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2012_
timestamp 1688980957
transform 1 0 32200 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2013_
timestamp 1688980957
transform 1 0 22724 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2014_
timestamp 1688980957
transform 1 0 20884 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _2015_
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2016_
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2017_
timestamp 1688980957
transform 1 0 24472 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2018_
timestamp 1688980957
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2019_
timestamp 1688980957
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2020_
timestamp 1688980957
transform 1 0 24472 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2021_
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2022_
timestamp 1688980957
transform 1 0 24196 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2023_
timestamp 1688980957
transform 1 0 23368 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2024_
timestamp 1688980957
transform 1 0 19780 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2025_
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2026_
timestamp 1688980957
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2027_
timestamp 1688980957
transform 1 0 19412 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2028_
timestamp 1688980957
transform 1 0 21252 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2029_
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2030_
timestamp 1688980957
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2031_
timestamp 1688980957
transform 1 0 30084 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2032_
timestamp 1688980957
transform 1 0 30084 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2033_
timestamp 1688980957
transform 1 0 32660 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2034_
timestamp 1688980957
transform 1 0 30452 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2035_
timestamp 1688980957
transform 1 0 33396 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2036_
timestamp 1688980957
transform 1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2037_
timestamp 1688980957
transform 1 0 29900 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2038_
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2039_
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2040_
timestamp 1688980957
transform 1 0 33580 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2041_
timestamp 1688980957
transform 1 0 30636 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2042_
timestamp 1688980957
transform 1 0 33488 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2043_
timestamp 1688980957
transform 1 0 29716 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2044_
timestamp 1688980957
transform 1 0 32752 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2045_
timestamp 1688980957
transform 1 0 30084 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2046_
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2047_
timestamp 1688980957
transform 1 0 33580 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2048_
timestamp 1688980957
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2049_
timestamp 1688980957
transform 1 0 28244 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2050_
timestamp 1688980957
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2051_
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2052_
timestamp 1688980957
transform 1 0 17572 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2053_
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2054_
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2055_
timestamp 1688980957
transform 1 0 32108 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2056_
timestamp 1688980957
transform 1 0 32384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2057_
timestamp 1688980957
transform 1 0 30452 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_4  _2058_
timestamp 1688980957
transform 1 0 15180 0 -1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2059_
timestamp 1688980957
transform 1 0 18124 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2060_
timestamp 1688980957
transform 1 0 10488 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2061_
timestamp 1688980957
transform 1 0 15088 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2062_
timestamp 1688980957
transform 1 0 18124 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2063_
timestamp 1688980957
transform 1 0 8004 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2064_
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2065_
timestamp 1688980957
transform 1 0 11868 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2066_
timestamp 1688980957
transform 1 0 8188 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_4  _2067_
timestamp 1688980957
transform 1 0 16836 0 -1 36992
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2068_
timestamp 1688980957
transform 1 0 16468 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2069_
timestamp 1688980957
transform 1 0 12144 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2070_
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2071_
timestamp 1688980957
transform 1 0 15088 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2072_
timestamp 1688980957
transform 1 0 4600 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2073_
timestamp 1688980957
transform 1 0 4600 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2074_
timestamp 1688980957
transform 1 0 12696 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2075_
timestamp 1688980957
transform 1 0 9108 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2076_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2077_
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2078_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2079_
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2080_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2081_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2082_
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2083_
timestamp 1688980957
transform 1 0 17296 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2084_
timestamp 1688980957
transform 1 0 9844 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2085_
timestamp 1688980957
transform 1 0 14628 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2086_
timestamp 1688980957
transform 1 0 14628 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2087_
timestamp 1688980957
transform 1 0 4232 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2088_
timestamp 1688980957
transform 1 0 4140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2089_
timestamp 1688980957
transform 1 0 12696 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2090_
timestamp 1688980957
transform 1 0 7360 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2091_
timestamp 1688980957
transform 1 0 24196 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2092_
timestamp 1688980957
transform 1 0 22632 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2093_
timestamp 1688980957
transform 1 0 27600 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2094_
timestamp 1688980957
transform 1 0 26036 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2095_
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2096_
timestamp 1688980957
transform 1 0 29072 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2097_
timestamp 1688980957
transform 1 0 31004 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2098_
timestamp 1688980957
transform 1 0 31924 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2099_
timestamp 1688980957
transform 1 0 18492 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2100_
timestamp 1688980957
transform 1 0 9844 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2101_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2102_
timestamp 1688980957
transform 1 0 16560 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2103_
timestamp 1688980957
transform 1 0 5704 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2104_
timestamp 1688980957
transform 1 0 6992 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2105_
timestamp 1688980957
transform 1 0 12144 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2106_
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2107_
timestamp 1688980957
transform 1 0 20240 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2108_
timestamp 1688980957
transform 1 0 1656 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2109_
timestamp 1688980957
transform 1 0 6348 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2110_
timestamp 1688980957
transform 1 0 13156 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2111_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _2112_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 -1 31552
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _2113_
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2114_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2115_
timestamp 1688980957
transform 1 0 4600 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2116_
timestamp 1688980957
transform 1 0 4600 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2117_
timestamp 1688980957
transform 1 0 1932 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2118_
timestamp 1688980957
transform 1 0 1840 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2119_
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2120_
timestamp 1688980957
transform 1 0 14444 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2121_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2122_
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2123_
timestamp 1688980957
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2124_
timestamp 1688980957
transform 1 0 5888 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2125_
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2126_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2127_
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2128_
timestamp 1688980957
transform 1 0 9292 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2129_
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2130_
timestamp 1688980957
transform 1 0 7360 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2131_
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2132_
timestamp 1688980957
transform 1 0 2300 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2133_
timestamp 1688980957
transform 1 0 2024 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2134_
timestamp 1688980957
transform 1 0 2576 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2135_
timestamp 1688980957
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2136_
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2137_
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2138_
timestamp 1688980957
transform 1 0 1840 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2139_
timestamp 1688980957
transform 1 0 1748 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2149_
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1688980957
transform 1 0 16376 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1688980957
transform 1 0 29348 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1688980957
transform 1 0 30452 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1688980957
transform 1 0 27416 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1688980957
transform 1 0 30176 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1688980957
transform 1 0 20148 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _2160_
timestamp 1688980957
transform 1 0 29440 0 -1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _2161_
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2162_
timestamp 1688980957
transform 1 0 14996 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2163_
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2164_
timestamp 1688980957
transform 1 0 17112 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2165_
timestamp 1688980957
transform 1 0 14812 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2166_
timestamp 1688980957
transform 1 0 22724 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1688980957
transform 1 0 24932 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1688980957
transform 1 0 22448 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2169_
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1688980957
transform 1 0 25208 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1688980957
transform 1 0 29992 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1688980957
transform 1 0 27416 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2173_
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2175_
timestamp 1688980957
transform 1 0 32384 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2177_
timestamp 1688980957
transform 1 0 22540 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2178_
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1688980957
transform 1 0 21988 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1688980957
transform 1 0 20884 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1688980957
transform 1 0 19596 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2182_
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2183_
timestamp 1688980957
transform 1 0 22816 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1688980957
transform 1 0 29072 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2185_
timestamp 1688980957
transform 1 0 29808 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1688980957
transform 1 0 19596 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2188_
timestamp 1688980957
transform 1 0 17940 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2189_
timestamp 1688980957
transform 1 0 29624 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2190_
timestamp 1688980957
transform 1 0 22080 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2191_
timestamp 1688980957
transform 1 0 19780 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2192_
timestamp 1688980957
transform 1 0 30820 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2193_
timestamp 1688980957
transform 1 0 19688 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2194_
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2195_
timestamp 1688980957
transform 1 0 17664 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2196_
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2197_
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2198_
timestamp 1688980957
transform 1 0 30544 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2199_
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2200_
timestamp 1688980957
transform 1 0 30176 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2201_
timestamp 1688980957
transform 1 0 32016 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2202_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2203_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2204_
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2205_
timestamp 1688980957
transform 1 0 28704 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2206_
timestamp 1688980957
transform 1 0 29532 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2207_
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2208_
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2209_
timestamp 1688980957
transform 1 0 17204 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2210_
timestamp 1688980957
transform 1 0 30912 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2211_
timestamp 1688980957
transform 1 0 17664 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2212_
timestamp 1688980957
transform 1 0 9844 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2213_
timestamp 1688980957
transform 1 0 14720 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2214_
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2215_
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2216_
timestamp 1688980957
transform 1 0 5520 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2217_
timestamp 1688980957
transform 1 0 12144 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2218_
timestamp 1688980957
transform 1 0 7544 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2219_
timestamp 1688980957
transform 1 0 16836 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2220_
timestamp 1688980957
transform 1 0 9752 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2221_
timestamp 1688980957
transform 1 0 11960 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2222_
timestamp 1688980957
transform 1 0 14628 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2223_
timestamp 1688980957
transform 1 0 4232 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2224_
timestamp 1688980957
transform 1 0 4140 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2225_
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2226_
timestamp 1688980957
transform 1 0 7636 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25576 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1688980957
transform 1 0 16928 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B
timestamp 1688980957
transform 1 0 18308 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__D
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A2
timestamp 1688980957
transform 1 0 18216 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A2
timestamp 1688980957
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1688980957
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__S
timestamp 1688980957
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B2
timestamp 1688980957
transform 1 0 7360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__B2
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__S
timestamp 1688980957
transform 1 0 33580 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B2
timestamp 1688980957
transform 1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__S
timestamp 1688980957
transform 1 0 33028 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__B2
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__S
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__B2
timestamp 1688980957
transform 1 0 8280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__S
timestamp 1688980957
transform 1 0 30912 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B2
timestamp 1688980957
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__S
timestamp 1688980957
transform 1 0 31280 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B2
timestamp 1688980957
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A1
timestamp 1688980957
transform 1 0 11776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__S
timestamp 1688980957
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B2
timestamp 1688980957
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__S
timestamp 1688980957
transform 1 0 27140 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1688980957
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A2
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A1
timestamp 1688980957
transform 1 0 3220 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A2
timestamp 1688980957
transform 1 0 5796 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A2
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A2
timestamp 1688980957
transform 1 0 8188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A2
timestamp 1688980957
transform 1 0 7912 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1
timestamp 1688980957
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A2
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A2
timestamp 1688980957
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A2
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1688980957
transform 1 0 16100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1688980957
transform 1 0 24840 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__C1
timestamp 1688980957
transform 1 0 41860 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__B
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B
timestamp 1688980957
transform 1 0 25208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1688980957
transform 1 0 23092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B2
timestamp 1688980957
transform 1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1
timestamp 1688980957
transform 1 0 15364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1688980957
transform 1 0 15180 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A0
timestamp 1688980957
transform 1 0 31924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 1688980957
transform 1 0 26496 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A0
timestamp 1688980957
transform 1 0 30912 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1688980957
transform 1 0 28428 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A
timestamp 1688980957
transform 1 0 28888 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A0
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A
timestamp 1688980957
transform 1 0 25208 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A
timestamp 1688980957
transform 1 0 26588 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A0
timestamp 1688980957
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1688980957
transform 1 0 24840 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A0
timestamp 1688980957
transform 1 0 32660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A0
timestamp 1688980957
transform 1 0 32292 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A
timestamp 1688980957
transform 1 0 27876 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1688980957
transform 1 0 27508 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A0
timestamp 1688980957
transform 1 0 22264 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1688980957
transform 1 0 23276 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A0
timestamp 1688980957
transform 1 0 33028 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A
timestamp 1688980957
transform 1 0 31740 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A
timestamp 1688980957
transform 1 0 29256 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1688980957
transform 1 0 29072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1688980957
transform 1 0 25576 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1688980957
transform 1 0 24380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A1
timestamp 1688980957
transform 1 0 25300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__B
timestamp 1688980957
transform 1 0 18308 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__B2
timestamp 1688980957
transform 1 0 23460 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B1
timestamp 1688980957
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1688980957
transform 1 0 27232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A0
timestamp 1688980957
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A1
timestamp 1688980957
transform 1 0 18676 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A2
timestamp 1688980957
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A3
timestamp 1688980957
transform 1 0 15824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__B
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__B
timestamp 1688980957
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__B1
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__A1
timestamp 1688980957
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A1
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__B2
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__B2
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__B2
timestamp 1688980957
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__B2
timestamp 1688980957
transform 1 0 10488 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B2
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1688980957
transform 1 0 16468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__B2
timestamp 1688980957
transform 1 0 6532 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__B2
timestamp 1688980957
transform 1 0 7912 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__B2
timestamp 1688980957
transform 1 0 6992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__B
timestamp 1688980957
transform 1 0 13432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__B
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A2
timestamp 1688980957
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__A2
timestamp 1688980957
transform 1 0 14720 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__D
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__C
timestamp 1688980957
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A2
timestamp 1688980957
transform 1 0 4416 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__B2
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A2
timestamp 1688980957
transform 1 0 22724 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__C
timestamp 1688980957
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__B
timestamp 1688980957
transform 1 0 14168 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__A2
timestamp 1688980957
transform 1 0 3220 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__B1
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__A1
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__B1
timestamp 1688980957
transform 1 0 23736 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A2
timestamp 1688980957
transform 1 0 31280 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__B1
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1688980957
transform 1 0 22724 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__S
timestamp 1688980957
transform 1 0 1840 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__C
timestamp 1688980957
transform 1 0 17480 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A1
timestamp 1688980957
transform 1 0 15088 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__B1
timestamp 1688980957
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__A
timestamp 1688980957
transform 1 0 20516 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__A
timestamp 1688980957
transform 1 0 11684 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__A
timestamp 1688980957
transform 1 0 13156 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__B
timestamp 1688980957
transform 1 0 13524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A2
timestamp 1688980957
transform 1 0 15824 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__B1
timestamp 1688980957
transform 1 0 10488 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__A1
timestamp 1688980957
transform 1 0 10396 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__A2
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__A
timestamp 1688980957
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A
timestamp 1688980957
transform 1 0 10856 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A
timestamp 1688980957
transform 1 0 10856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__B
timestamp 1688980957
transform 1 0 10396 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__A1
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1688980957
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__B1
timestamp 1688980957
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__A1
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__A2
timestamp 1688980957
transform 1 0 11592 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__A
timestamp 1688980957
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__B
timestamp 1688980957
transform 1 0 10212 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__A2
timestamp 1688980957
transform 1 0 8004 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1530__B
timestamp 1688980957
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__A1
timestamp 1688980957
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__A
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A1
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A2
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__A0
timestamp 1688980957
transform 1 0 10120 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__S
timestamp 1688980957
transform 1 0 9568 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__A
timestamp 1688980957
transform 1 0 11684 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__B
timestamp 1688980957
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__A1
timestamp 1688980957
transform 1 0 8280 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__A
timestamp 1688980957
transform 1 0 7360 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__A1
timestamp 1688980957
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__A2
timestamp 1688980957
transform 1 0 7176 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__B1
timestamp 1688980957
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__S
timestamp 1688980957
transform 1 0 20700 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__A2
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__B1
timestamp 1688980957
transform 1 0 4048 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__A2
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__B2
timestamp 1688980957
transform 1 0 5428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A2
timestamp 1688980957
transform 1 0 6808 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__B1
timestamp 1688980957
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A2
timestamp 1688980957
transform 1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__B2
timestamp 1688980957
transform 1 0 4784 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__A2
timestamp 1688980957
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__B1
timestamp 1688980957
transform 1 0 7912 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__A2
timestamp 1688980957
transform 1 0 8648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__B2
timestamp 1688980957
transform 1 0 7912 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__A2
timestamp 1688980957
transform 1 0 10212 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__B1
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__A1
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__A2
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__B2
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__A2
timestamp 1688980957
transform 1 0 9844 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__B1
timestamp 1688980957
transform 1 0 8280 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__B1
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__A2
timestamp 1688980957
transform 1 0 14260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__B2
timestamp 1688980957
transform 1 0 13248 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A2
timestamp 1688980957
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B1
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__A2
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__B2
timestamp 1688980957
transform 1 0 14444 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1664__A2
timestamp 1688980957
transform 1 0 9752 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1664__B2
timestamp 1688980957
transform 1 0 9384 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1678__C1
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__C1
timestamp 1688980957
transform 1 0 5520 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1699__A0
timestamp 1688980957
transform 1 0 3956 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1699__S
timestamp 1688980957
transform 1 0 4324 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1700__S
timestamp 1688980957
transform 1 0 10304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1702__S
timestamp 1688980957
transform 1 0 12696 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1703__S
timestamp 1688980957
transform 1 0 10948 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1704__S
timestamp 1688980957
transform 1 0 10120 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1705__A
timestamp 1688980957
transform 1 0 7912 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1706__A1
timestamp 1688980957
transform 1 0 8280 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1706__A2
timestamp 1688980957
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__A
timestamp 1688980957
transform 1 0 6532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1709__B2
timestamp 1688980957
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1710__S
timestamp 1688980957
transform 1 0 5796 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1711__S
timestamp 1688980957
transform 1 0 4416 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1712__A0
timestamp 1688980957
transform 1 0 6164 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1712__S
timestamp 1688980957
transform 1 0 1932 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__S
timestamp 1688980957
transform 1 0 3128 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1717__A
timestamp 1688980957
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1717__B
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1718__A
timestamp 1688980957
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1718__B
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1720__B
timestamp 1688980957
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1722__B1
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1728__B
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1729__B1
timestamp 1688980957
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1731__A2
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1738__A1
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1740__A
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1743__A1
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1744__A1
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__B1
timestamp 1688980957
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1750__A1
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1752__B1
timestamp 1688980957
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1756__A1
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1758__B1
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1762__A1
timestamp 1688980957
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1764__B1
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1768__A1
timestamp 1688980957
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__A1
timestamp 1688980957
transform 1 0 5888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__C1
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1773__A1
timestamp 1688980957
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1776__A
timestamp 1688980957
transform 1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1777__A2
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1777__C1
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1778__A
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1781__A1
timestamp 1688980957
transform 1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1783__A2
timestamp 1688980957
transform 1 0 10580 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1783__C1
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1784__A
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1787__A1
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1789__A1
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1789__A2
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1789__C1
timestamp 1688980957
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1790__A
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1793__A1
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1795__A2
timestamp 1688980957
transform 1 0 7544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1795__C1
timestamp 1688980957
transform 1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1796__A
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1799__A1
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1801__A2
timestamp 1688980957
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1801__C1
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__A
timestamp 1688980957
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1805__A1
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1807__A2
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1807__C1
timestamp 1688980957
transform 1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1808__A
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__A1
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1812__A2
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1812__C1
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1813__A1
timestamp 1688980957
transform 1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1815__B1_N
timestamp 1688980957
transform 1 0 1564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A1
timestamp 1688980957
transform 1 0 4416 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A2
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__C1
timestamp 1688980957
transform 1 0 6624 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1818__A1
timestamp 1688980957
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1820__B2
timestamp 1688980957
transform 1 0 5428 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1824__B
timestamp 1688980957
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1826__D
timestamp 1688980957
transform 1 0 20516 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1830__A
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1830__D
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1832__S
timestamp 1688980957
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1833__A
timestamp 1688980957
transform 1 0 2024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1834__S
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1835__A
timestamp 1688980957
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1836__S
timestamp 1688980957
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1837__A
timestamp 1688980957
transform 1 0 3680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1838__S
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1839__A
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1840__S
timestamp 1688980957
transform 1 0 4048 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1841__A
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1842__S
timestamp 1688980957
transform 1 0 2024 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1843__A
timestamp 1688980957
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1844__S
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1845__A
timestamp 1688980957
transform 1 0 4508 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1846__S
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1847__A
timestamp 1688980957
transform 1 0 1656 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__S
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__A
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1850__S
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1851__A
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1852__S
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1853__A
timestamp 1688980957
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1854__S
timestamp 1688980957
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1855__A
timestamp 1688980957
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1856__S
timestamp 1688980957
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1857__A
timestamp 1688980957
transform 1 0 7268 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1858__S
timestamp 1688980957
transform 1 0 7636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1859__A
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1860__S
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1861__A
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1862__S
timestamp 1688980957
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1863__A
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__B
timestamp 1688980957
transform 1 0 21160 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1865__B
timestamp 1688980957
transform 1 0 21344 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1866__B
timestamp 1688980957
transform 1 0 32476 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1868__B
timestamp 1688980957
transform 1 0 32292 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1869__A
timestamp 1688980957
transform 1 0 27876 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1870__A
timestamp 1688980957
transform 1 0 32292 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1870__B
timestamp 1688980957
transform 1 0 32660 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1871__A
timestamp 1688980957
transform 1 0 20884 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1871__B
timestamp 1688980957
transform 1 0 20148 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__A
timestamp 1688980957
transform 1 0 33396 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1876__S
timestamp 1688980957
transform 1 0 26036 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__A1
timestamp 1688980957
transform 1 0 26128 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1878__A1
timestamp 1688980957
transform 1 0 23368 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__A
timestamp 1688980957
transform 1 0 28796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1883__C1
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1886__A2
timestamp 1688980957
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1888__A
timestamp 1688980957
transform 1 0 13248 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1888__D
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1891__B1
timestamp 1688980957
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1893__A2
timestamp 1688980957
transform 1 0 13432 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1895__A
timestamp 1688980957
transform 1 0 14352 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1896__A0
timestamp 1688980957
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1896__A1
timestamp 1688980957
transform 1 0 14352 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1898__A
timestamp 1688980957
transform 1 0 12604 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1899__B2
timestamp 1688980957
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1901__A1
timestamp 1688980957
transform 1 0 19412 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1902__A1
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1904__C1
timestamp 1688980957
transform 1 0 19412 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1905__A1
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1906__A1
timestamp 1688980957
transform 1 0 17020 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1906__S
timestamp 1688980957
transform 1 0 17020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1909__A
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1912__A
timestamp 1688980957
transform 1 0 32568 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1914__B2
timestamp 1688980957
transform 1 0 12420 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1915__A2
timestamp 1688980957
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1916__A0
timestamp 1688980957
transform 1 0 13156 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1916__S
timestamp 1688980957
transform 1 0 12788 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1918__A
timestamp 1688980957
transform 1 0 13892 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1919__A
timestamp 1688980957
transform 1 0 33028 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1919__B
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__A
timestamp 1688980957
transform 1 0 25852 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__B
timestamp 1688980957
transform 1 0 27140 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1921__A
timestamp 1688980957
transform 1 0 21896 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1922__A
timestamp 1688980957
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1922__B
timestamp 1688980957
transform 1 0 25852 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__B1
timestamp 1688980957
transform 1 0 27784 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1926__C1
timestamp 1688980957
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1927__A1
timestamp 1688980957
transform 1 0 22816 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1927__A3
timestamp 1688980957
transform 1 0 22448 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1927__B1
timestamp 1688980957
transform 1 0 22080 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1930__C1
timestamp 1688980957
transform 1 0 33396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1931__A1
timestamp 1688980957
transform 1 0 26220 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1931__A3
timestamp 1688980957
transform 1 0 30544 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1931__B1
timestamp 1688980957
transform 1 0 23552 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1934__C1
timestamp 1688980957
transform 1 0 33028 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1935__A1
timestamp 1688980957
transform 1 0 30176 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1935__A3
timestamp 1688980957
transform 1 0 29256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1935__B1
timestamp 1688980957
transform 1 0 28336 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1937__A1
timestamp 1688980957
transform 1 0 33028 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1937__A3
timestamp 1688980957
transform 1 0 31648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1939__A1
timestamp 1688980957
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1939__A3
timestamp 1688980957
transform 1 0 25760 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1939__B1
timestamp 1688980957
transform 1 0 25024 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1941__A
timestamp 1688980957
transform 1 0 34040 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1941__B
timestamp 1688980957
transform 1 0 34408 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1942__B1
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1969__B1
timestamp 1688980957
transform 1 0 23552 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1975__C1
timestamp 1688980957
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1983__C1
timestamp 1688980957
transform 1 0 27140 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1987__C1
timestamp 1688980957
transform 1 0 29716 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1994__A
timestamp 1688980957
transform 1 0 17480 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2003__A
timestamp 1688980957
transform 1 0 29716 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2014__C1
timestamp 1688980957
transform 1 0 25944 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2023__C1
timestamp 1688980957
transform 1 0 24564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__A
timestamp 1688980957
transform 1 0 34040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2038__C1
timestamp 1688980957
transform 1 0 34224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2045__A
timestamp 1688980957
transform 1 0 29716 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2047__A
timestamp 1688980957
transform 1 0 33764 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2051__A1
timestamp 1688980957
transform 1 0 29256 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2051__C1
timestamp 1688980957
transform 1 0 29624 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2053__B2
timestamp 1688980957
transform 1 0 13248 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2055__C_N
timestamp 1688980957
transform 1 0 32936 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2056__A1
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2057__A
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2058__B1
timestamp 1688980957
transform 1 0 16376 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2067__B1
timestamp 1688980957
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 7820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 4140 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 4048 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 13892 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 35236 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 32752 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 22632 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 21528 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 29164 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_A
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout63_A
timestamp 1688980957
transform 1 0 22448 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout73_A
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_A
timestamp 1688980957
transform 1 0 24288 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp 1688980957
transform 1 0 34500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout76_A
timestamp 1688980957
transform 1 0 34132 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout77_A
timestamp 1688980957
transform 1 0 33396 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_A
timestamp 1688980957
transform 1 0 32660 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold147_A
timestamp 1688980957
transform 1 0 15364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold160_A
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold167_A
timestamp 1688980957
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold191_A
timestamp 1688980957
transform 1 0 4508 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold200_A
timestamp 1688980957
transform 1 0 11500 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold214_A
timestamp 1688980957
transform 1 0 17848 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold217_A
timestamp 1688980957
transform 1 0 34224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold223_A
timestamp 1688980957
transform 1 0 28888 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold225_A
timestamp 1688980957
transform 1 0 22448 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold229_A
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold232_A
timestamp 1688980957
transform 1 0 12052 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold234_A
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold236_A
timestamp 1688980957
transform 1 0 29992 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output15_A
timestamp 1688980957
transform 1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output16_A
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1688980957
transform 1 0 1656 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1688980957
transform 1 0 3036 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1688980957
transform 1 0 3036 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1688980957
transform 1 0 6440 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1688980957
transform 1 0 6808 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1688980957
transform 1 0 7820 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1688980957
transform 1 0 15916 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1688980957
transform 1 0 28060 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1688980957
transform 1 0 35420 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1688980957
transform 1 0 32936 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1688980957
transform 1 0 20700 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1688980957
transform 1 0 28060 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout48 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout52
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout53
timestamp 1688980957
transform 1 0 22264 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout54
timestamp 1688980957
transform 1 0 15548 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout55 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout56
timestamp 1688980957
transform 1 0 22632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout58
timestamp 1688980957
transform 1 0 23644 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout60
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout61
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1688980957
transform 1 0 23092 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1688980957
transform 1 0 23092 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout64
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout65 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout66
timestamp 1688980957
transform 1 0 19780 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout67
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout68
timestamp 1688980957
transform 1 0 20608 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1688980957
transform 1 0 23460 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout70
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout71
timestamp 1688980957
transform 1 0 22448 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout72
timestamp 1688980957
transform 1 0 23092 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout74
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 1688980957
transform 1 0 33396 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout77
timestamp 1688980957
transform 1 0 32844 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout78
timestamp 1688980957
transform 1 0 31096 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout79
timestamp 1688980957
transform 1 0 31464 0 1 38080
box -38 -48 866 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_257
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_19
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1688980957
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_461
timestamp 1688980957
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 1688980957
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_461
timestamp 1688980957
transform 1 0 43516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_19
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_23
timestamp 1688980957
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_461
timestamp 1688980957
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_461
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_461
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_461
timestamp 1688980957
transform 1 0 43516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1688980957
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1688980957
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1688980957
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 1688980957
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1688980957
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_457
timestamp 1688980957
transform 1 0 43148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_461
timestamp 1688980957
transform 1 0 43516 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1688980957
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 1688980957
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 1688980957
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 1688980957
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_461
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_19
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 1688980957
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 1688980957
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_457
timestamp 1688980957
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_461
timestamp 1688980957
transform 1 0 43516 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1688980957
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1688980957
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 1688980957
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 1688980957
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_19
timestamp 1688980957
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1688980957
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1688980957
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1688980957
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_457
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_461
timestamp 1688980957
transform 1 0 43516 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_36
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_48
timestamp 1688980957
transform 1 0 5520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_61
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_73
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_85
timestamp 1688980957
transform 1 0 8924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_97
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1688980957
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 1688980957
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 1688980957
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1688980957
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_461
timestamp 1688980957
transform 1 0 43516 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_19
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_25
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_36
timestamp 1688980957
transform 1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_40
timestamp 1688980957
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_45
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_49
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_54
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_64
timestamp 1688980957
transform 1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_74
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 1688980957
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 1688980957
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 1688980957
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 1688980957
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 1688980957
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_457
timestamp 1688980957
transform 1 0 43148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_461
timestamp 1688980957
transform 1 0 43516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_12
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_26
timestamp 1688980957
transform 1 0 3496 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_34
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_38
timestamp 1688980957
transform 1 0 4600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_46
timestamp 1688980957
transform 1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_74
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_78
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_99
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1688980957
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1688980957
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 1688980957
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 1688980957
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_461
timestamp 1688980957
transform 1 0 43516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_19
timestamp 1688980957
transform 1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_24
timestamp 1688980957
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_34
timestamp 1688980957
transform 1 0 4232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_39
timestamp 1688980957
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_44
timestamp 1688980957
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_90
timestamp 1688980957
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_96
timestamp 1688980957
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_108
timestamp 1688980957
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_114
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_126
timestamp 1688980957
transform 1 0 12696 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_157
timestamp 1688980957
transform 1 0 15548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_169
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_181
timestamp 1688980957
transform 1 0 17756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1688980957
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1688980957
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1688980957
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_461
timestamp 1688980957
transform 1 0 43516 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_8
timestamp 1688980957
transform 1 0 1840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_28
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_102
timestamp 1688980957
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_129
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_152
timestamp 1688980957
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1688980957
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 1688980957
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 1688980957
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 1688980957
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_461
timestamp 1688980957
transform 1 0 43516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_19
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_67
timestamp 1688980957
transform 1 0 7268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_71
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_102
timestamp 1688980957
transform 1 0 10488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_158
timestamp 1688980957
transform 1 0 15640 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_163
timestamp 1688980957
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_167
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_173
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 1688980957
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_217
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1688980957
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 1688980957
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 1688980957
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_457
timestamp 1688980957
transform 1 0 43148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_461
timestamp 1688980957
transform 1 0 43516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_35
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_71
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_79
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_96
timestamp 1688980957
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_100
timestamp 1688980957
transform 1 0 10304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_107
timestamp 1688980957
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_122
timestamp 1688980957
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_127
timestamp 1688980957
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_143
timestamp 1688980957
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1688980957
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_180
timestamp 1688980957
transform 1 0 17664 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_184
timestamp 1688980957
transform 1 0 18032 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_192
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_201
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_207
timestamp 1688980957
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_241
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_253
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_265
timestamp 1688980957
transform 1 0 25484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1688980957
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 1688980957
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1688980957
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1688980957
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 1688980957
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1688980957
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_461
timestamp 1688980957
transform 1 0 43516 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_50
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_88
timestamp 1688980957
transform 1 0 9200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_163
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_167
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_171
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_175
timestamp 1688980957
transform 1 0 17204 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_180
timestamp 1688980957
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_208
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_216
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_220
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_244
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1688980957
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1688980957
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1688980957
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1688980957
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1688980957
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_457
timestamp 1688980957
transform 1 0 43148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_461
timestamp 1688980957
transform 1 0 43516 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_160
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1688980957
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_214
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_255
timestamp 1688980957
transform 1 0 24564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_267
timestamp 1688980957
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1688980957
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 1688980957
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 1688980957
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 1688980957
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_455
timestamp 1688980957
transform 1 0 42964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_64
timestamp 1688980957
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_112
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_123
timestamp 1688980957
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_180
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_224
timestamp 1688980957
transform 1 0 21712 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_237
timestamp 1688980957
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_261
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_280
timestamp 1688980957
transform 1 0 26864 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_292
timestamp 1688980957
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_304
timestamp 1688980957
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 1688980957
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 1688980957
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1688980957
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_457
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_461
timestamp 1688980957
transform 1 0 43516 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_31
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_42
timestamp 1688980957
transform 1 0 4968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_71
timestamp 1688980957
transform 1 0 7636 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_77
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_91
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_101
timestamp 1688980957
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_108
timestamp 1688980957
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_153
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_202
timestamp 1688980957
transform 1 0 19688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_212
timestamp 1688980957
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_248
timestamp 1688980957
transform 1 0 23920 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_272
timestamp 1688980957
transform 1 0 26128 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_298
timestamp 1688980957
transform 1 0 28520 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_310
timestamp 1688980957
transform 1 0 29624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_322
timestamp 1688980957
transform 1 0 30728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_334
timestamp 1688980957
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 1688980957
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1688980957
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 1688980957
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 1688980957
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 1688980957
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_69
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_72
timestamp 1688980957
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_76
timestamp 1688980957
transform 1 0 8096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_80
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_89
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_105
timestamp 1688980957
transform 1 0 10764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_118
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_123
timestamp 1688980957
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_163
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_174
timestamp 1688980957
transform 1 0 17112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_256
timestamp 1688980957
transform 1 0 24656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_260
timestamp 1688980957
transform 1 0 25024 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_285
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 1688980957
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 1688980957
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1688980957
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 1688980957
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_457
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_461
timestamp 1688980957
transform 1 0 43516 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_60
timestamp 1688980957
transform 1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_68
timestamp 1688980957
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_94
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_109
timestamp 1688980957
transform 1 0 11132 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_152
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_172
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_215
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1688980957
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_236
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_255
timestamp 1688980957
transform 1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_265
timestamp 1688980957
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1688980957
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_300
timestamp 1688980957
transform 1 0 28704 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_312
timestamp 1688980957
transform 1 0 29808 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_324
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 1688980957
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 1688980957
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1688980957
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_461
timestamp 1688980957
transform 1 0 43516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_52
timestamp 1688980957
transform 1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_174
timestamp 1688980957
transform 1 0 17112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_208
timestamp 1688980957
transform 1 0 20240 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_241
timestamp 1688980957
transform 1 0 23276 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_262
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_269
timestamp 1688980957
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 1688980957
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 1688980957
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1688980957
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1688980957
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_457
timestamp 1688980957
transform 1 0 43148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_461
timestamp 1688980957
transform 1 0 43516 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_141
timestamp 1688980957
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_174
timestamp 1688980957
transform 1 0 17112 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_194
timestamp 1688980957
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_201
timestamp 1688980957
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_209
timestamp 1688980957
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_213
timestamp 1688980957
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_220
timestamp 1688980957
transform 1 0 21344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_238
timestamp 1688980957
transform 1 0 23000 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_247
timestamp 1688980957
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_251
timestamp 1688980957
transform 1 0 24196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_255
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_265
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_300
timestamp 1688980957
transform 1 0 28704 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_312
timestamp 1688980957
transform 1 0 29808 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_324
timestamp 1688980957
transform 1 0 30912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 1688980957
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_429
timestamp 1688980957
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 1688980957
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_461
timestamp 1688980957
transform 1 0 43516 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_19
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_113
timestamp 1688980957
transform 1 0 11500 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_118
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_150
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_185
timestamp 1688980957
transform 1 0 18124 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_190
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1688980957
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_203
timestamp 1688980957
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_232
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_267
timestamp 1688980957
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_281
timestamp 1688980957
transform 1 0 26956 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_303
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_326
timestamp 1688980957
transform 1 0 31096 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_338
timestamp 1688980957
transform 1 0 32200 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_350
timestamp 1688980957
transform 1 0 33304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_362
timestamp 1688980957
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 1688980957
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 1688980957
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_457
timestamp 1688980957
transform 1 0 43148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_461
timestamp 1688980957
transform 1 0 43516 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_83
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_92
timestamp 1688980957
transform 1 0 9568 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_96
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_99
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_103
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_117
timestamp 1688980957
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_157
timestamp 1688980957
transform 1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_200
timestamp 1688980957
transform 1 0 19504 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_243
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_251
timestamp 1688980957
transform 1 0 24196 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_259
timestamp 1688980957
transform 1 0 24932 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_271
timestamp 1688980957
transform 1 0 26036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1688980957
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_287
timestamp 1688980957
transform 1 0 27508 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_300
timestamp 1688980957
transform 1 0 28704 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_312
timestamp 1688980957
transform 1 0 29808 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_324
timestamp 1688980957
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1688980957
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 1688980957
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 1688980957
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 1688980957
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_461
timestamp 1688980957
transform 1 0 43516 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_80
timestamp 1688980957
transform 1 0 8464 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_110
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_126
timestamp 1688980957
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_169
timestamp 1688980957
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_178
timestamp 1688980957
transform 1 0 17480 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_204
timestamp 1688980957
transform 1 0 19872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_211
timestamp 1688980957
transform 1 0 20516 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_223
timestamp 1688980957
transform 1 0 21620 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_227
timestamp 1688980957
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_231
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_247
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 1688980957
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1688980957
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 1688980957
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 1688980957
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_457
timestamp 1688980957
transform 1 0 43148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_461
timestamp 1688980957
transform 1 0 43516 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_35
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_45
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_79
timestamp 1688980957
transform 1 0 8372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 1688980957
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_128
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_159
timestamp 1688980957
transform 1 0 15732 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_163
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_178
timestamp 1688980957
transform 1 0 17480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_212
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_220
timestamp 1688980957
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_231
timestamp 1688980957
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_252
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_260
timestamp 1688980957
transform 1 0 25024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_264
timestamp 1688980957
transform 1 0 25392 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_271
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_307
timestamp 1688980957
transform 1 0 29348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_319
timestamp 1688980957
transform 1 0 30452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_331
timestamp 1688980957
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_417
timestamp 1688980957
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_429
timestamp 1688980957
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_441
timestamp 1688980957
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 1688980957
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_461
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_58
timestamp 1688980957
transform 1 0 6440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_62
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_71
timestamp 1688980957
transform 1 0 7636 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_76
timestamp 1688980957
transform 1 0 8096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_80
timestamp 1688980957
transform 1 0 8464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_151
timestamp 1688980957
transform 1 0 14996 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_160
timestamp 1688980957
transform 1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_169
timestamp 1688980957
transform 1 0 16652 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_257
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_264
timestamp 1688980957
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_283
timestamp 1688980957
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_287
timestamp 1688980957
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_304
timestamp 1688980957
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_344
timestamp 1688980957
transform 1 0 32752 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_348
timestamp 1688980957
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_360
timestamp 1688980957
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1688980957
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 1688980957
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 1688980957
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1688980957
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 1688980957
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 1688980957
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_457
timestamp 1688980957
transform 1 0 43148 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_461
timestamp 1688980957
transform 1 0 43516 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_34
timestamp 1688980957
transform 1 0 4232 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_44
timestamp 1688980957
transform 1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_52
timestamp 1688980957
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_62
timestamp 1688980957
transform 1 0 6808 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_66
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_70
timestamp 1688980957
transform 1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_75
timestamp 1688980957
transform 1 0 8004 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_79
timestamp 1688980957
transform 1 0 8372 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_88
timestamp 1688980957
transform 1 0 9200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_95
timestamp 1688980957
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_99
timestamp 1688980957
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_118
timestamp 1688980957
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_122
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_126
timestamp 1688980957
transform 1 0 12696 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_141
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_144
timestamp 1688980957
transform 1 0 14352 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_234
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_238
timestamp 1688980957
transform 1 0 23000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_253
timestamp 1688980957
transform 1 0 24380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_274
timestamp 1688980957
transform 1 0 26312 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_295
timestamp 1688980957
transform 1 0 28244 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_299
timestamp 1688980957
transform 1 0 28612 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_327
timestamp 1688980957
transform 1 0 31188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_334
timestamp 1688980957
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1688980957
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 1688980957
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_461
timestamp 1688980957
transform 1 0 43516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_51
timestamp 1688980957
transform 1 0 5796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_61
timestamp 1688980957
transform 1 0 6716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_72
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_101
timestamp 1688980957
transform 1 0 10396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_118
timestamp 1688980957
transform 1 0 11960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_123
timestamp 1688980957
transform 1 0 12420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_151
timestamp 1688980957
transform 1 0 14996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_232
timestamp 1688980957
transform 1 0 22448 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_240
timestamp 1688980957
transform 1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_261
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_281
timestamp 1688980957
transform 1 0 26956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 1688980957
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_313
timestamp 1688980957
transform 1 0 29900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_356
timestamp 1688980957
transform 1 0 33856 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 1688980957
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 1688980957
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1688980957
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_461
timestamp 1688980957
transform 1 0 43516 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_47
timestamp 1688980957
transform 1 0 5428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_76
timestamp 1688980957
transform 1 0 8096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_95
timestamp 1688980957
transform 1 0 9844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_121
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_142
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_213
timestamp 1688980957
transform 1 0 20700 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_230
timestamp 1688980957
transform 1 0 22264 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_285
timestamp 1688980957
transform 1 0 27324 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_356
timestamp 1688980957
transform 1 0 33856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_360
timestamp 1688980957
transform 1 0 34224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_364
timestamp 1688980957
transform 1 0 34592 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_376
timestamp 1688980957
transform 1 0 35696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_388
timestamp 1688980957
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1688980957
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 1688980957
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 1688980957
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 1688980957
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_24
timestamp 1688980957
transform 1 0 3312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_37
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_72
timestamp 1688980957
transform 1 0 7728 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_92
timestamp 1688980957
transform 1 0 9568 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_116
timestamp 1688980957
transform 1 0 11776 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_120
timestamp 1688980957
transform 1 0 12144 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_163
timestamp 1688980957
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_173
timestamp 1688980957
transform 1 0 17020 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_191
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_203
timestamp 1688980957
transform 1 0 19780 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_214
timestamp 1688980957
transform 1 0 20792 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_220
timestamp 1688980957
transform 1 0 21344 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_225
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_263
timestamp 1688980957
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_275
timestamp 1688980957
transform 1 0 26404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_312
timestamp 1688980957
transform 1 0 29808 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_344
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_348
timestamp 1688980957
transform 1 0 33120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_353
timestamp 1688980957
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_361
timestamp 1688980957
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_461
timestamp 1688980957
transform 1 0 43516 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_25
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_50
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_68
timestamp 1688980957
transform 1 0 7360 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_72
timestamp 1688980957
transform 1 0 7728 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_76
timestamp 1688980957
transform 1 0 8096 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_80
timestamp 1688980957
transform 1 0 8464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_88
timestamp 1688980957
transform 1 0 9200 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_92
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_96
timestamp 1688980957
transform 1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_101
timestamp 1688980957
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_117
timestamp 1688980957
transform 1 0 11868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_121
timestamp 1688980957
transform 1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_129
timestamp 1688980957
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_140
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_144
timestamp 1688980957
transform 1 0 14352 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_151
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_165
timestamp 1688980957
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_172
timestamp 1688980957
transform 1 0 16928 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_176
timestamp 1688980957
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_185
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_197
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_220
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_256
timestamp 1688980957
transform 1 0 24656 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_260
timestamp 1688980957
transform 1 0 25024 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_264
timestamp 1688980957
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_268
timestamp 1688980957
transform 1 0 25760 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_276
timestamp 1688980957
transform 1 0 26496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_292
timestamp 1688980957
transform 1 0 27968 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_325
timestamp 1688980957
transform 1 0 31004 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_353
timestamp 1688980957
transform 1 0 33580 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_365
timestamp 1688980957
transform 1 0 34684 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_377
timestamp 1688980957
transform 1 0 35788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 1688980957
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_19
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_24
timestamp 1688980957
transform 1 0 3312 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_34
timestamp 1688980957
transform 1 0 4232 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_38
timestamp 1688980957
transform 1 0 4600 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_60
timestamp 1688980957
transform 1 0 6624 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_64
timestamp 1688980957
transform 1 0 6992 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_75
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_79
timestamp 1688980957
transform 1 0 8372 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_91
timestamp 1688980957
transform 1 0 9476 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_99
timestamp 1688980957
transform 1 0 10212 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_104
timestamp 1688980957
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_108
timestamp 1688980957
transform 1 0 11040 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_111
timestamp 1688980957
transform 1 0 11316 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_115
timestamp 1688980957
transform 1 0 11684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_127
timestamp 1688980957
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_131
timestamp 1688980957
transform 1 0 13156 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_167
timestamp 1688980957
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_171
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_184
timestamp 1688980957
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_228
timestamp 1688980957
transform 1 0 22080 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_232
timestamp 1688980957
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_240
timestamp 1688980957
transform 1 0 23184 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_262
timestamp 1688980957
transform 1 0 25208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_271
timestamp 1688980957
transform 1 0 26036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_331
timestamp 1688980957
transform 1 0 31556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_349
timestamp 1688980957
transform 1 0 33212 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_353
timestamp 1688980957
transform 1 0 33580 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_461
timestamp 1688980957
transform 1 0 43516 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_19
timestamp 1688980957
transform 1 0 2852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_35
timestamp 1688980957
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_47
timestamp 1688980957
transform 1 0 5428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_66
timestamp 1688980957
transform 1 0 7176 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_76
timestamp 1688980957
transform 1 0 8096 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_95
timestamp 1688980957
transform 1 0 9844 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_101
timestamp 1688980957
transform 1 0 10396 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_123
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_127
timestamp 1688980957
transform 1 0 12788 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_135
timestamp 1688980957
transform 1 0 13524 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_152
timestamp 1688980957
transform 1 0 15088 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_173
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_232
timestamp 1688980957
transform 1 0 22448 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_265
timestamp 1688980957
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_270
timestamp 1688980957
transform 1 0 25944 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_274
timestamp 1688980957
transform 1 0 26312 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_294
timestamp 1688980957
transform 1 0 28152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_298
timestamp 1688980957
transform 1 0 28520 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_302
timestamp 1688980957
transform 1 0 28888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_308
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_358
timestamp 1688980957
transform 1 0 34040 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_362
timestamp 1688980957
transform 1 0 34408 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_374
timestamp 1688980957
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_386
timestamp 1688980957
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_19
timestamp 1688980957
transform 1 0 2852 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_51
timestamp 1688980957
transform 1 0 5796 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_55
timestamp 1688980957
transform 1 0 6164 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_59
timestamp 1688980957
transform 1 0 6532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_80
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_92
timestamp 1688980957
transform 1 0 9568 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_148
timestamp 1688980957
transform 1 0 14720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_170
timestamp 1688980957
transform 1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_191
timestamp 1688980957
transform 1 0 18676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_259
timestamp 1688980957
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_273
timestamp 1688980957
transform 1 0 26220 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_295
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_299
timestamp 1688980957
transform 1 0 28612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_319
timestamp 1688980957
transform 1 0 30452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_356
timestamp 1688980957
transform 1 0 33856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_360
timestamp 1688980957
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 1688980957
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 1688980957
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 1688980957
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_457
timestamp 1688980957
transform 1 0 43148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_461
timestamp 1688980957
transform 1 0 43516 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_29
timestamp 1688980957
transform 1 0 3772 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_37
timestamp 1688980957
transform 1 0 4508 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_62
timestamp 1688980957
transform 1 0 6808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_66
timestamp 1688980957
transform 1 0 7176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_73
timestamp 1688980957
transform 1 0 7820 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_85
timestamp 1688980957
transform 1 0 8924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1688980957
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_116
timestamp 1688980957
transform 1 0 11776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_139
timestamp 1688980957
transform 1 0 13892 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_143
timestamp 1688980957
transform 1 0 14260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_153
timestamp 1688980957
transform 1 0 15180 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 1688980957
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_218
timestamp 1688980957
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_253
timestamp 1688980957
transform 1 0 24380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_257
timestamp 1688980957
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_269
timestamp 1688980957
transform 1 0 25852 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_276
timestamp 1688980957
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_294
timestamp 1688980957
transform 1 0 28152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_325
timestamp 1688980957
transform 1 0 31004 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_358
timestamp 1688980957
transform 1 0 34040 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_370
timestamp 1688980957
transform 1 0 35144 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_382
timestamp 1688980957
transform 1 0 36248 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_390
timestamp 1688980957
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 1688980957
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 1688980957
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 1688980957
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 1688980957
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_449
timestamp 1688980957
transform 1 0 42412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_25
timestamp 1688980957
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_34
timestamp 1688980957
transform 1 0 4232 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_38
timestamp 1688980957
transform 1 0 4600 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_49
timestamp 1688980957
transform 1 0 5612 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_57
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_68
timestamp 1688980957
transform 1 0 7360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_72
timestamp 1688980957
transform 1 0 7728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_82
timestamp 1688980957
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_91
timestamp 1688980957
transform 1 0 9476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_105
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_120
timestamp 1688980957
transform 1 0 12144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_124
timestamp 1688980957
transform 1 0 12512 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_146
timestamp 1688980957
transform 1 0 14536 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_150
timestamp 1688980957
transform 1 0 14904 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_154
timestamp 1688980957
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_158
timestamp 1688980957
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_178
timestamp 1688980957
transform 1 0 17480 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_235
timestamp 1688980957
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1688980957
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_261
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_269
timestamp 1688980957
transform 1 0 25852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_278
timestamp 1688980957
transform 1 0 26680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_291
timestamp 1688980957
transform 1 0 27876 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_298
timestamp 1688980957
transform 1 0 28520 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_315
timestamp 1688980957
transform 1 0 30084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 1688980957
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 1688980957
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 1688980957
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_433
timestamp 1688980957
transform 1 0 40940 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_441
timestamp 1688980957
transform 1 0 41676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_460
timestamp 1688980957
transform 1 0 43424 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_35
timestamp 1688980957
transform 1 0 4324 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_46
timestamp 1688980957
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1688980957
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_61
timestamp 1688980957
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_77
timestamp 1688980957
transform 1 0 8188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_95
timestamp 1688980957
transform 1 0 9844 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_103
timestamp 1688980957
transform 1 0 10580 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_140
timestamp 1688980957
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_146
timestamp 1688980957
transform 1 0 14536 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_183
timestamp 1688980957
transform 1 0 17940 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_197
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_222
timestamp 1688980957
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_241
timestamp 1688980957
transform 1 0 23276 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_268
timestamp 1688980957
transform 1 0 25760 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_272
timestamp 1688980957
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_297
timestamp 1688980957
transform 1 0 28428 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_314
timestamp 1688980957
transform 1 0 29992 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_320
timestamp 1688980957
transform 1 0 30544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_357
timestamp 1688980957
transform 1 0 33948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_365
timestamp 1688980957
transform 1 0 34684 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_377
timestamp 1688980957
transform 1 0 35788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_389
timestamp 1688980957
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 1688980957
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 1688980957
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 1688980957
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 1688980957
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 1688980957
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_461
timestamp 1688980957
transform 1 0 43516 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_19
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_38
timestamp 1688980957
transform 1 0 4600 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_52
timestamp 1688980957
transform 1 0 5888 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_73
timestamp 1688980957
transform 1 0 7820 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_92
timestamp 1688980957
transform 1 0 9568 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_102
timestamp 1688980957
transform 1 0 10488 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_164
timestamp 1688980957
transform 1 0 16192 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_175
timestamp 1688980957
transform 1 0 17204 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_249
timestamp 1688980957
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_259
timestamp 1688980957
transform 1 0 24932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_263
timestamp 1688980957
transform 1 0 25300 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_267
timestamp 1688980957
transform 1 0 25668 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_278
timestamp 1688980957
transform 1 0 26680 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_293
timestamp 1688980957
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_332
timestamp 1688980957
transform 1 0 31648 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_341
timestamp 1688980957
transform 1 0 32476 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_384
timestamp 1688980957
transform 1 0 36432 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_396
timestamp 1688980957
transform 1 0 37536 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_408
timestamp 1688980957
transform 1 0 38640 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1688980957
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 1688980957
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_457
timestamp 1688980957
transform 1 0 43148 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_461
timestamp 1688980957
transform 1 0 43516 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_52
timestamp 1688980957
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_67
timestamp 1688980957
transform 1 0 7268 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_74
timestamp 1688980957
transform 1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_91
timestamp 1688980957
transform 1 0 9476 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_97
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_107
timestamp 1688980957
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_118
timestamp 1688980957
transform 1 0 11960 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_123
timestamp 1688980957
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_130
timestamp 1688980957
transform 1 0 13064 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_164
timestamp 1688980957
transform 1 0 16192 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_194
timestamp 1688980957
transform 1 0 18952 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_201
timestamp 1688980957
transform 1 0 19596 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_233
timestamp 1688980957
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_252
timestamp 1688980957
transform 1 0 24288 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_260
timestamp 1688980957
transform 1 0 25024 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_286
timestamp 1688980957
transform 1 0 27416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_296
timestamp 1688980957
transform 1 0 28336 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_300
timestamp 1688980957
transform 1 0 28704 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_353
timestamp 1688980957
transform 1 0 33580 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_365
timestamp 1688980957
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_377
timestamp 1688980957
transform 1 0 35788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_389
timestamp 1688980957
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 1688980957
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 1688980957
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 1688980957
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 1688980957
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 1688980957
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_461
timestamp 1688980957
transform 1 0 43516 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_33
timestamp 1688980957
transform 1 0 4140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_57
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_64
timestamp 1688980957
transform 1 0 6992 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_75
timestamp 1688980957
transform 1 0 8004 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_80
timestamp 1688980957
transform 1 0 8464 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_102
timestamp 1688980957
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_106
timestamp 1688980957
transform 1 0 10856 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_131
timestamp 1688980957
transform 1 0 13156 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_136
timestamp 1688980957
transform 1 0 13616 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_150
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_163
timestamp 1688980957
transform 1 0 16100 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1688980957
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_206
timestamp 1688980957
transform 1 0 20056 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_213
timestamp 1688980957
transform 1 0 20700 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_244
timestamp 1688980957
transform 1 0 23552 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_248
timestamp 1688980957
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_267
timestamp 1688980957
transform 1 0 25668 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_275
timestamp 1688980957
transform 1 0 26404 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_283
timestamp 1688980957
transform 1 0 27140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_298
timestamp 1688980957
transform 1 0 28520 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_306
timestamp 1688980957
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_313
timestamp 1688980957
transform 1 0 29900 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_322
timestamp 1688980957
transform 1 0 30728 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_347
timestamp 1688980957
transform 1 0 33028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_359
timestamp 1688980957
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 1688980957
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 1688980957
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1688980957
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1688980957
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1688980957
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_457
timestamp 1688980957
transform 1 0 43148 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_461
timestamp 1688980957
transform 1 0 43516 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_26
timestamp 1688980957
transform 1 0 3496 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_37
timestamp 1688980957
transform 1 0 4508 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_46
timestamp 1688980957
transform 1 0 5336 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_50
timestamp 1688980957
transform 1 0 5704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_70
timestamp 1688980957
transform 1 0 7544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_90
timestamp 1688980957
transform 1 0 9384 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_130
timestamp 1688980957
transform 1 0 13064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_148
timestamp 1688980957
transform 1 0 14720 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_174
timestamp 1688980957
transform 1 0 17112 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_184
timestamp 1688980957
transform 1 0 18032 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_201
timestamp 1688980957
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_208
timestamp 1688980957
transform 1 0 20240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_214
timestamp 1688980957
transform 1 0 20792 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_246
timestamp 1688980957
transform 1 0 23736 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_287
timestamp 1688980957
transform 1 0 27508 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_302
timestamp 1688980957
transform 1 0 28888 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_306
timestamp 1688980957
transform 1 0 29256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_326
timestamp 1688980957
transform 1 0 31096 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_330
timestamp 1688980957
transform 1 0 31464 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_334
timestamp 1688980957
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1688980957
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 1688980957
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 1688980957
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 1688980957
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 1688980957
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_461
timestamp 1688980957
transform 1 0 43516 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_23
timestamp 1688980957
transform 1 0 3220 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_38
timestamp 1688980957
transform 1 0 4600 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_49
timestamp 1688980957
transform 1 0 5612 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_60
timestamp 1688980957
transform 1 0 6624 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_69
timestamp 1688980957
transform 1 0 7452 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_73
timestamp 1688980957
transform 1 0 7820 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_79
timestamp 1688980957
transform 1 0 8372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_102
timestamp 1688980957
transform 1 0 10488 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_111
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_115
timestamp 1688980957
transform 1 0 11684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_122
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_128
timestamp 1688980957
transform 1 0 12880 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_132
timestamp 1688980957
transform 1 0 13248 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_136
timestamp 1688980957
transform 1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_156
timestamp 1688980957
transform 1 0 15456 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_194
timestamp 1688980957
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_224
timestamp 1688980957
transform 1 0 21712 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_259
timestamp 1688980957
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_284
timestamp 1688980957
transform 1 0 27232 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_297
timestamp 1688980957
transform 1 0 28428 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 1688980957
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_313
timestamp 1688980957
transform 1 0 29900 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_348
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_360
timestamp 1688980957
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 1688980957
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 1688980957
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 1688980957
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1688980957
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1688980957
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1688980957
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_457
timestamp 1688980957
transform 1 0 43148 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_461
timestamp 1688980957
transform 1 0 43516 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_98
timestamp 1688980957
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_102
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_108
timestamp 1688980957
transform 1 0 11040 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_117
timestamp 1688980957
transform 1 0 11868 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_121
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_129
timestamp 1688980957
transform 1 0 12972 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_133
timestamp 1688980957
transform 1 0 13340 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_162
timestamp 1688980957
transform 1 0 16008 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_174
timestamp 1688980957
transform 1 0 17112 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_221
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_229
timestamp 1688980957
transform 1 0 22172 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_269
timestamp 1688980957
transform 1 0 25852 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_307
timestamp 1688980957
transform 1 0 29348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_318
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_340
timestamp 1688980957
transform 1 0 32384 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_344
timestamp 1688980957
transform 1 0 32752 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_356
timestamp 1688980957
transform 1 0 33856 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_368
timestamp 1688980957
transform 1 0 34960 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_380
timestamp 1688980957
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1688980957
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 1688980957
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 1688980957
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1688980957
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_461
timestamp 1688980957
transform 1 0 43516 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_6
timestamp 1688980957
transform 1 0 1656 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_24
timestamp 1688980957
transform 1 0 3312 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_33
timestamp 1688980957
transform 1 0 4140 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_55
timestamp 1688980957
transform 1 0 6164 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_73
timestamp 1688980957
transform 1 0 7820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_107
timestamp 1688980957
transform 1 0 10948 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_128
timestamp 1688980957
transform 1 0 12880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_174
timestamp 1688980957
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_239
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_268
timestamp 1688980957
transform 1 0 25760 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_283
timestamp 1688980957
transform 1 0 27140 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_295
timestamp 1688980957
transform 1 0 28244 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_299
timestamp 1688980957
transform 1 0 28612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_328
timestamp 1688980957
transform 1 0 31280 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_340
timestamp 1688980957
transform 1 0 32384 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_352
timestamp 1688980957
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1688980957
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1688980957
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 1688980957
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1688980957
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_457
timestamp 1688980957
transform 1 0 43148 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_461
timestamp 1688980957
transform 1 0 43516 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_7
timestamp 1688980957
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_35
timestamp 1688980957
transform 1 0 4324 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_65
timestamp 1688980957
transform 1 0 7084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_75
timestamp 1688980957
transform 1 0 8004 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_96
timestamp 1688980957
transform 1 0 9936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_100
timestamp 1688980957
transform 1 0 10304 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_135
timestamp 1688980957
transform 1 0 13524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_150
timestamp 1688980957
transform 1 0 14904 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_179
timestamp 1688980957
transform 1 0 17572 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_199
timestamp 1688980957
transform 1 0 19412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_252
timestamp 1688980957
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_267
timestamp 1688980957
transform 1 0 25668 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_274
timestamp 1688980957
transform 1 0 26312 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_278
timestamp 1688980957
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_285
timestamp 1688980957
transform 1 0 27324 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_289
timestamp 1688980957
transform 1 0 27692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_300
timestamp 1688980957
transform 1 0 28704 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_304
timestamp 1688980957
transform 1 0 29072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_322
timestamp 1688980957
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_334
timestamp 1688980957
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1688980957
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1688980957
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 1688980957
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 1688980957
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1688980957
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_461
timestamp 1688980957
transform 1 0 43516 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_6
timestamp 1688980957
transform 1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_26
timestamp 1688980957
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_52
timestamp 1688980957
transform 1 0 5888 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_80
timestamp 1688980957
transform 1 0 8464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_94
timestamp 1688980957
transform 1 0 9752 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_99
timestamp 1688980957
transform 1 0 10212 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_103
timestamp 1688980957
transform 1 0 10580 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_111
timestamp 1688980957
transform 1 0 11316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_126
timestamp 1688980957
transform 1 0 12696 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_137
timestamp 1688980957
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_172
timestamp 1688980957
transform 1 0 16928 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_232
timestamp 1688980957
transform 1 0 22448 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_322
timestamp 1688980957
transform 1 0 30728 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_326
timestamp 1688980957
transform 1 0 31096 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_330
timestamp 1688980957
transform 1 0 31464 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_342
timestamp 1688980957
transform 1 0 32568 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_354
timestamp 1688980957
transform 1 0 33672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_362
timestamp 1688980957
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1688980957
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1688980957
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_457
timestamp 1688980957
transform 1 0 43148 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_461
timestamp 1688980957
transform 1 0 43516 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_8
timestamp 1688980957
transform 1 0 1840 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_50
timestamp 1688980957
transform 1 0 5704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_73
timestamp 1688980957
transform 1 0 7820 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_100
timestamp 1688980957
transform 1 0 10304 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_104
timestamp 1688980957
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_108
timestamp 1688980957
transform 1 0 11040 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_158
timestamp 1688980957
transform 1 0 15640 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_187
timestamp 1688980957
transform 1 0 18308 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_204
timestamp 1688980957
transform 1 0 19872 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_245
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_255
timestamp 1688980957
transform 1 0 24564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_267
timestamp 1688980957
transform 1 0 25668 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_271
timestamp 1688980957
transform 1 0 26036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_303
timestamp 1688980957
transform 1 0 28980 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_331
timestamp 1688980957
transform 1 0 31556 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_341
timestamp 1688980957
transform 1 0 32476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_353
timestamp 1688980957
transform 1 0 33580 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_365
timestamp 1688980957
transform 1 0 34684 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_377
timestamp 1688980957
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_389
timestamp 1688980957
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 1688980957
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 1688980957
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_461
timestamp 1688980957
transform 1 0 43516 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_24
timestamp 1688980957
transform 1 0 3312 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_66
timestamp 1688980957
transform 1 0 7176 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_120
timestamp 1688980957
transform 1 0 12144 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_192
timestamp 1688980957
transform 1 0 18768 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_236
timestamp 1688980957
transform 1 0 22816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_242
timestamp 1688980957
transform 1 0 23368 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_246
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_256
timestamp 1688980957
transform 1 0 24656 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_260
timestamp 1688980957
transform 1 0 25024 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_274
timestamp 1688980957
transform 1 0 26312 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_295
timestamp 1688980957
transform 1 0 28244 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_306
timestamp 1688980957
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_319
timestamp 1688980957
transform 1 0 30452 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_339
timestamp 1688980957
transform 1 0 32292 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_343
timestamp 1688980957
transform 1 0 32660 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_347
timestamp 1688980957
transform 1 0 33028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_359
timestamp 1688980957
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1688980957
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1688980957
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1688980957
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_457
timestamp 1688980957
transform 1 0 43148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_461
timestamp 1688980957
transform 1 0 43516 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_97
timestamp 1688980957
transform 1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_103
timestamp 1688980957
transform 1 0 10580 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_134
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_164
timestamp 1688980957
transform 1 0 16192 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_250
timestamp 1688980957
transform 1 0 24104 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_275
timestamp 1688980957
transform 1 0 26404 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_316
timestamp 1688980957
transform 1 0 30176 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_345
timestamp 1688980957
transform 1 0 32844 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1688980957
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1688980957
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_93
timestamp 1688980957
transform 1 0 9660 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_108
timestamp 1688980957
transform 1 0 11040 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_117
timestamp 1688980957
transform 1 0 11868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_150
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_184
timestamp 1688980957
transform 1 0 18032 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_206
timestamp 1688980957
transform 1 0 20056 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_288
timestamp 1688980957
transform 1 0 27600 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_341
timestamp 1688980957
transform 1 0 32476 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_349
timestamp 1688980957
transform 1 0 33212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_361
timestamp 1688980957
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1688980957
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_457
timestamp 1688980957
transform 1 0 43148 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_461
timestamp 1688980957
transform 1 0 43516 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_23
timestamp 1688980957
transform 1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_49
timestamp 1688980957
transform 1 0 5612 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_53
timestamp 1688980957
transform 1 0 5980 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_87
timestamp 1688980957
transform 1 0 9108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_91
timestamp 1688980957
transform 1 0 9476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_122
timestamp 1688980957
transform 1 0 12328 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_152
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_238
timestamp 1688980957
transform 1 0 23000 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_258
timestamp 1688980957
transform 1 0 24840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_312
timestamp 1688980957
transform 1 0 29808 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_330
timestamp 1688980957
transform 1 0 31464 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_334
timestamp 1688980957
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_345
timestamp 1688980957
transform 1 0 32844 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_353
timestamp 1688980957
transform 1 0 33580 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_365
timestamp 1688980957
transform 1 0 34684 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_377
timestamp 1688980957
transform 1 0 35788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_389
timestamp 1688980957
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 1688980957
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 1688980957
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_461
timestamp 1688980957
transform 1 0 43516 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_19
timestamp 1688980957
transform 1 0 2852 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_23
timestamp 1688980957
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_49
timestamp 1688980957
transform 1 0 5612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_64
timestamp 1688980957
transform 1 0 6992 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_94
timestamp 1688980957
transform 1 0 9752 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_146
timestamp 1688980957
transform 1 0 14536 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_163
timestamp 1688980957
transform 1 0 16100 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_211
timestamp 1688980957
transform 1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_223
timestamp 1688980957
transform 1 0 21620 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_286
timestamp 1688980957
transform 1 0 27416 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 1688980957
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_318
timestamp 1688980957
transform 1 0 30360 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_334
timestamp 1688980957
transform 1 0 31832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_351
timestamp 1688980957
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_355
timestamp 1688980957
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1688980957
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 1688980957
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_457
timestamp 1688980957
transform 1 0 43148 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_461
timestamp 1688980957
transform 1 0 43516 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_67
timestamp 1688980957
transform 1 0 7268 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_96
timestamp 1688980957
transform 1 0 9936 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_110
timestamp 1688980957
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_122
timestamp 1688980957
transform 1 0 12328 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_142
timestamp 1688980957
transform 1 0 14168 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_206
timestamp 1688980957
transform 1 0 20056 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_213
timestamp 1688980957
transform 1 0 20700 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_221
timestamp 1688980957
transform 1 0 21436 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_229
timestamp 1688980957
transform 1 0 22172 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_248
timestamp 1688980957
transform 1 0 23920 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_285
timestamp 1688980957
transform 1 0 27324 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_332
timestamp 1688980957
transform 1 0 31648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_345
timestamp 1688980957
transform 1 0 32844 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_358
timestamp 1688980957
transform 1 0 34040 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_362
timestamp 1688980957
transform 1 0 34408 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_374
timestamp 1688980957
transform 1 0 35512 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_386
timestamp 1688980957
transform 1 0 36616 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 1688980957
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 1688980957
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_461
timestamp 1688980957
transform 1 0 43516 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_19
timestamp 1688980957
transform 1 0 2852 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_23
timestamp 1688980957
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_80
timestamp 1688980957
transform 1 0 8464 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_111
timestamp 1688980957
transform 1 0 11316 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_137
timestamp 1688980957
transform 1 0 13708 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_210
timestamp 1688980957
transform 1 0 20424 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_250
timestamp 1688980957
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_304
timestamp 1688980957
transform 1 0 29072 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_328
timestamp 1688980957
transform 1 0 31280 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_355
timestamp 1688980957
transform 1 0 33764 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 1688980957
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_457
timestamp 1688980957
transform 1 0 43148 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_461
timestamp 1688980957
transform 1 0 43516 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_47
timestamp 1688980957
transform 1 0 5428 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_66
timestamp 1688980957
transform 1 0 7176 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_144
timestamp 1688980957
transform 1 0 14352 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_163
timestamp 1688980957
transform 1 0 16100 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_202
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_206
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_209
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_213
timestamp 1688980957
transform 1 0 20700 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_220
timestamp 1688980957
transform 1 0 21344 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_259
timestamp 1688980957
transform 1 0 24932 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_277
timestamp 1688980957
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_322
timestamp 1688980957
transform 1 0 30728 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_345
timestamp 1688980957
transform 1 0 32844 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 1688980957
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 1688980957
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_461
timestamp 1688980957
transform 1 0 43516 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_19
timestamp 1688980957
transform 1 0 2852 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_23
timestamp 1688980957
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_49
timestamp 1688980957
transform 1 0 5612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_94
timestamp 1688980957
transform 1 0 9752 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_111
timestamp 1688980957
transform 1 0 11316 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_136
timestamp 1688980957
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_163
timestamp 1688980957
transform 1 0 16100 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_192
timestamp 1688980957
transform 1 0 18768 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_217
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_222
timestamp 1688980957
transform 1 0 21528 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_230
timestamp 1688980957
transform 1 0 22264 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_250
timestamp 1688980957
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_266
timestamp 1688980957
transform 1 0 25576 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_270
timestamp 1688980957
transform 1 0 25944 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_303
timestamp 1688980957
transform 1 0 28980 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_341
timestamp 1688980957
transform 1 0 32476 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1688980957
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1688980957
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1688980957
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 1688980957
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_457
timestamp 1688980957
transform 1 0 43148 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_74
timestamp 1688980957
transform 1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_86
timestamp 1688980957
transform 1 0 9016 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_97
timestamp 1688980957
transform 1 0 10028 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_110
timestamp 1688980957
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_119
timestamp 1688980957
transform 1 0 12052 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_179
timestamp 1688980957
transform 1 0 17572 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_188
timestamp 1688980957
transform 1 0 18400 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_200
timestamp 1688980957
transform 1 0 19504 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_212
timestamp 1688980957
transform 1 0 20608 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_231
timestamp 1688980957
transform 1 0 22356 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_234
timestamp 1688980957
transform 1 0 22632 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_238
timestamp 1688980957
transform 1 0 23000 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_267
timestamp 1688980957
transform 1 0 25668 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_271
timestamp 1688980957
transform 1 0 26036 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_275
timestamp 1688980957
transform 1 0 26404 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_281
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_285
timestamp 1688980957
transform 1 0 27324 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_333
timestamp 1688980957
transform 1 0 31740 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_341
timestamp 1688980957
transform 1 0 32476 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_345
timestamp 1688980957
transform 1 0 32844 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_357
timestamp 1688980957
transform 1 0 33948 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_369
timestamp 1688980957
transform 1 0 35052 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_381
timestamp 1688980957
transform 1 0 36156 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_389
timestamp 1688980957
transform 1 0 36892 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 1688980957
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 1688980957
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_461
timestamp 1688980957
transform 1 0 43516 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_6
timestamp 1688980957
transform 1 0 1656 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_18
timestamp 1688980957
transform 1 0 2760 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_26
timestamp 1688980957
transform 1 0 3496 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_73
timestamp 1688980957
transform 1 0 7820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_99
timestamp 1688980957
transform 1 0 10212 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_108
timestamp 1688980957
transform 1 0 11040 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_134
timestamp 1688980957
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_149
timestamp 1688980957
transform 1 0 14812 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_168
timestamp 1688980957
transform 1 0 16560 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_180
timestamp 1688980957
transform 1 0 17664 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_192
timestamp 1688980957
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1688980957
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1688980957
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_245
timestamp 1688980957
transform 1 0 23644 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_249
timestamp 1688980957
transform 1 0 24012 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_258
timestamp 1688980957
transform 1 0 24840 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_262
timestamp 1688980957
transform 1 0 25208 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_266
timestamp 1688980957
transform 1 0 25576 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_274
timestamp 1688980957
transform 1 0 26312 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_289
timestamp 1688980957
transform 1 0 27692 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_293
timestamp 1688980957
transform 1 0 28060 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_302
timestamp 1688980957
transform 1 0 28888 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1688980957
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1688980957
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1688980957
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_457
timestamp 1688980957
transform 1 0 43148 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_461
timestamp 1688980957
transform 1 0 43516 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_83
timestamp 1688980957
transform 1 0 8740 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_95
timestamp 1688980957
transform 1 0 9844 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_119
timestamp 1688980957
transform 1 0 12052 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_136
timestamp 1688980957
transform 1 0 13616 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_148
timestamp 1688980957
transform 1 0 14720 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_160
timestamp 1688980957
transform 1 0 15824 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1688980957
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1688980957
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1688980957
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1688980957
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1688980957
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_314
timestamp 1688980957
transform 1 0 29992 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_318
timestamp 1688980957
transform 1 0 30360 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_330
timestamp 1688980957
transform 1 0 31464 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1688980957
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1688980957
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1688980957
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1688980957
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_461
timestamp 1688980957
transform 1 0 43516 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_6
timestamp 1688980957
transform 1 0 1656 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_18
timestamp 1688980957
transform 1 0 2760 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_26
timestamp 1688980957
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1688980957
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1688980957
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1688980957
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1688980957
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1688980957
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_301
timestamp 1688980957
transform 1 0 28796 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_304
timestamp 1688980957
transform 1 0 29072 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1688980957
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1688980957
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1688980957
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1688980957
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_457
timestamp 1688980957
transform 1 0 43148 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_461
timestamp 1688980957
transform 1 0 43516 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_29
timestamp 1688980957
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_41
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_53
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_85
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_97
timestamp 1688980957
transform 1 0 10028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_109
timestamp 1688980957
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_141
timestamp 1688980957
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_153
timestamp 1688980957
transform 1 0 15180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_165
timestamp 1688980957
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_197
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_209
timestamp 1688980957
transform 1 0 20332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_221
timestamp 1688980957
transform 1 0 21436 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_256
timestamp 1688980957
transform 1 0 24656 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_264
timestamp 1688980957
transform 1 0 25392 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_268
timestamp 1688980957
transform 1 0 25760 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_284
timestamp 1688980957
transform 1 0 27232 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_290
timestamp 1688980957
transform 1 0 27784 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_294
timestamp 1688980957
transform 1 0 28152 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_302
timestamp 1688980957
transform 1 0 28888 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_307
timestamp 1688980957
transform 1 0 29348 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_309
timestamp 1688980957
transform 1 0 29532 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_320
timestamp 1688980957
transform 1 0 30544 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_328
timestamp 1688980957
transform 1 0 31280 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_333
timestamp 1688980957
transform 1 0 31740 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_346
timestamp 1688980957
transform 1 0 32936 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_358
timestamp 1688980957
transform 1 0 34040 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_365
timestamp 1688980957
transform 1 0 34684 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_381
timestamp 1688980957
transform 1 0 36156 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 1688980957
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1688980957
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_398
timestamp 1688980957
transform 1 0 37720 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_410
timestamp 1688980957
transform 1 0 38824 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_418
timestamp 1688980957
transform 1 0 39560 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_421
timestamp 1688980957
transform 1 0 39836 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_433
timestamp 1688980957
transform 1 0 40940 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_445
timestamp 1688980957
transform 1 0 42044 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_461
timestamp 1688980957
transform 1 0 43516 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 26128 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 24104 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 23368 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 9108 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 6624 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 24104 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 22908 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 9752 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 3864 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 4324 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 10304 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 6624 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 5888 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 9292 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 12144 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 9016 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 6440 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 5888 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 3864 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 4048 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 32292 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 29992 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 12880 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 11868 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 5520 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 7176 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 15824 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 14352 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 18768 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 16836 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 12512 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 13248 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 3404 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 4784 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 16008 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 15088 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 8096 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 8004 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 13616 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 11408 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 10672 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 9936 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 11868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 15548 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 14260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 20700 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 22356 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 7360 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 18400 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 11500 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 18952 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 16836 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 17664 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 18032 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 17204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 16468 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 14444 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 14444 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 18400 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 19228 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 20148 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 19872 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 17296 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 18216 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 3496 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 1932 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 20516 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 8096 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 7268 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 2760 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 2024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold93 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 27508 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 26680 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold100
timestamp 1688980957
transform 1 0 13800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 30544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 31004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 5704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform 1 0 28888 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 4048 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold114
timestamp 1688980957
transform 1 0 18124 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 17204 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold118
timestamp 1688980957
transform 1 0 5612 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 23460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold122
timestamp 1688980957
transform 1 0 19044 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 20148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform 1 0 5060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 4232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 4232 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 25208 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 23828 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold135
timestamp 1688980957
transform 1 0 15824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold139
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform 1 0 6256 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 20792 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 30728 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 32292 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 15548 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold149 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28612 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 30544 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold151
timestamp 1688980957
transform 1 0 31096 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  hold152
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 29992 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform 1 0 32016 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 31280 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold156
timestamp 1688980957
transform 1 0 31556 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform 1 0 22356 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 18216 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold160
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 27048 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform 1 0 27508 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform 1 0 32476 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold166
timestamp 1688980957
transform 1 0 31004 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform 1 0 20056 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold169
timestamp 1688980957
transform 1 0 20148 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold171
timestamp 1688980957
transform 1 0 8096 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 6716 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold173 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform 1 0 23000 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold175
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform 1 0 14904 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold177
timestamp 1688980957
transform 1 0 12052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform 1 0 4968 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold180
timestamp 1688980957
transform 1 0 6072 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform 1 0 4876 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold185
timestamp 1688980957
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold188
timestamp 1688980957
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold191 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 2852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold193
timestamp 1688980957
transform 1 0 3680 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold194
timestamp 1688980957
transform 1 0 9200 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform 1 0 6532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold198
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 17848 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform 1 0 10580 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 22264 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 30636 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform 1 0 3496 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 1840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold213
timestamp 1688980957
transform 1 0 31096 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 33028 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold217
timestamp 1688980957
transform 1 0 33304 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 25392 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform 1 0 30820 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 29256 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform 1 0 28152 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold225
timestamp 1688980957
transform 1 0 22448 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform 1 0 2944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 28244 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold229
timestamp 1688980957
transform 1 0 26496 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform 1 0 2208 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform 1 0 16376 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 15640 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform 1 0 14352 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform 1 0 27968 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform 1 0 26956 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 25392 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform 1 0 29624 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 31464 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform 1 0 24196 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 43332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 43332 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 25484 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 27876 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 29072 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 30268 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 31464 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 32660 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 35052 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 36248 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 37444 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1688980957
transform 1 0 43056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap47
timestamp 1688980957
transform 1 0 13248 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  output15 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output16
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output17
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output18
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output19
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output20
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output35
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output36
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output37
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 43884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 43884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 43884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 43884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 43884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 43884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 43884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 43884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 43884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 43884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 43884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 43884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 43884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 43884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 43884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 43884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 43884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 43884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 43884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 43884 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 43884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 43884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 43884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 43884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 43884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 43884 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 43884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 43884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 43884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 43884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 43884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 43884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 43884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 43884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 43884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 43884 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 43884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 43884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 43884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 43884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 43884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 43884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 43884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 43884 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 43884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 43884 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 43884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 43884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 43884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 43884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 43884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 43884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 43884 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 43884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 43884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 43884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 43884 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 43884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 43884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 43884 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 34592 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire51
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_80 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_81
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_82
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_83
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapped_6502_84
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 314 592
<< labels >>
flabel metal3 s 44200 28024 45000 28144 0 FreeSans 480 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 44200 39176 45000 39296 0 FreeSans 480 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal2 s 1490 44200 1546 45000 0 FreeSans 224 90 0 0 io_in[0]
port 2 nsew signal input
flabel metal2 s 13450 44200 13506 45000 0 FreeSans 224 90 0 0 io_in[10]
port 3 nsew signal input
flabel metal2 s 14646 44200 14702 45000 0 FreeSans 224 90 0 0 io_in[11]
port 4 nsew signal input
flabel metal2 s 15842 44200 15898 45000 0 FreeSans 224 90 0 0 io_in[12]
port 5 nsew signal input
flabel metal2 s 17038 44200 17094 45000 0 FreeSans 224 90 0 0 io_in[13]
port 6 nsew signal input
flabel metal2 s 18234 44200 18290 45000 0 FreeSans 224 90 0 0 io_in[14]
port 7 nsew signal input
flabel metal2 s 19430 44200 19486 45000 0 FreeSans 224 90 0 0 io_in[15]
port 8 nsew signal input
flabel metal2 s 20626 44200 20682 45000 0 FreeSans 224 90 0 0 io_in[16]
port 9 nsew signal input
flabel metal2 s 21822 44200 21878 45000 0 FreeSans 224 90 0 0 io_in[17]
port 10 nsew signal input
flabel metal2 s 23018 44200 23074 45000 0 FreeSans 224 90 0 0 io_in[18]
port 11 nsew signal input
flabel metal2 s 24214 44200 24270 45000 0 FreeSans 224 90 0 0 io_in[19]
port 12 nsew signal input
flabel metal2 s 2686 44200 2742 45000 0 FreeSans 224 90 0 0 io_in[1]
port 13 nsew signal input
flabel metal2 s 25410 44200 25466 45000 0 FreeSans 224 90 0 0 io_in[20]
port 14 nsew signal input
flabel metal2 s 26606 44200 26662 45000 0 FreeSans 224 90 0 0 io_in[21]
port 15 nsew signal input
flabel metal2 s 27802 44200 27858 45000 0 FreeSans 224 90 0 0 io_in[22]
port 16 nsew signal input
flabel metal2 s 28998 44200 29054 45000 0 FreeSans 224 90 0 0 io_in[23]
port 17 nsew signal input
flabel metal2 s 30194 44200 30250 45000 0 FreeSans 224 90 0 0 io_in[24]
port 18 nsew signal input
flabel metal2 s 31390 44200 31446 45000 0 FreeSans 224 90 0 0 io_in[25]
port 19 nsew signal input
flabel metal2 s 32586 44200 32642 45000 0 FreeSans 224 90 0 0 io_in[26]
port 20 nsew signal input
flabel metal2 s 33782 44200 33838 45000 0 FreeSans 224 90 0 0 io_in[27]
port 21 nsew signal input
flabel metal2 s 34978 44200 35034 45000 0 FreeSans 224 90 0 0 io_in[28]
port 22 nsew signal input
flabel metal2 s 36174 44200 36230 45000 0 FreeSans 224 90 0 0 io_in[29]
port 23 nsew signal input
flabel metal2 s 3882 44200 3938 45000 0 FreeSans 224 90 0 0 io_in[2]
port 24 nsew signal input
flabel metal2 s 37370 44200 37426 45000 0 FreeSans 224 90 0 0 io_in[30]
port 25 nsew signal input
flabel metal2 s 38566 44200 38622 45000 0 FreeSans 224 90 0 0 io_in[31]
port 26 nsew signal input
flabel metal2 s 39762 44200 39818 45000 0 FreeSans 224 90 0 0 io_in[32]
port 27 nsew signal input
flabel metal2 s 40958 44200 41014 45000 0 FreeSans 224 90 0 0 io_in[33]
port 28 nsew signal input
flabel metal2 s 42154 44200 42210 45000 0 FreeSans 224 90 0 0 io_in[34]
port 29 nsew signal input
flabel metal2 s 43350 44200 43406 45000 0 FreeSans 224 90 0 0 io_in[35]
port 30 nsew signal input
flabel metal2 s 5078 44200 5134 45000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 6274 44200 6330 45000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 7470 44200 7526 45000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 8666 44200 8722 45000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 9862 44200 9918 45000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 11058 44200 11114 45000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 12254 44200 12310 45000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 io_oeb
port 38 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 io_out[0]
port 39 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_out[10]
port 40 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_out[11]
port 41 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 io_out[12]
port 42 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 io_out[13]
port 43 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 io_out[14]
port 44 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 io_out[15]
port 45 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_out[16]
port 46 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 io_out[17]
port 47 nsew signal tristate
flabel metal3 s 0 22856 800 22976 0 FreeSans 480 0 0 0 io_out[18]
port 48 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 io_out[19]
port 49 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_out[1]
port 50 nsew signal tristate
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 io_out[20]
port 51 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[21]
port 52 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 io_out[22]
port 53 nsew signal tristate
flabel metal3 s 0 28296 800 28416 0 FreeSans 480 0 0 0 io_out[23]
port 54 nsew signal tristate
flabel metal3 s 0 29384 800 29504 0 FreeSans 480 0 0 0 io_out[24]
port 55 nsew signal tristate
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 io_out[25]
port 56 nsew signal tristate
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 io_out[26]
port 57 nsew signal tristate
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 io_out[27]
port 58 nsew signal tristate
flabel metal3 s 0 33736 800 33856 0 FreeSans 480 0 0 0 io_out[28]
port 59 nsew signal tristate
flabel metal3 s 0 34824 800 34944 0 FreeSans 480 0 0 0 io_out[29]
port 60 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 io_out[2]
port 61 nsew signal tristate
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 io_out[30]
port 62 nsew signal tristate
flabel metal3 s 0 37000 800 37120 0 FreeSans 480 0 0 0 io_out[31]
port 63 nsew signal tristate
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_out[32]
port 64 nsew signal tristate
flabel metal3 s 0 39176 800 39296 0 FreeSans 480 0 0 0 io_out[33]
port 65 nsew signal tristate
flabel metal3 s 0 40264 800 40384 0 FreeSans 480 0 0 0 io_out[34]
port 66 nsew signal tristate
flabel metal3 s 0 41352 800 41472 0 FreeSans 480 0 0 0 io_out[35]
port 67 nsew signal tristate
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 io_out[3]
port 68 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 io_out[4]
port 69 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 io_out[5]
port 70 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[6]
port 71 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 io_out[7]
port 72 nsew signal tristate
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 io_out[8]
port 73 nsew signal tristate
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 io_out[9]
port 74 nsew signal tristate
flabel metal3 s 44200 16872 45000 16992 0 FreeSans 480 0 0 0 rst_n
port 75 nsew signal input
flabel metal4 s 4208 2128 4528 42480 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 2128 35248 42480 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 19568 2128 19888 42480 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal3 s 44200 5720 45000 5840 0 FreeSans 480 0 0 0 wb_clk_i
port 78 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 45000 45000
<< end >>
