VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_fgcaptest
  CLASS BLOCK ;
  FOREIGN top_fgcaptest ;
  ORIGIN 48.000 174.000 ;
  SIZE 681.000 BY 630.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 273.000 434.000 275.000 456.000 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 279.000 437.000 281.000 456.000 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 285.000 440.000 287.000 456.000 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 291.000 443.000 293.000 456.000 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 297.000 446.000 299.000 456.000 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 303.000 444.200 305.000 456.000 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 309.000 441.200 311.000 456.000 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 315.000 438.200 317.000 456.000 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.415000 ;
    PORT
      LAYER met3 ;
        RECT 321.000 435.200 323.000 456.000 ;
    END
  END addr[8]
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 629.000 -174.000 633.000 437.000 ;
    END
  END vssd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT -48.000 -174.000 -44.000 456.000 ;
    END
  END vccd2
  OBS
      LAYER nwell ;
        RECT 0.000 -157.065 599.830 446.230 ;
      LAYER li1 ;
        RECT 0.020 -156.935 599.810 446.210 ;
      LAYER met1 ;
        RECT 0.010 -160.375 599.820 446.220 ;
      LAYER met2 ;
        RECT 0.000 -171.175 602.420 446.230 ;
      LAYER met3 ;
        RECT 0.580 433.600 272.600 450.000 ;
        RECT 275.400 436.600 278.600 450.000 ;
        RECT 281.400 439.600 284.600 450.000 ;
        RECT 287.400 442.600 290.600 450.000 ;
        RECT 293.400 445.600 296.600 450.000 ;
        RECT 299.400 445.600 302.600 450.000 ;
        RECT 293.400 443.800 302.600 445.600 ;
        RECT 305.400 443.800 308.600 450.000 ;
        RECT 293.400 442.600 308.600 443.800 ;
        RECT 287.400 440.800 308.600 442.600 ;
        RECT 311.400 440.800 314.600 450.000 ;
        RECT 287.400 439.600 314.600 440.800 ;
        RECT 281.400 437.800 314.600 439.600 ;
        RECT 317.400 437.800 320.600 450.000 ;
        RECT 281.400 436.600 320.600 437.800 ;
        RECT 275.400 434.800 320.600 436.600 ;
        RECT 323.400 434.800 602.420 450.000 ;
        RECT 275.400 433.600 602.420 434.800 ;
        RECT 0.580 -173.675 602.420 433.600 ;
      LAYER met4 ;
        RECT -43.600 437.400 629.000 456.000 ;
        RECT -43.600 -174.000 628.600 437.400 ;
      LAYER met5 ;
        RECT -5.000 -174.000 604.600 456.000 ;
  END
END top_fgcaptest
END LIBRARY

