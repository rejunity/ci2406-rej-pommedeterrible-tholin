* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for execution_unit abstract view
.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_idx[5]
+ dest_mask[0] dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0]
+ dest_val[10] dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16]
+ dest_val[17] dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22]
+ dest_val[23] dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29]
+ dest_val[2] dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6]
+ dest_val[7] dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11]
+ instruction[12] instruction[13] instruction[14] instruction[15] instruction[16]
+ instruction[17] instruction[18] instruction[19] instruction[1] instruction[20] instruction[21]
+ instruction[22] instruction[23] instruction[24] instruction[25] instruction[26]
+ instruction[27] instruction[28] instruction[29] instruction[2] instruction[30] instruction[31]
+ instruction[32] instruction[33] instruction[34] instruction[35] instruction[36]
+ instruction[37] instruction[38] instruction[39] instruction[3] instruction[40] instruction[41]
+ instruction[4] instruction[5] instruction[6] instruction[7] instruction[8] instruction[9]
+ int_return is_load is_store loadstore_address[0] loadstore_address[10] loadstore_address[11]
+ loadstore_address[12] loadstore_address[13] loadstore_address[14] loadstore_address[15]
+ loadstore_address[16] loadstore_address[17] loadstore_address[18] loadstore_address[19]
+ loadstore_address[1] loadstore_address[20] loadstore_address[21] loadstore_address[22]
+ loadstore_address[23] loadstore_address[24] loadstore_address[25] loadstore_address[26]
+ loadstore_address[27] loadstore_address[28] loadstore_address[29] loadstore_address[2]
+ loadstore_address[30] loadstore_address[31] loadstore_address[3] loadstore_address[4]
+ loadstore_address[5] loadstore_address[6] loadstore_address[7] loadstore_address[8]
+ loadstore_address[9] loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3]
+ loadstore_dest[4] loadstore_dest[5] loadstore_size[0] loadstore_size[1] new_PC[0]
+ new_PC[10] new_PC[11] new_PC[12] new_PC[13] new_PC[14] new_PC[15] new_PC[16] new_PC[17]
+ new_PC[18] new_PC[19] new_PC[1] new_PC[20] new_PC[21] new_PC[22] new_PC[23] new_PC[24]
+ new_PC[25] new_PC[26] new_PC[27] new_PC[2] new_PC[3] new_PC[4] new_PC[5] new_PC[6]
+ new_PC[7] new_PC[8] new_PC[9] pred_idx[0] pred_idx[1] pred_idx[2] pred_val reg1_idx[0]
+ reg1_idx[1] reg1_idx[2] reg1_idx[3] reg1_idx[4] reg1_idx[5] reg1_val[0] reg1_val[10]
+ reg1_val[11] reg1_val[12] reg1_val[13] reg1_val[14] reg1_val[15] reg1_val[16] reg1_val[17]
+ reg1_val[18] reg1_val[19] reg1_val[1] reg1_val[20] reg1_val[21] reg1_val[22] reg1_val[23]
+ reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27] reg1_val[28] reg1_val[29] reg1_val[2]
+ reg1_val[30] reg1_val[31] reg1_val[3] reg1_val[4] reg1_val[5] reg1_val[6] reg1_val[7]
+ reg1_val[8] reg1_val[9] reg2_idx[0] reg2_idx[1] reg2_idx[2] reg2_idx[3] reg2_idx[4]
+ reg2_idx[5] reg2_val[0] reg2_val[10] reg2_val[11] reg2_val[12] reg2_val[13] reg2_val[14]
+ reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18] reg2_val[19] reg2_val[1] reg2_val[20]
+ reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24] reg2_val[25] reg2_val[26] reg2_val[27]
+ reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30] reg2_val[31] reg2_val[3] reg2_val[4]
+ reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8] reg2_val[9] rst sign_extend take_branch
+ vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for icache abstract view
.subckt icache cache_entry[0] cache_entry[100] cache_entry[101] cache_entry[102] cache_entry[103]
+ cache_entry[104] cache_entry[105] cache_entry[106] cache_entry[107] cache_entry[108]
+ cache_entry[109] cache_entry[10] cache_entry[110] cache_entry[111] cache_entry[112]
+ cache_entry[113] cache_entry[114] cache_entry[115] cache_entry[116] cache_entry[117]
+ cache_entry[118] cache_entry[119] cache_entry[11] cache_entry[120] cache_entry[121]
+ cache_entry[122] cache_entry[123] cache_entry[124] cache_entry[125] cache_entry[126]
+ cache_entry[127] cache_entry[12] cache_entry[13] cache_entry[14] cache_entry[15]
+ cache_entry[16] cache_entry[17] cache_entry[18] cache_entry[19] cache_entry[1] cache_entry[20]
+ cache_entry[21] cache_entry[22] cache_entry[23] cache_entry[24] cache_entry[25]
+ cache_entry[26] cache_entry[27] cache_entry[28] cache_entry[29] cache_entry[2] cache_entry[30]
+ cache_entry[31] cache_entry[32] cache_entry[33] cache_entry[34] cache_entry[35]
+ cache_entry[36] cache_entry[37] cache_entry[38] cache_entry[39] cache_entry[3] cache_entry[40]
+ cache_entry[41] cache_entry[42] cache_entry[43] cache_entry[44] cache_entry[45]
+ cache_entry[46] cache_entry[47] cache_entry[48] cache_entry[49] cache_entry[4] cache_entry[50]
+ cache_entry[51] cache_entry[52] cache_entry[53] cache_entry[54] cache_entry[55]
+ cache_entry[56] cache_entry[57] cache_entry[58] cache_entry[59] cache_entry[5] cache_entry[60]
+ cache_entry[61] cache_entry[62] cache_entry[63] cache_entry[64] cache_entry[65]
+ cache_entry[66] cache_entry[67] cache_entry[68] cache_entry[69] cache_entry[6] cache_entry[70]
+ cache_entry[71] cache_entry[72] cache_entry[73] cache_entry[74] cache_entry[75]
+ cache_entry[76] cache_entry[77] cache_entry[78] cache_entry[79] cache_entry[7] cache_entry[80]
+ cache_entry[81] cache_entry[82] cache_entry[83] cache_entry[84] cache_entry[85]
+ cache_entry[86] cache_entry[87] cache_entry[88] cache_entry[89] cache_entry[8] cache_entry[90]
+ cache_entry[91] cache_entry[92] cache_entry[93] cache_entry[94] cache_entry[95]
+ cache_entry[96] cache_entry[97] cache_entry[98] cache_entry[99] cache_entry[9] cache_hit
+ curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13] curr_PC[14] curr_PC[15]
+ curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1] curr_PC[20] curr_PC[21]
+ curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26] curr_PC[27] curr_PC[2]
+ curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8] curr_PC[9] entry_valid
+ invalidate new_entry[0] new_entry[100] new_entry[101] new_entry[102] new_entry[103]
+ new_entry[104] new_entry[105] new_entry[106] new_entry[107] new_entry[108] new_entry[109]
+ new_entry[10] new_entry[110] new_entry[111] new_entry[112] new_entry[113] new_entry[114]
+ new_entry[115] new_entry[116] new_entry[117] new_entry[118] new_entry[119] new_entry[11]
+ new_entry[120] new_entry[121] new_entry[122] new_entry[123] new_entry[124] new_entry[125]
+ new_entry[126] new_entry[127] new_entry[12] new_entry[13] new_entry[14] new_entry[15]
+ new_entry[16] new_entry[17] new_entry[18] new_entry[19] new_entry[1] new_entry[20]
+ new_entry[21] new_entry[22] new_entry[23] new_entry[24] new_entry[25] new_entry[26]
+ new_entry[27] new_entry[28] new_entry[29] new_entry[2] new_entry[30] new_entry[31]
+ new_entry[32] new_entry[33] new_entry[34] new_entry[35] new_entry[36] new_entry[37]
+ new_entry[38] new_entry[39] new_entry[3] new_entry[40] new_entry[41] new_entry[42]
+ new_entry[43] new_entry[44] new_entry[45] new_entry[46] new_entry[47] new_entry[48]
+ new_entry[49] new_entry[4] new_entry[50] new_entry[51] new_entry[52] new_entry[53]
+ new_entry[54] new_entry[55] new_entry[56] new_entry[57] new_entry[58] new_entry[59]
+ new_entry[5] new_entry[60] new_entry[61] new_entry[62] new_entry[63] new_entry[64]
+ new_entry[65] new_entry[66] new_entry[67] new_entry[68] new_entry[69] new_entry[6]
+ new_entry[70] new_entry[71] new_entry[72] new_entry[73] new_entry[74] new_entry[75]
+ new_entry[76] new_entry[77] new_entry[78] new_entry[79] new_entry[7] new_entry[80]
+ new_entry[81] new_entry[82] new_entry[83] new_entry[84] new_entry[85] new_entry[86]
+ new_entry[87] new_entry[88] new_entry[89] new_entry[8] new_entry[90] new_entry[91]
+ new_entry[92] new_entry[93] new_entry[94] new_entry[95] new_entry[96] new_entry[97]
+ new_entry[98] new_entry[99] new_entry[9] rst vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_8x305 abstract view
.subckt wrapped_8x305 custom_settings[0] custom_settings[1] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vccd1
+ vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for scrapcpu abstract view
.subckt scrapcpu io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for multiplexer abstract view
.subckt multiplexer cap_addr[0] cap_addr[1] cap_addr[2] cap_addr[3] cap_addr[4] cap_addr[5]
+ cap_addr[6] cap_addr[7] cap_addr[8] cap_io_in[0] cap_io_in[1] cap_io_in[2] cap_io_in[3]
+ cap_io_in[4] cap_io_in[5] cap_io_in[6] cap_io_in[7] cap_io_in[8] custom_settings[0]
+ custom_settings[10] custom_settings[11] custom_settings[12] custom_settings[13]
+ custom_settings[14] custom_settings[15] custom_settings[16] custom_settings[17]
+ custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20] custom_settings[21]
+ custom_settings[22] custom_settings[23] custom_settings[24] custom_settings[25]
+ custom_settings[26] custom_settings[27] custom_settings[28] custom_settings[29]
+ custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3] custom_settings[4]
+ custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8] custom_settings[9]
+ io_in_0 io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2]
+ io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_oeb_6502
+ io_oeb_8x305[0] io_oeb_8x305[1] io_oeb_8x305[2] io_oeb_8x305[3] io_oeb_8x305[4]
+ io_oeb_as1802 io_oeb_scrapcpu[0] io_oeb_scrapcpu[10] io_oeb_scrapcpu[11] io_oeb_scrapcpu[12]
+ io_oeb_scrapcpu[13] io_oeb_scrapcpu[14] io_oeb_scrapcpu[15] io_oeb_scrapcpu[16]
+ io_oeb_scrapcpu[17] io_oeb_scrapcpu[18] io_oeb_scrapcpu[19] io_oeb_scrapcpu[1] io_oeb_scrapcpu[20]
+ io_oeb_scrapcpu[21] io_oeb_scrapcpu[22] io_oeb_scrapcpu[23] io_oeb_scrapcpu[24]
+ io_oeb_scrapcpu[25] io_oeb_scrapcpu[26] io_oeb_scrapcpu[27] io_oeb_scrapcpu[28]
+ io_oeb_scrapcpu[29] io_oeb_scrapcpu[2] io_oeb_scrapcpu[30] io_oeb_scrapcpu[31] io_oeb_scrapcpu[32]
+ io_oeb_scrapcpu[33] io_oeb_scrapcpu[34] io_oeb_scrapcpu[35] io_oeb_scrapcpu[3] io_oeb_scrapcpu[4]
+ io_oeb_scrapcpu[5] io_oeb_scrapcpu[6] io_oeb_scrapcpu[7] io_oeb_scrapcpu[8] io_oeb_scrapcpu[9]
+ io_oeb_vliw[0] io_oeb_vliw[10] io_oeb_vliw[11] io_oeb_vliw[12] io_oeb_vliw[13] io_oeb_vliw[14]
+ io_oeb_vliw[15] io_oeb_vliw[16] io_oeb_vliw[17] io_oeb_vliw[18] io_oeb_vliw[19]
+ io_oeb_vliw[1] io_oeb_vliw[20] io_oeb_vliw[21] io_oeb_vliw[22] io_oeb_vliw[23] io_oeb_vliw[24]
+ io_oeb_vliw[25] io_oeb_vliw[26] io_oeb_vliw[27] io_oeb_vliw[28] io_oeb_vliw[29]
+ io_oeb_vliw[2] io_oeb_vliw[30] io_oeb_vliw[31] io_oeb_vliw[32] io_oeb_vliw[33] io_oeb_vliw[34]
+ io_oeb_vliw[35] io_oeb_vliw[3] io_oeb_vliw[4] io_oeb_vliw[5] io_oeb_vliw[6] io_oeb_vliw[7]
+ io_oeb_vliw[8] io_oeb_vliw[9] io_oeb_z80[0] io_oeb_z80[10] io_oeb_z80[11] io_oeb_z80[12]
+ io_oeb_z80[13] io_oeb_z80[14] io_oeb_z80[15] io_oeb_z80[16] io_oeb_z80[17] io_oeb_z80[18]
+ io_oeb_z80[19] io_oeb_z80[1] io_oeb_z80[20] io_oeb_z80[21] io_oeb_z80[22] io_oeb_z80[23]
+ io_oeb_z80[24] io_oeb_z80[25] io_oeb_z80[26] io_oeb_z80[27] io_oeb_z80[28] io_oeb_z80[29]
+ io_oeb_z80[2] io_oeb_z80[30] io_oeb_z80[31] io_oeb_z80[32] io_oeb_z80[33] io_oeb_z80[34]
+ io_oeb_z80[35] io_oeb_z80[3] io_oeb_z80[4] io_oeb_z80[5] io_oeb_z80[6] io_oeb_z80[7]
+ io_oeb_z80[8] io_oeb_z80[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8]
+ io_out[9] io_out_6502[0] io_out_6502[10] io_out_6502[11] io_out_6502[12] io_out_6502[13]
+ io_out_6502[14] io_out_6502[15] io_out_6502[16] io_out_6502[17] io_out_6502[18]
+ io_out_6502[19] io_out_6502[1] io_out_6502[20] io_out_6502[21] io_out_6502[22] io_out_6502[23]
+ io_out_6502[24] io_out_6502[25] io_out_6502[26] io_out_6502[27] io_out_6502[28]
+ io_out_6502[29] io_out_6502[2] io_out_6502[30] io_out_6502[31] io_out_6502[32] io_out_6502[33]
+ io_out_6502[34] io_out_6502[35] io_out_6502[3] io_out_6502[4] io_out_6502[5] io_out_6502[6]
+ io_out_6502[7] io_out_6502[8] io_out_6502[9] io_out_8x305[0] io_out_8x305[10] io_out_8x305[11]
+ io_out_8x305[12] io_out_8x305[13] io_out_8x305[14] io_out_8x305[15] io_out_8x305[16]
+ io_out_8x305[17] io_out_8x305[18] io_out_8x305[19] io_out_8x305[1] io_out_8x305[20]
+ io_out_8x305[21] io_out_8x305[22] io_out_8x305[23] io_out_8x305[24] io_out_8x305[25]
+ io_out_8x305[26] io_out_8x305[27] io_out_8x305[28] io_out_8x305[29] io_out_8x305[2]
+ io_out_8x305[30] io_out_8x305[31] io_out_8x305[32] io_out_8x305[33] io_out_8x305[34]
+ io_out_8x305[35] io_out_8x305[3] io_out_8x305[4] io_out_8x305[5] io_out_8x305[6]
+ io_out_8x305[7] io_out_8x305[8] io_out_8x305[9] io_out_as1802[0] io_out_as1802[10]
+ io_out_as1802[11] io_out_as1802[12] io_out_as1802[13] io_out_as1802[14] io_out_as1802[15]
+ io_out_as1802[16] io_out_as1802[17] io_out_as1802[18] io_out_as1802[19] io_out_as1802[1]
+ io_out_as1802[20] io_out_as1802[21] io_out_as1802[22] io_out_as1802[23] io_out_as1802[24]
+ io_out_as1802[25] io_out_as1802[26] io_out_as1802[27] io_out_as1802[28] io_out_as1802[29]
+ io_out_as1802[2] io_out_as1802[30] io_out_as1802[31] io_out_as1802[32] io_out_as1802[33]
+ io_out_as1802[34] io_out_as1802[35] io_out_as1802[3] io_out_as1802[4] io_out_as1802[5]
+ io_out_as1802[6] io_out_as1802[7] io_out_as1802[8] io_out_as1802[9] io_out_scrapcpu[0]
+ io_out_scrapcpu[10] io_out_scrapcpu[11] io_out_scrapcpu[12] io_out_scrapcpu[13]
+ io_out_scrapcpu[14] io_out_scrapcpu[15] io_out_scrapcpu[16] io_out_scrapcpu[17]
+ io_out_scrapcpu[18] io_out_scrapcpu[19] io_out_scrapcpu[1] io_out_scrapcpu[20] io_out_scrapcpu[21]
+ io_out_scrapcpu[22] io_out_scrapcpu[23] io_out_scrapcpu[24] io_out_scrapcpu[25]
+ io_out_scrapcpu[26] io_out_scrapcpu[27] io_out_scrapcpu[28] io_out_scrapcpu[29]
+ io_out_scrapcpu[2] io_out_scrapcpu[30] io_out_scrapcpu[31] io_out_scrapcpu[32] io_out_scrapcpu[33]
+ io_out_scrapcpu[34] io_out_scrapcpu[35] io_out_scrapcpu[3] io_out_scrapcpu[4] io_out_scrapcpu[5]
+ io_out_scrapcpu[6] io_out_scrapcpu[7] io_out_scrapcpu[8] io_out_scrapcpu[9] io_out_vliw[0]
+ io_out_vliw[10] io_out_vliw[11] io_out_vliw[12] io_out_vliw[13] io_out_vliw[14]
+ io_out_vliw[15] io_out_vliw[16] io_out_vliw[17] io_out_vliw[18] io_out_vliw[19]
+ io_out_vliw[1] io_out_vliw[20] io_out_vliw[21] io_out_vliw[22] io_out_vliw[23] io_out_vliw[24]
+ io_out_vliw[25] io_out_vliw[26] io_out_vliw[27] io_out_vliw[28] io_out_vliw[29]
+ io_out_vliw[2] io_out_vliw[30] io_out_vliw[31] io_out_vliw[32] io_out_vliw[33] io_out_vliw[34]
+ io_out_vliw[35] io_out_vliw[3] io_out_vliw[4] io_out_vliw[5] io_out_vliw[6] io_out_vliw[7]
+ io_out_vliw[8] io_out_vliw[9] io_out_z80[0] io_out_z80[10] io_out_z80[11] io_out_z80[12]
+ io_out_z80[13] io_out_z80[14] io_out_z80[15] io_out_z80[16] io_out_z80[17] io_out_z80[18]
+ io_out_z80[19] io_out_z80[1] io_out_z80[20] io_out_z80[21] io_out_z80[22] io_out_z80[23]
+ io_out_z80[24] io_out_z80[25] io_out_z80[26] io_out_z80[27] io_out_z80[28] io_out_z80[29]
+ io_out_z80[2] io_out_z80[30] io_out_z80[31] io_out_z80[32] io_out_z80[33] io_out_z80[34]
+ io_out_z80[35] io_out_z80[3] io_out_z80[4] io_out_z80[5] io_out_z80[6] io_out_z80[7]
+ io_out_z80[8] io_out_z80[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] rst_6502 rst_8x305 rst_as1802 rst_scrapcpu
+ rst_vliw rst_z80 vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for vliw abstract view
.subckt vliw cache_PC[0] cache_PC[10] cache_PC[11] cache_PC[12] cache_PC[13] cache_PC[14]
+ cache_PC[15] cache_PC[16] cache_PC[17] cache_PC[18] cache_PC[19] cache_PC[1] cache_PC[20]
+ cache_PC[21] cache_PC[22] cache_PC[23] cache_PC[24] cache_PC[25] cache_PC[26] cache_PC[27]
+ cache_PC[2] cache_PC[3] cache_PC[4] cache_PC[5] cache_PC[6] cache_PC[7] cache_PC[8]
+ cache_PC[9] cache_entry[0] cache_entry[100] cache_entry[101] cache_entry[102] cache_entry[103]
+ cache_entry[104] cache_entry[105] cache_entry[106] cache_entry[107] cache_entry[108]
+ cache_entry[109] cache_entry[10] cache_entry[110] cache_entry[111] cache_entry[112]
+ cache_entry[113] cache_entry[114] cache_entry[115] cache_entry[116] cache_entry[117]
+ cache_entry[118] cache_entry[119] cache_entry[11] cache_entry[120] cache_entry[121]
+ cache_entry[122] cache_entry[123] cache_entry[124] cache_entry[125] cache_entry[126]
+ cache_entry[127] cache_entry[12] cache_entry[13] cache_entry[14] cache_entry[15]
+ cache_entry[16] cache_entry[17] cache_entry[18] cache_entry[19] cache_entry[1] cache_entry[20]
+ cache_entry[21] cache_entry[22] cache_entry[23] cache_entry[24] cache_entry[25]
+ cache_entry[26] cache_entry[27] cache_entry[28] cache_entry[29] cache_entry[2] cache_entry[30]
+ cache_entry[31] cache_entry[32] cache_entry[33] cache_entry[34] cache_entry[35]
+ cache_entry[36] cache_entry[37] cache_entry[38] cache_entry[39] cache_entry[3] cache_entry[40]
+ cache_entry[41] cache_entry[42] cache_entry[43] cache_entry[44] cache_entry[45]
+ cache_entry[46] cache_entry[47] cache_entry[48] cache_entry[49] cache_entry[4] cache_entry[50]
+ cache_entry[51] cache_entry[52] cache_entry[53] cache_entry[54] cache_entry[55]
+ cache_entry[56] cache_entry[57] cache_entry[58] cache_entry[59] cache_entry[5] cache_entry[60]
+ cache_entry[61] cache_entry[62] cache_entry[63] cache_entry[64] cache_entry[65]
+ cache_entry[66] cache_entry[67] cache_entry[68] cache_entry[69] cache_entry[6] cache_entry[70]
+ cache_entry[71] cache_entry[72] cache_entry[73] cache_entry[74] cache_entry[75]
+ cache_entry[76] cache_entry[77] cache_entry[78] cache_entry[79] cache_entry[7] cache_entry[80]
+ cache_entry[81] cache_entry[82] cache_entry[83] cache_entry[84] cache_entry[85]
+ cache_entry[86] cache_entry[87] cache_entry[88] cache_entry[89] cache_entry[8] cache_entry[90]
+ cache_entry[91] cache_entry[92] cache_entry[93] cache_entry[94] cache_entry[95]
+ cache_entry[96] cache_entry[97] cache_entry[98] cache_entry[99] cache_entry[9] cache_entry_valid
+ cache_hit cache_invalidate cache_new_entry[0] cache_new_entry[100] cache_new_entry[101]
+ cache_new_entry[102] cache_new_entry[103] cache_new_entry[104] cache_new_entry[105]
+ cache_new_entry[106] cache_new_entry[107] cache_new_entry[108] cache_new_entry[109]
+ cache_new_entry[10] cache_new_entry[110] cache_new_entry[111] cache_new_entry[112]
+ cache_new_entry[113] cache_new_entry[114] cache_new_entry[115] cache_new_entry[116]
+ cache_new_entry[117] cache_new_entry[118] cache_new_entry[119] cache_new_entry[11]
+ cache_new_entry[120] cache_new_entry[121] cache_new_entry[122] cache_new_entry[123]
+ cache_new_entry[124] cache_new_entry[125] cache_new_entry[126] cache_new_entry[127]
+ cache_new_entry[12] cache_new_entry[13] cache_new_entry[14] cache_new_entry[15]
+ cache_new_entry[16] cache_new_entry[17] cache_new_entry[18] cache_new_entry[19]
+ cache_new_entry[1] cache_new_entry[20] cache_new_entry[21] cache_new_entry[22] cache_new_entry[23]
+ cache_new_entry[24] cache_new_entry[25] cache_new_entry[26] cache_new_entry[27]
+ cache_new_entry[28] cache_new_entry[29] cache_new_entry[2] cache_new_entry[30] cache_new_entry[31]
+ cache_new_entry[32] cache_new_entry[33] cache_new_entry[34] cache_new_entry[35]
+ cache_new_entry[36] cache_new_entry[37] cache_new_entry[38] cache_new_entry[39]
+ cache_new_entry[3] cache_new_entry[40] cache_new_entry[41] cache_new_entry[42] cache_new_entry[43]
+ cache_new_entry[44] cache_new_entry[45] cache_new_entry[46] cache_new_entry[47]
+ cache_new_entry[48] cache_new_entry[49] cache_new_entry[4] cache_new_entry[50] cache_new_entry[51]
+ cache_new_entry[52] cache_new_entry[53] cache_new_entry[54] cache_new_entry[55]
+ cache_new_entry[56] cache_new_entry[57] cache_new_entry[58] cache_new_entry[59]
+ cache_new_entry[5] cache_new_entry[60] cache_new_entry[61] cache_new_entry[62] cache_new_entry[63]
+ cache_new_entry[64] cache_new_entry[65] cache_new_entry[66] cache_new_entry[67]
+ cache_new_entry[68] cache_new_entry[69] cache_new_entry[6] cache_new_entry[70] cache_new_entry[71]
+ cache_new_entry[72] cache_new_entry[73] cache_new_entry[74] cache_new_entry[75]
+ cache_new_entry[76] cache_new_entry[77] cache_new_entry[78] cache_new_entry[79]
+ cache_new_entry[7] cache_new_entry[80] cache_new_entry[81] cache_new_entry[82] cache_new_entry[83]
+ cache_new_entry[84] cache_new_entry[85] cache_new_entry[86] cache_new_entry[87]
+ cache_new_entry[88] cache_new_entry[89] cache_new_entry[8] cache_new_entry[90] cache_new_entry[91]
+ cache_new_entry[92] cache_new_entry[93] cache_new_entry[94] cache_new_entry[95]
+ cache_new_entry[96] cache_new_entry[97] cache_new_entry[98] cache_new_entry[99]
+ cache_new_entry[9] cache_rst curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] custom_settings[0] custom_settings[1] custom_settings[2] custom_settings[3]
+ custom_settings[4] dest_idx0[0] dest_idx0[1] dest_idx0[2] dest_idx0[3] dest_idx0[4]
+ dest_idx0[5] dest_idx1[0] dest_idx1[1] dest_idx1[2] dest_idx1[3] dest_idx1[4] dest_idx1[5]
+ dest_idx2[0] dest_idx2[1] dest_idx2[2] dest_idx2[3] dest_idx2[4] dest_idx2[5] dest_mask0[0]
+ dest_mask0[1] dest_mask1[0] dest_mask1[1] dest_mask2[0] dest_mask2[1] dest_pred0[0]
+ dest_pred0[1] dest_pred0[2] dest_pred1[0] dest_pred1[1] dest_pred1[2] dest_pred2[0]
+ dest_pred2[1] dest_pred2[2] dest_pred_val0 dest_pred_val1 dest_pred_val2 dest_val0[0]
+ dest_val0[10] dest_val0[11] dest_val0[12] dest_val0[13] dest_val0[14] dest_val0[15]
+ dest_val0[16] dest_val0[17] dest_val0[18] dest_val0[19] dest_val0[1] dest_val0[20]
+ dest_val0[21] dest_val0[22] dest_val0[23] dest_val0[24] dest_val0[25] dest_val0[26]
+ dest_val0[27] dest_val0[28] dest_val0[29] dest_val0[2] dest_val0[30] dest_val0[31]
+ dest_val0[3] dest_val0[4] dest_val0[5] dest_val0[6] dest_val0[7] dest_val0[8] dest_val0[9]
+ dest_val1[0] dest_val1[10] dest_val1[11] dest_val1[12] dest_val1[13] dest_val1[14]
+ dest_val1[15] dest_val1[16] dest_val1[17] dest_val1[18] dest_val1[19] dest_val1[1]
+ dest_val1[20] dest_val1[21] dest_val1[22] dest_val1[23] dest_val1[24] dest_val1[25]
+ dest_val1[26] dest_val1[27] dest_val1[28] dest_val1[29] dest_val1[2] dest_val1[30]
+ dest_val1[31] dest_val1[3] dest_val1[4] dest_val1[5] dest_val1[6] dest_val1[7] dest_val1[8]
+ dest_val1[9] dest_val2[0] dest_val2[10] dest_val2[11] dest_val2[12] dest_val2[13]
+ dest_val2[14] dest_val2[15] dest_val2[16] dest_val2[17] dest_val2[18] dest_val2[19]
+ dest_val2[1] dest_val2[20] dest_val2[21] dest_val2[22] dest_val2[23] dest_val2[24]
+ dest_val2[25] dest_val2[26] dest_val2[27] dest_val2[28] dest_val2[29] dest_val2[2]
+ dest_val2[30] dest_val2[31] dest_val2[3] dest_val2[4] dest_val2[5] dest_val2[6]
+ dest_val2[7] dest_val2[8] dest_val2[9] eu0_busy eu0_instruction[0] eu0_instruction[10]
+ eu0_instruction[11] eu0_instruction[12] eu0_instruction[13] eu0_instruction[14]
+ eu0_instruction[15] eu0_instruction[16] eu0_instruction[17] eu0_instruction[18]
+ eu0_instruction[19] eu0_instruction[1] eu0_instruction[20] eu0_instruction[21] eu0_instruction[22]
+ eu0_instruction[23] eu0_instruction[24] eu0_instruction[25] eu0_instruction[26]
+ eu0_instruction[27] eu0_instruction[28] eu0_instruction[29] eu0_instruction[2] eu0_instruction[30]
+ eu0_instruction[31] eu0_instruction[32] eu0_instruction[33] eu0_instruction[34]
+ eu0_instruction[35] eu0_instruction[36] eu0_instruction[37] eu0_instruction[38]
+ eu0_instruction[39] eu0_instruction[3] eu0_instruction[40] eu0_instruction[41] eu0_instruction[4]
+ eu0_instruction[5] eu0_instruction[6] eu0_instruction[7] eu0_instruction[8] eu0_instruction[9]
+ eu1_busy eu1_instruction[0] eu1_instruction[10] eu1_instruction[11] eu1_instruction[12]
+ eu1_instruction[13] eu1_instruction[14] eu1_instruction[15] eu1_instruction[16]
+ eu1_instruction[17] eu1_instruction[18] eu1_instruction[19] eu1_instruction[1] eu1_instruction[20]
+ eu1_instruction[21] eu1_instruction[22] eu1_instruction[23] eu1_instruction[24]
+ eu1_instruction[25] eu1_instruction[26] eu1_instruction[27] eu1_instruction[28]
+ eu1_instruction[29] eu1_instruction[2] eu1_instruction[30] eu1_instruction[31] eu1_instruction[32]
+ eu1_instruction[33] eu1_instruction[34] eu1_instruction[35] eu1_instruction[36]
+ eu1_instruction[37] eu1_instruction[38] eu1_instruction[39] eu1_instruction[3] eu1_instruction[40]
+ eu1_instruction[41] eu1_instruction[4] eu1_instruction[5] eu1_instruction[6] eu1_instruction[7]
+ eu1_instruction[8] eu1_instruction[9] eu2_busy eu2_instruction[0] eu2_instruction[10]
+ eu2_instruction[11] eu2_instruction[12] eu2_instruction[13] eu2_instruction[14]
+ eu2_instruction[15] eu2_instruction[16] eu2_instruction[17] eu2_instruction[18]
+ eu2_instruction[19] eu2_instruction[1] eu2_instruction[20] eu2_instruction[21] eu2_instruction[22]
+ eu2_instruction[23] eu2_instruction[24] eu2_instruction[25] eu2_instruction[26]
+ eu2_instruction[27] eu2_instruction[28] eu2_instruction[29] eu2_instruction[2] eu2_instruction[30]
+ eu2_instruction[31] eu2_instruction[32] eu2_instruction[33] eu2_instruction[34]
+ eu2_instruction[35] eu2_instruction[36] eu2_instruction[37] eu2_instruction[38]
+ eu2_instruction[39] eu2_instruction[3] eu2_instruction[40] eu2_instruction[41] eu2_instruction[4]
+ eu2_instruction[5] eu2_instruction[6] eu2_instruction[7] eu2_instruction[8] eu2_instruction[9]
+ int_return0 int_return1 int_return2 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] is_load0 is_load1 is_load2 is_store0 is_store1
+ is_store2 loadstore_address0[0] loadstore_address0[10] loadstore_address0[11] loadstore_address0[12]
+ loadstore_address0[13] loadstore_address0[14] loadstore_address0[15] loadstore_address0[16]
+ loadstore_address0[17] loadstore_address0[18] loadstore_address0[19] loadstore_address0[1]
+ loadstore_address0[20] loadstore_address0[21] loadstore_address0[22] loadstore_address0[23]
+ loadstore_address0[24] loadstore_address0[25] loadstore_address0[26] loadstore_address0[27]
+ loadstore_address0[28] loadstore_address0[29] loadstore_address0[2] loadstore_address0[30]
+ loadstore_address0[31] loadstore_address0[3] loadstore_address0[4] loadstore_address0[5]
+ loadstore_address0[6] loadstore_address0[7] loadstore_address0[8] loadstore_address0[9]
+ loadstore_address1[0] loadstore_address1[10] loadstore_address1[11] loadstore_address1[12]
+ loadstore_address1[13] loadstore_address1[14] loadstore_address1[15] loadstore_address1[16]
+ loadstore_address1[17] loadstore_address1[18] loadstore_address1[19] loadstore_address1[1]
+ loadstore_address1[20] loadstore_address1[21] loadstore_address1[22] loadstore_address1[23]
+ loadstore_address1[24] loadstore_address1[25] loadstore_address1[26] loadstore_address1[27]
+ loadstore_address1[28] loadstore_address1[29] loadstore_address1[2] loadstore_address1[30]
+ loadstore_address1[31] loadstore_address1[3] loadstore_address1[4] loadstore_address1[5]
+ loadstore_address1[6] loadstore_address1[7] loadstore_address1[8] loadstore_address1[9]
+ loadstore_address2[0] loadstore_address2[10] loadstore_address2[11] loadstore_address2[12]
+ loadstore_address2[13] loadstore_address2[14] loadstore_address2[15] loadstore_address2[16]
+ loadstore_address2[17] loadstore_address2[18] loadstore_address2[19] loadstore_address2[1]
+ loadstore_address2[20] loadstore_address2[21] loadstore_address2[22] loadstore_address2[23]
+ loadstore_address2[24] loadstore_address2[25] loadstore_address2[26] loadstore_address2[27]
+ loadstore_address2[28] loadstore_address2[29] loadstore_address2[2] loadstore_address2[30]
+ loadstore_address2[31] loadstore_address2[3] loadstore_address2[4] loadstore_address2[5]
+ loadstore_address2[6] loadstore_address2[7] loadstore_address2[8] loadstore_address2[9]
+ loadstore_dest0[0] loadstore_dest0[1] loadstore_dest0[2] loadstore_dest0[3] loadstore_dest0[4]
+ loadstore_dest0[5] loadstore_dest1[0] loadstore_dest1[1] loadstore_dest1[2] loadstore_dest1[3]
+ loadstore_dest1[4] loadstore_dest1[5] loadstore_dest2[0] loadstore_dest2[1] loadstore_dest2[2]
+ loadstore_dest2[3] loadstore_dest2[4] loadstore_dest2[5] loadstore_size0[0] loadstore_size0[1]
+ loadstore_size1[0] loadstore_size1[1] loadstore_size2[0] loadstore_size2[1] new_PC0[0]
+ new_PC0[10] new_PC0[11] new_PC0[12] new_PC0[13] new_PC0[14] new_PC0[15] new_PC0[16]
+ new_PC0[17] new_PC0[18] new_PC0[19] new_PC0[1] new_PC0[20] new_PC0[21] new_PC0[22]
+ new_PC0[23] new_PC0[24] new_PC0[25] new_PC0[26] new_PC0[27] new_PC0[2] new_PC0[3]
+ new_PC0[4] new_PC0[5] new_PC0[6] new_PC0[7] new_PC0[8] new_PC0[9] new_PC1[0] new_PC1[10]
+ new_PC1[11] new_PC1[12] new_PC1[13] new_PC1[14] new_PC1[15] new_PC1[16] new_PC1[17]
+ new_PC1[18] new_PC1[19] new_PC1[1] new_PC1[20] new_PC1[21] new_PC1[22] new_PC1[23]
+ new_PC1[24] new_PC1[25] new_PC1[26] new_PC1[27] new_PC1[2] new_PC1[3] new_PC1[4]
+ new_PC1[5] new_PC1[6] new_PC1[7] new_PC1[8] new_PC1[9] new_PC2[0] new_PC2[10] new_PC2[11]
+ new_PC2[12] new_PC2[13] new_PC2[14] new_PC2[15] new_PC2[16] new_PC2[17] new_PC2[18]
+ new_PC2[19] new_PC2[1] new_PC2[20] new_PC2[21] new_PC2[22] new_PC2[23] new_PC2[24]
+ new_PC2[25] new_PC2[26] new_PC2[27] new_PC2[2] new_PC2[3] new_PC2[4] new_PC2[5]
+ new_PC2[6] new_PC2[7] new_PC2[8] new_PC2[9] pred_idx0[0] pred_idx0[1] pred_idx0[2]
+ pred_idx1[0] pred_idx1[1] pred_idx1[2] pred_idx2[0] pred_idx2[1] pred_idx2[2] pred_val0
+ pred_val1 pred_val2 reg1_idx0[0] reg1_idx0[1] reg1_idx0[2] reg1_idx0[3] reg1_idx0[4]
+ reg1_idx0[5] reg1_idx1[0] reg1_idx1[1] reg1_idx1[2] reg1_idx1[3] reg1_idx1[4] reg1_idx1[5]
+ reg1_idx2[0] reg1_idx2[1] reg1_idx2[2] reg1_idx2[3] reg1_idx2[4] reg1_idx2[5] reg1_val0[0]
+ reg1_val0[10] reg1_val0[11] reg1_val0[12] reg1_val0[13] reg1_val0[14] reg1_val0[15]
+ reg1_val0[16] reg1_val0[17] reg1_val0[18] reg1_val0[19] reg1_val0[1] reg1_val0[20]
+ reg1_val0[21] reg1_val0[22] reg1_val0[23] reg1_val0[24] reg1_val0[25] reg1_val0[26]
+ reg1_val0[27] reg1_val0[28] reg1_val0[29] reg1_val0[2] reg1_val0[30] reg1_val0[31]
+ reg1_val0[3] reg1_val0[4] reg1_val0[5] reg1_val0[6] reg1_val0[7] reg1_val0[8] reg1_val0[9]
+ reg1_val1[0] reg1_val1[10] reg1_val1[11] reg1_val1[12] reg1_val1[13] reg1_val1[14]
+ reg1_val1[15] reg1_val1[16] reg1_val1[17] reg1_val1[18] reg1_val1[19] reg1_val1[1]
+ reg1_val1[20] reg1_val1[21] reg1_val1[22] reg1_val1[23] reg1_val1[24] reg1_val1[25]
+ reg1_val1[26] reg1_val1[27] reg1_val1[28] reg1_val1[29] reg1_val1[2] reg1_val1[30]
+ reg1_val1[31] reg1_val1[3] reg1_val1[4] reg1_val1[5] reg1_val1[6] reg1_val1[7] reg1_val1[8]
+ reg1_val1[9] reg1_val2[0] reg1_val2[10] reg1_val2[11] reg1_val2[12] reg1_val2[13]
+ reg1_val2[14] reg1_val2[15] reg1_val2[16] reg1_val2[17] reg1_val2[18] reg1_val2[19]
+ reg1_val2[1] reg1_val2[20] reg1_val2[21] reg1_val2[22] reg1_val2[23] reg1_val2[24]
+ reg1_val2[25] reg1_val2[26] reg1_val2[27] reg1_val2[28] reg1_val2[29] reg1_val2[2]
+ reg1_val2[30] reg1_val2[31] reg1_val2[3] reg1_val2[4] reg1_val2[5] reg1_val2[6]
+ reg1_val2[7] reg1_val2[8] reg1_val2[9] reg2_idx0[0] reg2_idx0[1] reg2_idx0[2] reg2_idx0[3]
+ reg2_idx0[4] reg2_idx0[5] reg2_idx1[0] reg2_idx1[1] reg2_idx1[2] reg2_idx1[3] reg2_idx1[4]
+ reg2_idx1[5] reg2_idx2[0] reg2_idx2[1] reg2_idx2[2] reg2_idx2[3] reg2_idx2[4] reg2_idx2[5]
+ reg2_val0[0] reg2_val0[10] reg2_val0[11] reg2_val0[12] reg2_val0[13] reg2_val0[14]
+ reg2_val0[15] reg2_val0[16] reg2_val0[17] reg2_val0[18] reg2_val0[19] reg2_val0[1]
+ reg2_val0[20] reg2_val0[21] reg2_val0[22] reg2_val0[23] reg2_val0[24] reg2_val0[25]
+ reg2_val0[26] reg2_val0[27] reg2_val0[28] reg2_val0[29] reg2_val0[2] reg2_val0[30]
+ reg2_val0[31] reg2_val0[3] reg2_val0[4] reg2_val0[5] reg2_val0[6] reg2_val0[7] reg2_val0[8]
+ reg2_val0[9] reg2_val1[0] reg2_val1[10] reg2_val1[11] reg2_val1[12] reg2_val1[13]
+ reg2_val1[14] reg2_val1[15] reg2_val1[16] reg2_val1[17] reg2_val1[18] reg2_val1[19]
+ reg2_val1[1] reg2_val1[20] reg2_val1[21] reg2_val1[22] reg2_val1[23] reg2_val1[24]
+ reg2_val1[25] reg2_val1[26] reg2_val1[27] reg2_val1[28] reg2_val1[29] reg2_val1[2]
+ reg2_val1[30] reg2_val1[31] reg2_val1[3] reg2_val1[4] reg2_val1[5] reg2_val1[6]
+ reg2_val1[7] reg2_val1[8] reg2_val1[9] reg2_val2[0] reg2_val2[10] reg2_val2[11]
+ reg2_val2[12] reg2_val2[13] reg2_val2[14] reg2_val2[15] reg2_val2[16] reg2_val2[17]
+ reg2_val2[18] reg2_val2[19] reg2_val2[1] reg2_val2[20] reg2_val2[21] reg2_val2[22]
+ reg2_val2[23] reg2_val2[24] reg2_val2[25] reg2_val2[26] reg2_val2[27] reg2_val2[28]
+ reg2_val2[29] reg2_val2[2] reg2_val2[30] reg2_val2[31] reg2_val2[3] reg2_val2[4]
+ reg2_val2[5] reg2_val2[6] reg2_val2[7] reg2_val2[8] reg2_val2[9] rst_eu rst_n sign_extend0
+ sign_extend1 sign_extend2 take_branch0 take_branch1 take_branch2 vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_as1802 abstract view
.subckt wrapped_as1802 custom_settings[0] custom_settings[10] custom_settings[11]
+ custom_settings[12] custom_settings[13] custom_settings[14] custom_settings[15]
+ custom_settings[16] custom_settings[17] custom_settings[18] custom_settings[19]
+ custom_settings[1] custom_settings[20] custom_settings[21] custom_settings[22] custom_settings[23]
+ custom_settings[24] custom_settings[25] custom_settings[26] custom_settings[27]
+ custom_settings[28] custom_settings[29] custom_settings[2] custom_settings[3] custom_settings[4]
+ custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8] custom_settings[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9]
+ io_oeb io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_6502 abstract view
.subckt wrapped_6502 custom_settings[0] custom_settings[1] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24]
+ io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31]
+ io_out[32] io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for unused_tie abstract view
.subckt unused_tie irq[0] irq[1] irq[2] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[8] la_data_out[9] vccd1 vssd1 wb_clk_i wb_rst_i
.ends

* Black-box entry subcircuit for ci2406_z80 abstract view
.subckt ci2406_z80 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xeu1 eu1/busy eu2/curr_PC[0] eu2/curr_PC[10] eu2/curr_PC[11] eu2/curr_PC[12] eu2/curr_PC[13]
+ eu2/curr_PC[14] eu2/curr_PC[15] eu2/curr_PC[16] eu2/curr_PC[17] eu2/curr_PC[18]
+ eu2/curr_PC[19] eu2/curr_PC[1] eu2/curr_PC[20] eu2/curr_PC[21] eu2/curr_PC[22] eu2/curr_PC[23]
+ eu2/curr_PC[24] eu2/curr_PC[25] eu2/curr_PC[26] eu2/curr_PC[27] eu2/curr_PC[2] eu2/curr_PC[3]
+ eu2/curr_PC[4] eu2/curr_PC[5] eu2/curr_PC[6] eu2/curr_PC[7] eu2/curr_PC[8] eu2/curr_PC[9]
+ eu1/dest_idx[0] eu1/dest_idx[1] eu1/dest_idx[2] eu1/dest_idx[3] eu1/dest_idx[4]
+ eu1/dest_idx[5] eu1/dest_mask[0] eu1/dest_mask[1] eu1/dest_pred[0] eu1/dest_pred[1]
+ eu1/dest_pred[2] eu1/dest_pred_val eu1/dest_val[0] eu1/dest_val[10] eu1/dest_val[11]
+ eu1/dest_val[12] eu1/dest_val[13] eu1/dest_val[14] eu1/dest_val[15] eu1/dest_val[16]
+ eu1/dest_val[17] eu1/dest_val[18] eu1/dest_val[19] eu1/dest_val[1] eu1/dest_val[20]
+ eu1/dest_val[21] eu1/dest_val[22] eu1/dest_val[23] eu1/dest_val[24] eu1/dest_val[25]
+ eu1/dest_val[26] eu1/dest_val[27] eu1/dest_val[28] eu1/dest_val[29] eu1/dest_val[2]
+ eu1/dest_val[30] eu1/dest_val[31] eu1/dest_val[3] eu1/dest_val[4] eu1/dest_val[5]
+ eu1/dest_val[6] eu1/dest_val[7] eu1/dest_val[8] eu1/dest_val[9] eu1/instruction[0]
+ eu1/instruction[10] eu1/instruction[11] eu1/instruction[12] eu1/instruction[13]
+ eu1/instruction[14] eu1/instruction[15] eu1/instruction[16] eu1/instruction[17]
+ eu1/instruction[18] eu1/instruction[19] eu1/instruction[1] eu1/instruction[20] eu1/instruction[21]
+ eu1/instruction[22] eu1/instruction[23] eu1/instruction[24] eu1/instruction[25]
+ eu1/instruction[26] eu1/instruction[27] eu1/instruction[28] eu1/instruction[29]
+ eu1/instruction[2] eu1/instruction[30] eu1/instruction[31] eu1/instruction[32] eu1/instruction[33]
+ eu1/instruction[34] eu1/instruction[35] eu1/instruction[36] eu1/instruction[37]
+ eu1/instruction[38] eu1/instruction[39] eu1/instruction[3] eu1/instruction[40] eu1/instruction[41]
+ eu1/instruction[4] eu1/instruction[5] eu1/instruction[6] eu1/instruction[7] eu1/instruction[8]
+ eu1/instruction[9] eu1/int_return eu1/is_load eu1/is_store eu1/loadstore_address[0]
+ eu1/loadstore_address[10] eu1/loadstore_address[11] eu1/loadstore_address[12] eu1/loadstore_address[13]
+ eu1/loadstore_address[14] eu1/loadstore_address[15] eu1/loadstore_address[16] eu1/loadstore_address[17]
+ eu1/loadstore_address[18] eu1/loadstore_address[19] eu1/loadstore_address[1] eu1/loadstore_address[20]
+ eu1/loadstore_address[21] eu1/loadstore_address[22] eu1/loadstore_address[23] eu1/loadstore_address[24]
+ eu1/loadstore_address[25] eu1/loadstore_address[26] eu1/loadstore_address[27] eu1/loadstore_address[28]
+ eu1/loadstore_address[29] eu1/loadstore_address[2] eu1/loadstore_address[30] eu1/loadstore_address[31]
+ eu1/loadstore_address[3] eu1/loadstore_address[4] eu1/loadstore_address[5] eu1/loadstore_address[6]
+ eu1/loadstore_address[7] eu1/loadstore_address[8] eu1/loadstore_address[9] eu1/loadstore_dest[0]
+ eu1/loadstore_dest[1] eu1/loadstore_dest[2] eu1/loadstore_dest[3] eu1/loadstore_dest[4]
+ eu1/loadstore_dest[5] eu1/loadstore_size[0] eu1/loadstore_size[1] eu1/new_PC[0]
+ eu1/new_PC[10] eu1/new_PC[11] eu1/new_PC[12] eu1/new_PC[13] eu1/new_PC[14] eu1/new_PC[15]
+ eu1/new_PC[16] eu1/new_PC[17] eu1/new_PC[18] eu1/new_PC[19] eu1/new_PC[1] eu1/new_PC[20]
+ eu1/new_PC[21] eu1/new_PC[22] eu1/new_PC[23] eu1/new_PC[24] eu1/new_PC[25] eu1/new_PC[26]
+ eu1/new_PC[27] eu1/new_PC[2] eu1/new_PC[3] eu1/new_PC[4] eu1/new_PC[5] eu1/new_PC[6]
+ eu1/new_PC[7] eu1/new_PC[8] eu1/new_PC[9] eu1/pred_idx[0] eu1/pred_idx[1] eu1/pred_idx[2]
+ eu1/pred_val eu1/reg1_idx[0] eu1/reg1_idx[1] eu1/reg1_idx[2] eu1/reg1_idx[3] eu1/reg1_idx[4]
+ eu1/reg1_idx[5] eu1/reg1_val[0] eu1/reg1_val[10] eu1/reg1_val[11] eu1/reg1_val[12]
+ eu1/reg1_val[13] eu1/reg1_val[14] eu1/reg1_val[15] eu1/reg1_val[16] eu1/reg1_val[17]
+ eu1/reg1_val[18] eu1/reg1_val[19] eu1/reg1_val[1] eu1/reg1_val[20] eu1/reg1_val[21]
+ eu1/reg1_val[22] eu1/reg1_val[23] eu1/reg1_val[24] eu1/reg1_val[25] eu1/reg1_val[26]
+ eu1/reg1_val[27] eu1/reg1_val[28] eu1/reg1_val[29] eu1/reg1_val[2] eu1/reg1_val[30]
+ eu1/reg1_val[31] eu1/reg1_val[3] eu1/reg1_val[4] eu1/reg1_val[5] eu1/reg1_val[6]
+ eu1/reg1_val[7] eu1/reg1_val[8] eu1/reg1_val[9] eu1/reg2_idx[0] eu1/reg2_idx[1]
+ eu1/reg2_idx[2] eu1/reg2_idx[3] eu1/reg2_idx[4] eu1/reg2_idx[5] eu1/reg2_val[0]
+ eu1/reg2_val[10] eu1/reg2_val[11] eu1/reg2_val[12] eu1/reg2_val[13] eu1/reg2_val[14]
+ eu1/reg2_val[15] eu1/reg2_val[16] eu1/reg2_val[17] eu1/reg2_val[18] eu1/reg2_val[19]
+ eu1/reg2_val[1] eu1/reg2_val[20] eu1/reg2_val[21] eu1/reg2_val[22] eu1/reg2_val[23]
+ eu1/reg2_val[24] eu1/reg2_val[25] eu1/reg2_val[26] eu1/reg2_val[27] eu1/reg2_val[28]
+ eu1/reg2_val[29] eu1/reg2_val[2] eu1/reg2_val[30] eu1/reg2_val[31] eu1/reg2_val[3]
+ eu1/reg2_val[4] eu1/reg2_val[5] eu1/reg2_val[6] eu1/reg2_val[7] eu1/reg2_val[8]
+ eu1/reg2_val[9] eu2/rst eu1/sign_extend eu1/take_branch vccd1 vssd1 wb_clk_i execution_unit
Xeu0 eu0/busy eu2/curr_PC[0] eu2/curr_PC[10] eu2/curr_PC[11] eu2/curr_PC[12] eu2/curr_PC[13]
+ eu2/curr_PC[14] eu2/curr_PC[15] eu2/curr_PC[16] eu2/curr_PC[17] eu2/curr_PC[18]
+ eu2/curr_PC[19] eu2/curr_PC[1] eu2/curr_PC[20] eu2/curr_PC[21] eu2/curr_PC[22] eu2/curr_PC[23]
+ eu2/curr_PC[24] eu2/curr_PC[25] eu2/curr_PC[26] eu2/curr_PC[27] eu2/curr_PC[2] eu2/curr_PC[3]
+ eu2/curr_PC[4] eu2/curr_PC[5] eu2/curr_PC[6] eu2/curr_PC[7] eu2/curr_PC[8] eu2/curr_PC[9]
+ eu0/dest_idx[0] eu0/dest_idx[1] eu0/dest_idx[2] eu0/dest_idx[3] eu0/dest_idx[4]
+ eu0/dest_idx[5] eu0/dest_mask[0] eu0/dest_mask[1] eu0/dest_pred[0] eu0/dest_pred[1]
+ eu0/dest_pred[2] eu0/dest_pred_val eu0/dest_val[0] eu0/dest_val[10] eu0/dest_val[11]
+ eu0/dest_val[12] eu0/dest_val[13] eu0/dest_val[14] eu0/dest_val[15] eu0/dest_val[16]
+ eu0/dest_val[17] eu0/dest_val[18] eu0/dest_val[19] eu0/dest_val[1] eu0/dest_val[20]
+ eu0/dest_val[21] eu0/dest_val[22] eu0/dest_val[23] eu0/dest_val[24] eu0/dest_val[25]
+ eu0/dest_val[26] eu0/dest_val[27] eu0/dest_val[28] eu0/dest_val[29] eu0/dest_val[2]
+ eu0/dest_val[30] eu0/dest_val[31] eu0/dest_val[3] eu0/dest_val[4] eu0/dest_val[5]
+ eu0/dest_val[6] eu0/dest_val[7] eu0/dest_val[8] eu0/dest_val[9] eu0/instruction[0]
+ eu0/instruction[10] eu0/instruction[11] eu0/instruction[12] eu0/instruction[13]
+ eu0/instruction[14] eu0/instruction[15] eu0/instruction[16] eu0/instruction[17]
+ eu0/instruction[18] eu0/instruction[19] eu0/instruction[1] eu0/instruction[20] eu0/instruction[21]
+ eu0/instruction[22] eu0/instruction[23] eu0/instruction[24] eu0/instruction[25]
+ eu0/instruction[26] eu0/instruction[27] eu0/instruction[28] eu0/instruction[29]
+ eu0/instruction[2] eu0/instruction[30] eu0/instruction[31] eu0/instruction[32] eu0/instruction[33]
+ eu0/instruction[34] eu0/instruction[35] eu0/instruction[36] eu0/instruction[37]
+ eu0/instruction[38] eu0/instruction[39] eu0/instruction[3] eu0/instruction[40] eu0/instruction[41]
+ eu0/instruction[4] eu0/instruction[5] eu0/instruction[6] eu0/instruction[7] eu0/instruction[8]
+ eu0/instruction[9] eu0/int_return eu0/is_load eu0/is_store eu0/loadstore_address[0]
+ eu0/loadstore_address[10] eu0/loadstore_address[11] eu0/loadstore_address[12] eu0/loadstore_address[13]
+ eu0/loadstore_address[14] eu0/loadstore_address[15] eu0/loadstore_address[16] eu0/loadstore_address[17]
+ eu0/loadstore_address[18] eu0/loadstore_address[19] eu0/loadstore_address[1] eu0/loadstore_address[20]
+ eu0/loadstore_address[21] eu0/loadstore_address[22] eu0/loadstore_address[23] eu0/loadstore_address[24]
+ eu0/loadstore_address[25] eu0/loadstore_address[26] eu0/loadstore_address[27] eu0/loadstore_address[28]
+ eu0/loadstore_address[29] eu0/loadstore_address[2] eu0/loadstore_address[30] eu0/loadstore_address[31]
+ eu0/loadstore_address[3] eu0/loadstore_address[4] eu0/loadstore_address[5] eu0/loadstore_address[6]
+ eu0/loadstore_address[7] eu0/loadstore_address[8] eu0/loadstore_address[9] eu0/loadstore_dest[0]
+ eu0/loadstore_dest[1] eu0/loadstore_dest[2] eu0/loadstore_dest[3] eu0/loadstore_dest[4]
+ eu0/loadstore_dest[5] eu0/loadstore_size[0] eu0/loadstore_size[1] eu0/new_PC[0]
+ eu0/new_PC[10] eu0/new_PC[11] eu0/new_PC[12] eu0/new_PC[13] eu0/new_PC[14] eu0/new_PC[15]
+ eu0/new_PC[16] eu0/new_PC[17] eu0/new_PC[18] eu0/new_PC[19] eu0/new_PC[1] eu0/new_PC[20]
+ eu0/new_PC[21] eu0/new_PC[22] eu0/new_PC[23] eu0/new_PC[24] eu0/new_PC[25] eu0/new_PC[26]
+ eu0/new_PC[27] eu0/new_PC[2] eu0/new_PC[3] eu0/new_PC[4] eu0/new_PC[5] eu0/new_PC[6]
+ eu0/new_PC[7] eu0/new_PC[8] eu0/new_PC[9] eu0/pred_idx[0] eu0/pred_idx[1] eu0/pred_idx[2]
+ eu0/pred_val eu0/reg1_idx[0] eu0/reg1_idx[1] eu0/reg1_idx[2] eu0/reg1_idx[3] eu0/reg1_idx[4]
+ eu0/reg1_idx[5] eu0/reg1_val[0] eu0/reg1_val[10] eu0/reg1_val[11] eu0/reg1_val[12]
+ eu0/reg1_val[13] eu0/reg1_val[14] eu0/reg1_val[15] eu0/reg1_val[16] eu0/reg1_val[17]
+ eu0/reg1_val[18] eu0/reg1_val[19] eu0/reg1_val[1] eu0/reg1_val[20] eu0/reg1_val[21]
+ eu0/reg1_val[22] eu0/reg1_val[23] eu0/reg1_val[24] eu0/reg1_val[25] eu0/reg1_val[26]
+ eu0/reg1_val[27] eu0/reg1_val[28] eu0/reg1_val[29] eu0/reg1_val[2] eu0/reg1_val[30]
+ eu0/reg1_val[31] eu0/reg1_val[3] eu0/reg1_val[4] eu0/reg1_val[5] eu0/reg1_val[6]
+ eu0/reg1_val[7] eu0/reg1_val[8] eu0/reg1_val[9] eu0/reg2_idx[0] eu0/reg2_idx[1]
+ eu0/reg2_idx[2] eu0/reg2_idx[3] eu0/reg2_idx[4] eu0/reg2_idx[5] eu0/reg2_val[0]
+ eu0/reg2_val[10] eu0/reg2_val[11] eu0/reg2_val[12] eu0/reg2_val[13] eu0/reg2_val[14]
+ eu0/reg2_val[15] eu0/reg2_val[16] eu0/reg2_val[17] eu0/reg2_val[18] eu0/reg2_val[19]
+ eu0/reg2_val[1] eu0/reg2_val[20] eu0/reg2_val[21] eu0/reg2_val[22] eu0/reg2_val[23]
+ eu0/reg2_val[24] eu0/reg2_val[25] eu0/reg2_val[26] eu0/reg2_val[27] eu0/reg2_val[28]
+ eu0/reg2_val[29] eu0/reg2_val[2] eu0/reg2_val[30] eu0/reg2_val[31] eu0/reg2_val[3]
+ eu0/reg2_val[4] eu0/reg2_val[5] eu0/reg2_val[6] eu0/reg2_val[7] eu0/reg2_val[8]
+ eu0/reg2_val[9] eu2/rst eu0/sign_extend eu0/take_branch vccd1 vssd1 wb_clk_i execution_unit
Xeu2 eu2/busy eu2/curr_PC[0] eu2/curr_PC[10] eu2/curr_PC[11] eu2/curr_PC[12] eu2/curr_PC[13]
+ eu2/curr_PC[14] eu2/curr_PC[15] eu2/curr_PC[16] eu2/curr_PC[17] eu2/curr_PC[18]
+ eu2/curr_PC[19] eu2/curr_PC[1] eu2/curr_PC[20] eu2/curr_PC[21] eu2/curr_PC[22] eu2/curr_PC[23]
+ eu2/curr_PC[24] eu2/curr_PC[25] eu2/curr_PC[26] eu2/curr_PC[27] eu2/curr_PC[2] eu2/curr_PC[3]
+ eu2/curr_PC[4] eu2/curr_PC[5] eu2/curr_PC[6] eu2/curr_PC[7] eu2/curr_PC[8] eu2/curr_PC[9]
+ eu2/dest_idx[0] eu2/dest_idx[1] eu2/dest_idx[2] eu2/dest_idx[3] eu2/dest_idx[4]
+ eu2/dest_idx[5] eu2/dest_mask[0] eu2/dest_mask[1] eu2/dest_pred[0] eu2/dest_pred[1]
+ eu2/dest_pred[2] eu2/dest_pred_val eu2/dest_val[0] eu2/dest_val[10] eu2/dest_val[11]
+ eu2/dest_val[12] eu2/dest_val[13] eu2/dest_val[14] eu2/dest_val[15] eu2/dest_val[16]
+ eu2/dest_val[17] eu2/dest_val[18] eu2/dest_val[19] eu2/dest_val[1] eu2/dest_val[20]
+ eu2/dest_val[21] eu2/dest_val[22] eu2/dest_val[23] eu2/dest_val[24] eu2/dest_val[25]
+ eu2/dest_val[26] eu2/dest_val[27] eu2/dest_val[28] eu2/dest_val[29] eu2/dest_val[2]
+ eu2/dest_val[30] eu2/dest_val[31] eu2/dest_val[3] eu2/dest_val[4] eu2/dest_val[5]
+ eu2/dest_val[6] eu2/dest_val[7] eu2/dest_val[8] eu2/dest_val[9] eu2/instruction[0]
+ eu2/instruction[10] eu2/instruction[11] eu2/instruction[12] eu2/instruction[13]
+ eu2/instruction[14] eu2/instruction[15] eu2/instruction[16] eu2/instruction[17]
+ eu2/instruction[18] eu2/instruction[19] eu2/instruction[1] eu2/instruction[20] eu2/instruction[21]
+ eu2/instruction[22] eu2/instruction[23] eu2/instruction[24] eu2/instruction[25]
+ eu2/instruction[26] eu2/instruction[27] eu2/instruction[28] eu2/instruction[29]
+ eu2/instruction[2] eu2/instruction[30] eu2/instruction[31] eu2/instruction[32] eu2/instruction[33]
+ eu2/instruction[34] eu2/instruction[35] eu2/instruction[36] eu2/instruction[37]
+ eu2/instruction[38] eu2/instruction[39] eu2/instruction[3] eu2/instruction[40] eu2/instruction[41]
+ eu2/instruction[4] eu2/instruction[5] eu2/instruction[6] eu2/instruction[7] eu2/instruction[8]
+ eu2/instruction[9] eu2/int_return eu2/is_load eu2/is_store eu2/loadstore_address[0]
+ eu2/loadstore_address[10] eu2/loadstore_address[11] eu2/loadstore_address[12] eu2/loadstore_address[13]
+ eu2/loadstore_address[14] eu2/loadstore_address[15] eu2/loadstore_address[16] eu2/loadstore_address[17]
+ eu2/loadstore_address[18] eu2/loadstore_address[19] eu2/loadstore_address[1] eu2/loadstore_address[20]
+ eu2/loadstore_address[21] eu2/loadstore_address[22] eu2/loadstore_address[23] eu2/loadstore_address[24]
+ eu2/loadstore_address[25] eu2/loadstore_address[26] eu2/loadstore_address[27] eu2/loadstore_address[28]
+ eu2/loadstore_address[29] eu2/loadstore_address[2] eu2/loadstore_address[30] eu2/loadstore_address[31]
+ eu2/loadstore_address[3] eu2/loadstore_address[4] eu2/loadstore_address[5] eu2/loadstore_address[6]
+ eu2/loadstore_address[7] eu2/loadstore_address[8] eu2/loadstore_address[9] eu2/loadstore_dest[0]
+ eu2/loadstore_dest[1] eu2/loadstore_dest[2] eu2/loadstore_dest[3] eu2/loadstore_dest[4]
+ eu2/loadstore_dest[5] eu2/loadstore_size[0] eu2/loadstore_size[1] eu2/new_PC[0]
+ eu2/new_PC[10] eu2/new_PC[11] eu2/new_PC[12] eu2/new_PC[13] eu2/new_PC[14] eu2/new_PC[15]
+ eu2/new_PC[16] eu2/new_PC[17] eu2/new_PC[18] eu2/new_PC[19] eu2/new_PC[1] eu2/new_PC[20]
+ eu2/new_PC[21] eu2/new_PC[22] eu2/new_PC[23] eu2/new_PC[24] eu2/new_PC[25] eu2/new_PC[26]
+ eu2/new_PC[27] eu2/new_PC[2] eu2/new_PC[3] eu2/new_PC[4] eu2/new_PC[5] eu2/new_PC[6]
+ eu2/new_PC[7] eu2/new_PC[8] eu2/new_PC[9] eu2/pred_idx[0] eu2/pred_idx[1] eu2/pred_idx[2]
+ eu2/pred_val eu2/reg1_idx[0] eu2/reg1_idx[1] eu2/reg1_idx[2] eu2/reg1_idx[3] eu2/reg1_idx[4]
+ eu2/reg1_idx[5] eu2/reg1_val[0] eu2/reg1_val[10] eu2/reg1_val[11] eu2/reg1_val[12]
+ eu2/reg1_val[13] eu2/reg1_val[14] eu2/reg1_val[15] eu2/reg1_val[16] eu2/reg1_val[17]
+ eu2/reg1_val[18] eu2/reg1_val[19] eu2/reg1_val[1] eu2/reg1_val[20] eu2/reg1_val[21]
+ eu2/reg1_val[22] eu2/reg1_val[23] eu2/reg1_val[24] eu2/reg1_val[25] eu2/reg1_val[26]
+ eu2/reg1_val[27] eu2/reg1_val[28] eu2/reg1_val[29] eu2/reg1_val[2] eu2/reg1_val[30]
+ eu2/reg1_val[31] eu2/reg1_val[3] eu2/reg1_val[4] eu2/reg1_val[5] eu2/reg1_val[6]
+ eu2/reg1_val[7] eu2/reg1_val[8] eu2/reg1_val[9] eu2/reg2_idx[0] eu2/reg2_idx[1]
+ eu2/reg2_idx[2] eu2/reg2_idx[3] eu2/reg2_idx[4] eu2/reg2_idx[5] eu2/reg2_val[0]
+ eu2/reg2_val[10] eu2/reg2_val[11] eu2/reg2_val[12] eu2/reg2_val[13] eu2/reg2_val[14]
+ eu2/reg2_val[15] eu2/reg2_val[16] eu2/reg2_val[17] eu2/reg2_val[18] eu2/reg2_val[19]
+ eu2/reg2_val[1] eu2/reg2_val[20] eu2/reg2_val[21] eu2/reg2_val[22] eu2/reg2_val[23]
+ eu2/reg2_val[24] eu2/reg2_val[25] eu2/reg2_val[26] eu2/reg2_val[27] eu2/reg2_val[28]
+ eu2/reg2_val[29] eu2/reg2_val[2] eu2/reg2_val[30] eu2/reg2_val[31] eu2/reg2_val[3]
+ eu2/reg2_val[4] eu2/reg2_val[5] eu2/reg2_val[6] eu2/reg2_val[7] eu2/reg2_val[8]
+ eu2/reg2_val[9] eu2/rst eu2/sign_extend eu2/take_branch vccd1 vssd1 wb_clk_i execution_unit
Xicache vliw/cache_entry[0] vliw/cache_entry[100] vliw/cache_entry[101] vliw/cache_entry[102]
+ vliw/cache_entry[103] vliw/cache_entry[104] vliw/cache_entry[105] vliw/cache_entry[106]
+ vliw/cache_entry[107] vliw/cache_entry[108] vliw/cache_entry[109] vliw/cache_entry[10]
+ vliw/cache_entry[110] vliw/cache_entry[111] vliw/cache_entry[112] vliw/cache_entry[113]
+ vliw/cache_entry[114] vliw/cache_entry[115] vliw/cache_entry[116] vliw/cache_entry[117]
+ vliw/cache_entry[118] vliw/cache_entry[119] vliw/cache_entry[11] vliw/cache_entry[120]
+ vliw/cache_entry[121] vliw/cache_entry[122] vliw/cache_entry[123] vliw/cache_entry[124]
+ vliw/cache_entry[125] vliw/cache_entry[126] vliw/cache_entry[127] vliw/cache_entry[12]
+ vliw/cache_entry[13] vliw/cache_entry[14] vliw/cache_entry[15] vliw/cache_entry[16]
+ vliw/cache_entry[17] vliw/cache_entry[18] vliw/cache_entry[19] vliw/cache_entry[1]
+ vliw/cache_entry[20] vliw/cache_entry[21] vliw/cache_entry[22] vliw/cache_entry[23]
+ vliw/cache_entry[24] vliw/cache_entry[25] vliw/cache_entry[26] vliw/cache_entry[27]
+ vliw/cache_entry[28] vliw/cache_entry[29] vliw/cache_entry[2] vliw/cache_entry[30]
+ vliw/cache_entry[31] vliw/cache_entry[32] vliw/cache_entry[33] vliw/cache_entry[34]
+ vliw/cache_entry[35] vliw/cache_entry[36] vliw/cache_entry[37] vliw/cache_entry[38]
+ vliw/cache_entry[39] vliw/cache_entry[3] vliw/cache_entry[40] vliw/cache_entry[41]
+ vliw/cache_entry[42] vliw/cache_entry[43] vliw/cache_entry[44] vliw/cache_entry[45]
+ vliw/cache_entry[46] vliw/cache_entry[47] vliw/cache_entry[48] vliw/cache_entry[49]
+ vliw/cache_entry[4] vliw/cache_entry[50] vliw/cache_entry[51] vliw/cache_entry[52]
+ vliw/cache_entry[53] vliw/cache_entry[54] vliw/cache_entry[55] vliw/cache_entry[56]
+ vliw/cache_entry[57] vliw/cache_entry[58] vliw/cache_entry[59] vliw/cache_entry[5]
+ vliw/cache_entry[60] vliw/cache_entry[61] vliw/cache_entry[62] vliw/cache_entry[63]
+ vliw/cache_entry[64] vliw/cache_entry[65] vliw/cache_entry[66] vliw/cache_entry[67]
+ vliw/cache_entry[68] vliw/cache_entry[69] vliw/cache_entry[6] vliw/cache_entry[70]
+ vliw/cache_entry[71] vliw/cache_entry[72] vliw/cache_entry[73] vliw/cache_entry[74]
+ vliw/cache_entry[75] vliw/cache_entry[76] vliw/cache_entry[77] vliw/cache_entry[78]
+ vliw/cache_entry[79] vliw/cache_entry[7] vliw/cache_entry[80] vliw/cache_entry[81]
+ vliw/cache_entry[82] vliw/cache_entry[83] vliw/cache_entry[84] vliw/cache_entry[85]
+ vliw/cache_entry[86] vliw/cache_entry[87] vliw/cache_entry[88] vliw/cache_entry[89]
+ vliw/cache_entry[8] vliw/cache_entry[90] vliw/cache_entry[91] vliw/cache_entry[92]
+ vliw/cache_entry[93] vliw/cache_entry[94] vliw/cache_entry[95] vliw/cache_entry[96]
+ vliw/cache_entry[97] vliw/cache_entry[98] vliw/cache_entry[99] vliw/cache_entry[9]
+ vliw/cache_hit vliw/cache_PC[0] vliw/cache_PC[10] vliw/cache_PC[11] vliw/cache_PC[12]
+ vliw/cache_PC[13] vliw/cache_PC[14] vliw/cache_PC[15] vliw/cache_PC[16] vliw/cache_PC[17]
+ vliw/cache_PC[18] vliw/cache_PC[19] vliw/cache_PC[1] vliw/cache_PC[20] vliw/cache_PC[21]
+ vliw/cache_PC[22] vliw/cache_PC[23] vliw/cache_PC[24] vliw/cache_PC[25] vliw/cache_PC[26]
+ vliw/cache_PC[27] vliw/cache_PC[2] vliw/cache_PC[3] vliw/cache_PC[4] vliw/cache_PC[5]
+ vliw/cache_PC[6] vliw/cache_PC[7] vliw/cache_PC[8] vliw/cache_PC[9] icache/entry_valid
+ icache/invalidate icache/new_entry[0] icache/new_entry[100] icache/new_entry[101]
+ icache/new_entry[102] icache/new_entry[103] icache/new_entry[104] icache/new_entry[105]
+ icache/new_entry[106] icache/new_entry[107] icache/new_entry[108] icache/new_entry[109]
+ icache/new_entry[10] icache/new_entry[110] icache/new_entry[111] icache/new_entry[112]
+ icache/new_entry[113] icache/new_entry[114] icache/new_entry[115] icache/new_entry[116]
+ icache/new_entry[117] icache/new_entry[118] icache/new_entry[119] icache/new_entry[11]
+ icache/new_entry[120] icache/new_entry[121] icache/new_entry[122] icache/new_entry[123]
+ icache/new_entry[124] icache/new_entry[125] icache/new_entry[126] icache/new_entry[127]
+ icache/new_entry[12] icache/new_entry[13] icache/new_entry[14] icache/new_entry[15]
+ icache/new_entry[16] icache/new_entry[17] icache/new_entry[18] icache/new_entry[19]
+ icache/new_entry[1] icache/new_entry[20] icache/new_entry[21] icache/new_entry[22]
+ icache/new_entry[23] icache/new_entry[24] icache/new_entry[25] icache/new_entry[26]
+ icache/new_entry[27] icache/new_entry[28] icache/new_entry[29] icache/new_entry[2]
+ icache/new_entry[30] icache/new_entry[31] icache/new_entry[32] icache/new_entry[33]
+ icache/new_entry[34] icache/new_entry[35] icache/new_entry[36] icache/new_entry[37]
+ icache/new_entry[38] icache/new_entry[39] icache/new_entry[3] icache/new_entry[40]
+ icache/new_entry[41] icache/new_entry[42] icache/new_entry[43] icache/new_entry[44]
+ icache/new_entry[45] icache/new_entry[46] icache/new_entry[47] icache/new_entry[48]
+ icache/new_entry[49] icache/new_entry[4] icache/new_entry[50] icache/new_entry[51]
+ icache/new_entry[52] icache/new_entry[53] icache/new_entry[54] icache/new_entry[55]
+ icache/new_entry[56] icache/new_entry[57] icache/new_entry[58] icache/new_entry[59]
+ icache/new_entry[5] icache/new_entry[60] icache/new_entry[61] icache/new_entry[62]
+ icache/new_entry[63] icache/new_entry[64] icache/new_entry[65] icache/new_entry[66]
+ icache/new_entry[67] icache/new_entry[68] icache/new_entry[69] icache/new_entry[6]
+ icache/new_entry[70] icache/new_entry[71] icache/new_entry[72] icache/new_entry[73]
+ icache/new_entry[74] icache/new_entry[75] icache/new_entry[76] icache/new_entry[77]
+ icache/new_entry[78] icache/new_entry[79] icache/new_entry[7] icache/new_entry[80]
+ icache/new_entry[81] icache/new_entry[82] icache/new_entry[83] icache/new_entry[84]
+ icache/new_entry[85] icache/new_entry[86] icache/new_entry[87] icache/new_entry[88]
+ icache/new_entry[89] icache/new_entry[8] icache/new_entry[90] icache/new_entry[91]
+ icache/new_entry[92] icache/new_entry[93] icache/new_entry[94] icache/new_entry[95]
+ icache/new_entry[96] icache/new_entry[97] icache/new_entry[98] icache/new_entry[99]
+ icache/new_entry[9] icache/rst vccd1 vssd1 wb_clk_i icache
Xwrapped_8x305 vliw/custom_settings[0] vliw/custom_settings[1] io_in[1] io_in[12]
+ io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20]
+ io_in[21] io_in[2] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28]
+ io_in[29] io_in[30] io_in[31] io_in[4] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36]
+ io_in[37] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] io_in[11] wrapped_8x305/io_oeb[0]
+ wrapped_8x305/io_oeb[1] wrapped_8x305/io_oeb[2] wrapped_8x305/io_oeb[3] wrapped_8x305/io_oeb[4]
+ wrapped_8x305/io_out[0] wrapped_8x305/io_out[10] wrapped_8x305/io_out[11] wrapped_8x305/io_out[12]
+ wrapped_8x305/io_out[13] wrapped_8x305/io_out[14] wrapped_8x305/io_out[15] wrapped_8x305/io_out[16]
+ wrapped_8x305/io_out[17] wrapped_8x305/io_out[18] wrapped_8x305/io_out[19] wrapped_8x305/io_out[1]
+ wrapped_8x305/io_out[20] wrapped_8x305/io_out[21] wrapped_8x305/io_out[22] wrapped_8x305/io_out[23]
+ wrapped_8x305/io_out[24] wrapped_8x305/io_out[25] wrapped_8x305/io_out[26] wrapped_8x305/io_out[27]
+ wrapped_8x305/io_out[28] wrapped_8x305/io_out[29] wrapped_8x305/io_out[2] wrapped_8x305/io_out[30]
+ wrapped_8x305/io_out[31] wrapped_8x305/io_out[32] wrapped_8x305/io_out[33] wrapped_8x305/io_out[34]
+ wrapped_8x305/io_out[35] wrapped_8x305/io_out[3] wrapped_8x305/io_out[4] wrapped_8x305/io_out[5]
+ wrapped_8x305/io_out[6] wrapped_8x305/io_out[7] wrapped_8x305/io_out[8] wrapped_8x305/io_out[9]
+ wrapped_8x305/rst_n vccd1 vssd1 wb_clk_i wrapped_8x305
Xscrapcpu io_in[1] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] io_in[21] io_in[2] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[27] io_in[28] io_in[29] io_in[30] io_in[31] io_in[4] io_in[32] io_in[33] io_in[34]
+ io_in[35] io_in[36] io_in[37] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10]
+ io_in[11] scrapcpu/io_oeb[0] scrapcpu/io_oeb[10] scrapcpu/io_oeb[11] scrapcpu/io_oeb[12]
+ scrapcpu/io_oeb[13] scrapcpu/io_oeb[14] scrapcpu/io_oeb[15] scrapcpu/io_oeb[16]
+ scrapcpu/io_oeb[17] scrapcpu/io_oeb[18] scrapcpu/io_oeb[19] scrapcpu/io_oeb[1] scrapcpu/io_oeb[20]
+ scrapcpu/io_oeb[21] scrapcpu/io_oeb[22] scrapcpu/io_oeb[23] scrapcpu/io_oeb[24]
+ scrapcpu/io_oeb[25] scrapcpu/io_oeb[26] scrapcpu/io_oeb[27] scrapcpu/io_oeb[28]
+ scrapcpu/io_oeb[29] scrapcpu/io_oeb[2] scrapcpu/io_oeb[30] scrapcpu/io_oeb[31] scrapcpu/io_oeb[32]
+ scrapcpu/io_oeb[33] scrapcpu/io_oeb[34] scrapcpu/io_oeb[35] scrapcpu/io_oeb[3] scrapcpu/io_oeb[4]
+ scrapcpu/io_oeb[5] scrapcpu/io_oeb[6] scrapcpu/io_oeb[7] scrapcpu/io_oeb[8] scrapcpu/io_oeb[9]
+ scrapcpu/io_out[0] scrapcpu/io_out[10] scrapcpu/io_out[11] scrapcpu/io_out[12] scrapcpu/io_out[13]
+ scrapcpu/io_out[14] scrapcpu/io_out[15] scrapcpu/io_out[16] scrapcpu/io_out[17]
+ scrapcpu/io_out[18] scrapcpu/io_out[19] scrapcpu/io_out[1] scrapcpu/io_out[20] scrapcpu/io_out[21]
+ scrapcpu/io_out[22] scrapcpu/io_out[23] scrapcpu/io_out[24] scrapcpu/io_out[25]
+ scrapcpu/io_out[26] scrapcpu/io_out[27] scrapcpu/io_out[28] scrapcpu/io_out[29]
+ scrapcpu/io_out[2] scrapcpu/io_out[30] scrapcpu/io_out[31] scrapcpu/io_out[32] scrapcpu/io_out[33]
+ scrapcpu/io_out[34] scrapcpu/io_out[35] scrapcpu/io_out[3] scrapcpu/io_out[4] scrapcpu/io_out[5]
+ scrapcpu/io_out[6] scrapcpu/io_out[7] scrapcpu/io_out[8] scrapcpu/io_out[9] scrapcpu/rst_n
+ vccd1 vssd1 wb_clk_i scrapcpu
Xmultiplexer multiplexer/cap_addr[0] multiplexer/cap_addr[1] multiplexer/cap_addr[2]
+ multiplexer/cap_addr[3] multiplexer/cap_addr[4] multiplexer/cap_addr[5] multiplexer/cap_addr[6]
+ multiplexer/cap_addr[7] multiplexer/cap_addr[8] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] vliw/custom_settings[0] multiplexer/custom_settings[10]
+ multiplexer/custom_settings[11] multiplexer/custom_settings[12] multiplexer/custom_settings[13]
+ multiplexer/custom_settings[14] multiplexer/custom_settings[15] multiplexer/custom_settings[16]
+ multiplexer/custom_settings[17] multiplexer/custom_settings[18] multiplexer/custom_settings[19]
+ vliw/custom_settings[1] multiplexer/custom_settings[20] multiplexer/custom_settings[21]
+ multiplexer/custom_settings[22] multiplexer/custom_settings[23] multiplexer/custom_settings[24]
+ multiplexer/custom_settings[25] multiplexer/custom_settings[26] multiplexer/custom_settings[27]
+ multiplexer/custom_settings[28] multiplexer/custom_settings[29] vliw/custom_settings[2]
+ multiplexer/custom_settings[30] multiplexer/custom_settings[31] vliw/custom_settings[3]
+ vliw/custom_settings[4] multiplexer/custom_settings[5] multiplexer/custom_settings[6]
+ multiplexer/custom_settings[7] multiplexer/custom_settings[8] multiplexer/custom_settings[9]
+ io_in[0] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2]
+ io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37]
+ io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] wrapped_6502/io_oeb
+ wrapped_8x305/io_oeb[0] wrapped_8x305/io_oeb[1] wrapped_8x305/io_oeb[2] wrapped_8x305/io_oeb[3]
+ wrapped_8x305/io_oeb[4] wrapped_as1802/io_oeb scrapcpu/io_oeb[0] scrapcpu/io_oeb[10]
+ scrapcpu/io_oeb[11] scrapcpu/io_oeb[12] scrapcpu/io_oeb[13] scrapcpu/io_oeb[14]
+ scrapcpu/io_oeb[15] scrapcpu/io_oeb[16] scrapcpu/io_oeb[17] scrapcpu/io_oeb[18]
+ scrapcpu/io_oeb[19] scrapcpu/io_oeb[1] scrapcpu/io_oeb[20] scrapcpu/io_oeb[21] scrapcpu/io_oeb[22]
+ scrapcpu/io_oeb[23] scrapcpu/io_oeb[24] scrapcpu/io_oeb[25] scrapcpu/io_oeb[26]
+ scrapcpu/io_oeb[27] scrapcpu/io_oeb[28] scrapcpu/io_oeb[29] scrapcpu/io_oeb[2] scrapcpu/io_oeb[30]
+ scrapcpu/io_oeb[31] scrapcpu/io_oeb[32] scrapcpu/io_oeb[33] scrapcpu/io_oeb[34]
+ scrapcpu/io_oeb[35] scrapcpu/io_oeb[3] scrapcpu/io_oeb[4] scrapcpu/io_oeb[5] scrapcpu/io_oeb[6]
+ scrapcpu/io_oeb[7] scrapcpu/io_oeb[8] scrapcpu/io_oeb[9] vliw/io_oeb[0] vliw/io_oeb[10]
+ vliw/io_oeb[11] vliw/io_oeb[12] vliw/io_oeb[13] vliw/io_oeb[14] vliw/io_oeb[15]
+ vliw/io_oeb[16] vliw/io_oeb[17] vliw/io_oeb[18] vliw/io_oeb[19] vliw/io_oeb[1] vliw/io_oeb[20]
+ vliw/io_oeb[21] vliw/io_oeb[22] vliw/io_oeb[23] vliw/io_oeb[24] vliw/io_oeb[25]
+ vliw/io_oeb[26] vliw/io_oeb[27] vliw/io_oeb[28] vliw/io_oeb[29] vliw/io_oeb[2] vliw/io_oeb[30]
+ vliw/io_oeb[31] vliw/io_oeb[32] vliw/io_oeb[33] vliw/io_oeb[34] vliw/io_oeb[35]
+ vliw/io_oeb[3] vliw/io_oeb[4] vliw/io_oeb[5] vliw/io_oeb[6] vliw/io_oeb[7] vliw/io_oeb[8]
+ vliw/io_oeb[9] ci2406_z80/io_oeb[0] ci2406_z80/io_oeb[10] ci2406_z80/io_oeb[11]
+ ci2406_z80/io_oeb[12] ci2406_z80/io_oeb[13] ci2406_z80/io_oeb[14] ci2406_z80/io_oeb[15]
+ ci2406_z80/io_oeb[16] ci2406_z80/io_oeb[17] ci2406_z80/io_oeb[18] ci2406_z80/io_oeb[19]
+ ci2406_z80/io_oeb[1] ci2406_z80/io_oeb[20] ci2406_z80/io_oeb[21] ci2406_z80/io_oeb[22]
+ ci2406_z80/io_oeb[23] ci2406_z80/io_oeb[24] ci2406_z80/io_oeb[25] ci2406_z80/io_oeb[26]
+ ci2406_z80/io_oeb[27] ci2406_z80/io_oeb[28] ci2406_z80/io_oeb[29] ci2406_z80/io_oeb[2]
+ ci2406_z80/io_oeb[30] ci2406_z80/io_oeb[31] ci2406_z80/io_oeb[32] ci2406_z80/io_oeb[33]
+ ci2406_z80/io_oeb[34] ci2406_z80/io_oeb[35] ci2406_z80/io_oeb[3] ci2406_z80/io_oeb[4]
+ ci2406_z80/io_oeb[5] ci2406_z80/io_oeb[6] ci2406_z80/io_oeb[7] ci2406_z80/io_oeb[8]
+ ci2406_z80/io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ wrapped_6502/io_out[0] wrapped_6502/io_out[10] wrapped_6502/io_out[11] wrapped_6502/io_out[12]
+ wrapped_6502/io_out[13] wrapped_6502/io_out[14] wrapped_6502/io_out[15] wrapped_6502/io_out[16]
+ wrapped_6502/io_out[17] wrapped_6502/io_out[18] wrapped_6502/io_out[19] wrapped_6502/io_out[1]
+ wrapped_6502/io_out[20] wrapped_6502/io_out[21] wrapped_6502/io_out[22] wrapped_6502/io_out[23]
+ wrapped_6502/io_out[24] wrapped_6502/io_out[25] wrapped_6502/io_out[26] wrapped_6502/io_out[27]
+ wrapped_6502/io_out[28] wrapped_6502/io_out[29] wrapped_6502/io_out[2] wrapped_6502/io_out[30]
+ wrapped_6502/io_out[31] wrapped_6502/io_out[32] wrapped_6502/io_out[33] wrapped_6502/io_out[34]
+ wrapped_6502/io_out[35] wrapped_6502/io_out[3] wrapped_6502/io_out[4] wrapped_6502/io_out[5]
+ wrapped_6502/io_out[6] wrapped_6502/io_out[7] wrapped_6502/io_out[8] wrapped_6502/io_out[9]
+ wrapped_8x305/io_out[0] wrapped_8x305/io_out[10] wrapped_8x305/io_out[11] wrapped_8x305/io_out[12]
+ wrapped_8x305/io_out[13] wrapped_8x305/io_out[14] wrapped_8x305/io_out[15] wrapped_8x305/io_out[16]
+ wrapped_8x305/io_out[17] wrapped_8x305/io_out[18] wrapped_8x305/io_out[19] wrapped_8x305/io_out[1]
+ wrapped_8x305/io_out[20] wrapped_8x305/io_out[21] wrapped_8x305/io_out[22] wrapped_8x305/io_out[23]
+ wrapped_8x305/io_out[24] wrapped_8x305/io_out[25] wrapped_8x305/io_out[26] wrapped_8x305/io_out[27]
+ wrapped_8x305/io_out[28] wrapped_8x305/io_out[29] wrapped_8x305/io_out[2] wrapped_8x305/io_out[30]
+ wrapped_8x305/io_out[31] wrapped_8x305/io_out[32] wrapped_8x305/io_out[33] wrapped_8x305/io_out[34]
+ wrapped_8x305/io_out[35] wrapped_8x305/io_out[3] wrapped_8x305/io_out[4] wrapped_8x305/io_out[5]
+ wrapped_8x305/io_out[6] wrapped_8x305/io_out[7] wrapped_8x305/io_out[8] wrapped_8x305/io_out[9]
+ wrapped_as1802/io_out[0] wrapped_as1802/io_out[10] wrapped_as1802/io_out[11] wrapped_as1802/io_out[12]
+ wrapped_as1802/io_out[13] wrapped_as1802/io_out[14] wrapped_as1802/io_out[15] wrapped_as1802/io_out[16]
+ wrapped_as1802/io_out[17] wrapped_as1802/io_out[18] wrapped_as1802/io_out[19] wrapped_as1802/io_out[1]
+ wrapped_as1802/io_out[20] wrapped_as1802/io_out[21] wrapped_as1802/io_out[22] wrapped_as1802/io_out[23]
+ wrapped_as1802/io_out[24] wrapped_as1802/io_out[25] wrapped_as1802/io_out[26] wrapped_as1802/io_out[27]
+ wrapped_as1802/io_out[28] wrapped_as1802/io_out[29] wrapped_as1802/io_out[2] wrapped_as1802/io_out[30]
+ wrapped_as1802/io_out[31] wrapped_as1802/io_out[32] wrapped_as1802/io_out[33] wrapped_as1802/io_out[34]
+ wrapped_as1802/io_out[35] wrapped_as1802/io_out[3] wrapped_as1802/io_out[4] wrapped_as1802/io_out[5]
+ wrapped_as1802/io_out[6] wrapped_as1802/io_out[7] wrapped_as1802/io_out[8] wrapped_as1802/io_out[9]
+ scrapcpu/io_out[0] scrapcpu/io_out[10] scrapcpu/io_out[11] scrapcpu/io_out[12] scrapcpu/io_out[13]
+ scrapcpu/io_out[14] scrapcpu/io_out[15] scrapcpu/io_out[16] scrapcpu/io_out[17]
+ scrapcpu/io_out[18] scrapcpu/io_out[19] scrapcpu/io_out[1] scrapcpu/io_out[20] scrapcpu/io_out[21]
+ scrapcpu/io_out[22] scrapcpu/io_out[23] scrapcpu/io_out[24] scrapcpu/io_out[25]
+ scrapcpu/io_out[26] scrapcpu/io_out[27] scrapcpu/io_out[28] scrapcpu/io_out[29]
+ scrapcpu/io_out[2] scrapcpu/io_out[30] scrapcpu/io_out[31] scrapcpu/io_out[32] scrapcpu/io_out[33]
+ scrapcpu/io_out[34] scrapcpu/io_out[35] scrapcpu/io_out[3] scrapcpu/io_out[4] scrapcpu/io_out[5]
+ scrapcpu/io_out[6] scrapcpu/io_out[7] scrapcpu/io_out[8] scrapcpu/io_out[9] vliw/io_out[0]
+ vliw/io_out[10] vliw/io_out[11] vliw/io_out[12] vliw/io_out[13] vliw/io_out[14]
+ vliw/io_out[15] vliw/io_out[16] vliw/io_out[17] vliw/io_out[18] vliw/io_out[19]
+ vliw/io_out[1] vliw/io_out[20] vliw/io_out[21] vliw/io_out[22] vliw/io_out[23] vliw/io_out[24]
+ vliw/io_out[25] vliw/io_out[26] vliw/io_out[27] vliw/io_out[28] vliw/io_out[29]
+ vliw/io_out[2] vliw/io_out[30] vliw/io_out[31] vliw/io_out[32] vliw/io_out[33] vliw/io_out[34]
+ vliw/io_out[35] vliw/io_out[3] vliw/io_out[4] vliw/io_out[5] vliw/io_out[6] vliw/io_out[7]
+ vliw/io_out[8] vliw/io_out[9] ci2406_z80/io_out[0] ci2406_z80/io_out[10] ci2406_z80/io_out[11]
+ ci2406_z80/io_out[12] ci2406_z80/io_out[13] ci2406_z80/io_out[14] ci2406_z80/io_out[15]
+ ci2406_z80/io_out[16] ci2406_z80/io_out[17] ci2406_z80/io_out[18] ci2406_z80/io_out[19]
+ ci2406_z80/io_out[1] ci2406_z80/io_out[20] ci2406_z80/io_out[21] ci2406_z80/io_out[22]
+ ci2406_z80/io_out[23] ci2406_z80/io_out[24] ci2406_z80/io_out[25] ci2406_z80/io_out[26]
+ ci2406_z80/io_out[27] ci2406_z80/io_out[28] ci2406_z80/io_out[29] ci2406_z80/io_out[2]
+ ci2406_z80/io_out[30] ci2406_z80/io_out[31] ci2406_z80/io_out[32] ci2406_z80/io_out[33]
+ ci2406_z80/io_out[34] ci2406_z80/io_out[35] ci2406_z80/io_out[3] ci2406_z80/io_out[4]
+ ci2406_z80/io_out[5] ci2406_z80/io_out[6] ci2406_z80/io_out[7] ci2406_z80/io_out[8]
+ ci2406_z80/io_out[9] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] wrapped_6502/rst_n wrapped_8x305/rst_n
+ wrapped_as1802/rst_n scrapcpu/rst_n vliw/rst_n ci2406_z80/rst_n vccd1 vssd1 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i
+ wbs_we_i multiplexer
Xvliw vliw/cache_PC[0] vliw/cache_PC[10] vliw/cache_PC[11] vliw/cache_PC[12] vliw/cache_PC[13]
+ vliw/cache_PC[14] vliw/cache_PC[15] vliw/cache_PC[16] vliw/cache_PC[17] vliw/cache_PC[18]
+ vliw/cache_PC[19] vliw/cache_PC[1] vliw/cache_PC[20] vliw/cache_PC[21] vliw/cache_PC[22]
+ vliw/cache_PC[23] vliw/cache_PC[24] vliw/cache_PC[25] vliw/cache_PC[26] vliw/cache_PC[27]
+ vliw/cache_PC[2] vliw/cache_PC[3] vliw/cache_PC[4] vliw/cache_PC[5] vliw/cache_PC[6]
+ vliw/cache_PC[7] vliw/cache_PC[8] vliw/cache_PC[9] vliw/cache_entry[0] vliw/cache_entry[100]
+ vliw/cache_entry[101] vliw/cache_entry[102] vliw/cache_entry[103] vliw/cache_entry[104]
+ vliw/cache_entry[105] vliw/cache_entry[106] vliw/cache_entry[107] vliw/cache_entry[108]
+ vliw/cache_entry[109] vliw/cache_entry[10] vliw/cache_entry[110] vliw/cache_entry[111]
+ vliw/cache_entry[112] vliw/cache_entry[113] vliw/cache_entry[114] vliw/cache_entry[115]
+ vliw/cache_entry[116] vliw/cache_entry[117] vliw/cache_entry[118] vliw/cache_entry[119]
+ vliw/cache_entry[11] vliw/cache_entry[120] vliw/cache_entry[121] vliw/cache_entry[122]
+ vliw/cache_entry[123] vliw/cache_entry[124] vliw/cache_entry[125] vliw/cache_entry[126]
+ vliw/cache_entry[127] vliw/cache_entry[12] vliw/cache_entry[13] vliw/cache_entry[14]
+ vliw/cache_entry[15] vliw/cache_entry[16] vliw/cache_entry[17] vliw/cache_entry[18]
+ vliw/cache_entry[19] vliw/cache_entry[1] vliw/cache_entry[20] vliw/cache_entry[21]
+ vliw/cache_entry[22] vliw/cache_entry[23] vliw/cache_entry[24] vliw/cache_entry[25]
+ vliw/cache_entry[26] vliw/cache_entry[27] vliw/cache_entry[28] vliw/cache_entry[29]
+ vliw/cache_entry[2] vliw/cache_entry[30] vliw/cache_entry[31] vliw/cache_entry[32]
+ vliw/cache_entry[33] vliw/cache_entry[34] vliw/cache_entry[35] vliw/cache_entry[36]
+ vliw/cache_entry[37] vliw/cache_entry[38] vliw/cache_entry[39] vliw/cache_entry[3]
+ vliw/cache_entry[40] vliw/cache_entry[41] vliw/cache_entry[42] vliw/cache_entry[43]
+ vliw/cache_entry[44] vliw/cache_entry[45] vliw/cache_entry[46] vliw/cache_entry[47]
+ vliw/cache_entry[48] vliw/cache_entry[49] vliw/cache_entry[4] vliw/cache_entry[50]
+ vliw/cache_entry[51] vliw/cache_entry[52] vliw/cache_entry[53] vliw/cache_entry[54]
+ vliw/cache_entry[55] vliw/cache_entry[56] vliw/cache_entry[57] vliw/cache_entry[58]
+ vliw/cache_entry[59] vliw/cache_entry[5] vliw/cache_entry[60] vliw/cache_entry[61]
+ vliw/cache_entry[62] vliw/cache_entry[63] vliw/cache_entry[64] vliw/cache_entry[65]
+ vliw/cache_entry[66] vliw/cache_entry[67] vliw/cache_entry[68] vliw/cache_entry[69]
+ vliw/cache_entry[6] vliw/cache_entry[70] vliw/cache_entry[71] vliw/cache_entry[72]
+ vliw/cache_entry[73] vliw/cache_entry[74] vliw/cache_entry[75] vliw/cache_entry[76]
+ vliw/cache_entry[77] vliw/cache_entry[78] vliw/cache_entry[79] vliw/cache_entry[7]
+ vliw/cache_entry[80] vliw/cache_entry[81] vliw/cache_entry[82] vliw/cache_entry[83]
+ vliw/cache_entry[84] vliw/cache_entry[85] vliw/cache_entry[86] vliw/cache_entry[87]
+ vliw/cache_entry[88] vliw/cache_entry[89] vliw/cache_entry[8] vliw/cache_entry[90]
+ vliw/cache_entry[91] vliw/cache_entry[92] vliw/cache_entry[93] vliw/cache_entry[94]
+ vliw/cache_entry[95] vliw/cache_entry[96] vliw/cache_entry[97] vliw/cache_entry[98]
+ vliw/cache_entry[99] vliw/cache_entry[9] icache/entry_valid vliw/cache_hit icache/invalidate
+ icache/new_entry[0] icache/new_entry[100] icache/new_entry[101] icache/new_entry[102]
+ icache/new_entry[103] icache/new_entry[104] icache/new_entry[105] icache/new_entry[106]
+ icache/new_entry[107] icache/new_entry[108] icache/new_entry[109] icache/new_entry[10]
+ icache/new_entry[110] icache/new_entry[111] icache/new_entry[112] icache/new_entry[113]
+ icache/new_entry[114] icache/new_entry[115] icache/new_entry[116] icache/new_entry[117]
+ icache/new_entry[118] icache/new_entry[119] icache/new_entry[11] icache/new_entry[120]
+ icache/new_entry[121] icache/new_entry[122] icache/new_entry[123] icache/new_entry[124]
+ icache/new_entry[125] icache/new_entry[126] icache/new_entry[127] icache/new_entry[12]
+ icache/new_entry[13] icache/new_entry[14] icache/new_entry[15] icache/new_entry[16]
+ icache/new_entry[17] icache/new_entry[18] icache/new_entry[19] icache/new_entry[1]
+ icache/new_entry[20] icache/new_entry[21] icache/new_entry[22] icache/new_entry[23]
+ icache/new_entry[24] icache/new_entry[25] icache/new_entry[26] icache/new_entry[27]
+ icache/new_entry[28] icache/new_entry[29] icache/new_entry[2] icache/new_entry[30]
+ icache/new_entry[31] icache/new_entry[32] icache/new_entry[33] icache/new_entry[34]
+ icache/new_entry[35] icache/new_entry[36] icache/new_entry[37] icache/new_entry[38]
+ icache/new_entry[39] icache/new_entry[3] icache/new_entry[40] icache/new_entry[41]
+ icache/new_entry[42] icache/new_entry[43] icache/new_entry[44] icache/new_entry[45]
+ icache/new_entry[46] icache/new_entry[47] icache/new_entry[48] icache/new_entry[49]
+ icache/new_entry[4] icache/new_entry[50] icache/new_entry[51] icache/new_entry[52]
+ icache/new_entry[53] icache/new_entry[54] icache/new_entry[55] icache/new_entry[56]
+ icache/new_entry[57] icache/new_entry[58] icache/new_entry[59] icache/new_entry[5]
+ icache/new_entry[60] icache/new_entry[61] icache/new_entry[62] icache/new_entry[63]
+ icache/new_entry[64] icache/new_entry[65] icache/new_entry[66] icache/new_entry[67]
+ icache/new_entry[68] icache/new_entry[69] icache/new_entry[6] icache/new_entry[70]
+ icache/new_entry[71] icache/new_entry[72] icache/new_entry[73] icache/new_entry[74]
+ icache/new_entry[75] icache/new_entry[76] icache/new_entry[77] icache/new_entry[78]
+ icache/new_entry[79] icache/new_entry[7] icache/new_entry[80] icache/new_entry[81]
+ icache/new_entry[82] icache/new_entry[83] icache/new_entry[84] icache/new_entry[85]
+ icache/new_entry[86] icache/new_entry[87] icache/new_entry[88] icache/new_entry[89]
+ icache/new_entry[8] icache/new_entry[90] icache/new_entry[91] icache/new_entry[92]
+ icache/new_entry[93] icache/new_entry[94] icache/new_entry[95] icache/new_entry[96]
+ icache/new_entry[97] icache/new_entry[98] icache/new_entry[99] icache/new_entry[9]
+ icache/rst eu2/curr_PC[0] eu2/curr_PC[10] eu2/curr_PC[11] eu2/curr_PC[12] eu2/curr_PC[13]
+ eu2/curr_PC[14] eu2/curr_PC[15] eu2/curr_PC[16] eu2/curr_PC[17] eu2/curr_PC[18]
+ eu2/curr_PC[19] eu2/curr_PC[1] eu2/curr_PC[20] eu2/curr_PC[21] eu2/curr_PC[22] eu2/curr_PC[23]
+ eu2/curr_PC[24] eu2/curr_PC[25] eu2/curr_PC[26] eu2/curr_PC[27] eu2/curr_PC[2] eu2/curr_PC[3]
+ eu2/curr_PC[4] eu2/curr_PC[5] eu2/curr_PC[6] eu2/curr_PC[7] eu2/curr_PC[8] eu2/curr_PC[9]
+ vliw/custom_settings[0] vliw/custom_settings[1] vliw/custom_settings[2] vliw/custom_settings[3]
+ vliw/custom_settings[4] eu0/dest_idx[0] eu0/dest_idx[1] eu0/dest_idx[2] eu0/dest_idx[3]
+ eu0/dest_idx[4] eu0/dest_idx[5] eu1/dest_idx[0] eu1/dest_idx[1] eu1/dest_idx[2]
+ eu1/dest_idx[3] eu1/dest_idx[4] eu1/dest_idx[5] eu2/dest_idx[0] eu2/dest_idx[1]
+ eu2/dest_idx[2] eu2/dest_idx[3] eu2/dest_idx[4] eu2/dest_idx[5] eu0/dest_mask[0]
+ eu0/dest_mask[1] eu1/dest_mask[0] eu1/dest_mask[1] eu2/dest_mask[0] eu2/dest_mask[1]
+ eu0/dest_pred[0] eu0/dest_pred[1] eu0/dest_pred[2] eu1/dest_pred[0] eu1/dest_pred[1]
+ eu1/dest_pred[2] eu2/dest_pred[0] eu2/dest_pred[1] eu2/dest_pred[2] eu0/dest_pred_val
+ eu1/dest_pred_val eu2/dest_pred_val eu0/dest_val[0] eu0/dest_val[10] eu0/dest_val[11]
+ eu0/dest_val[12] eu0/dest_val[13] eu0/dest_val[14] eu0/dest_val[15] eu0/dest_val[16]
+ eu0/dest_val[17] eu0/dest_val[18] eu0/dest_val[19] eu0/dest_val[1] eu0/dest_val[20]
+ eu0/dest_val[21] eu0/dest_val[22] eu0/dest_val[23] eu0/dest_val[24] eu0/dest_val[25]
+ eu0/dest_val[26] eu0/dest_val[27] eu0/dest_val[28] eu0/dest_val[29] eu0/dest_val[2]
+ eu0/dest_val[30] eu0/dest_val[31] eu0/dest_val[3] eu0/dest_val[4] eu0/dest_val[5]
+ eu0/dest_val[6] eu0/dest_val[7] eu0/dest_val[8] eu0/dest_val[9] eu1/dest_val[0]
+ eu1/dest_val[10] eu1/dest_val[11] eu1/dest_val[12] eu1/dest_val[13] eu1/dest_val[14]
+ eu1/dest_val[15] eu1/dest_val[16] eu1/dest_val[17] eu1/dest_val[18] eu1/dest_val[19]
+ eu1/dest_val[1] eu1/dest_val[20] eu1/dest_val[21] eu1/dest_val[22] eu1/dest_val[23]
+ eu1/dest_val[24] eu1/dest_val[25] eu1/dest_val[26] eu1/dest_val[27] eu1/dest_val[28]
+ eu1/dest_val[29] eu1/dest_val[2] eu1/dest_val[30] eu1/dest_val[31] eu1/dest_val[3]
+ eu1/dest_val[4] eu1/dest_val[5] eu1/dest_val[6] eu1/dest_val[7] eu1/dest_val[8]
+ eu1/dest_val[9] eu2/dest_val[0] eu2/dest_val[10] eu2/dest_val[11] eu2/dest_val[12]
+ eu2/dest_val[13] eu2/dest_val[14] eu2/dest_val[15] eu2/dest_val[16] eu2/dest_val[17]
+ eu2/dest_val[18] eu2/dest_val[19] eu2/dest_val[1] eu2/dest_val[20] eu2/dest_val[21]
+ eu2/dest_val[22] eu2/dest_val[23] eu2/dest_val[24] eu2/dest_val[25] eu2/dest_val[26]
+ eu2/dest_val[27] eu2/dest_val[28] eu2/dest_val[29] eu2/dest_val[2] eu2/dest_val[30]
+ eu2/dest_val[31] eu2/dest_val[3] eu2/dest_val[4] eu2/dest_val[5] eu2/dest_val[6]
+ eu2/dest_val[7] eu2/dest_val[8] eu2/dest_val[9] eu0/busy eu0/instruction[0] eu0/instruction[10]
+ eu0/instruction[11] eu0/instruction[12] eu0/instruction[13] eu0/instruction[14]
+ eu0/instruction[15] eu0/instruction[16] eu0/instruction[17] eu0/instruction[18]
+ eu0/instruction[19] eu0/instruction[1] eu0/instruction[20] eu0/instruction[21] eu0/instruction[22]
+ eu0/instruction[23] eu0/instruction[24] eu0/instruction[25] eu0/instruction[26]
+ eu0/instruction[27] eu0/instruction[28] eu0/instruction[29] eu0/instruction[2] eu0/instruction[30]
+ eu0/instruction[31] eu0/instruction[32] eu0/instruction[33] eu0/instruction[34]
+ eu0/instruction[35] eu0/instruction[36] eu0/instruction[37] eu0/instruction[38]
+ eu0/instruction[39] eu0/instruction[3] eu0/instruction[40] eu0/instruction[41] eu0/instruction[4]
+ eu0/instruction[5] eu0/instruction[6] eu0/instruction[7] eu0/instruction[8] eu0/instruction[9]
+ eu1/busy eu1/instruction[0] eu1/instruction[10] eu1/instruction[11] eu1/instruction[12]
+ eu1/instruction[13] eu1/instruction[14] eu1/instruction[15] eu1/instruction[16]
+ eu1/instruction[17] eu1/instruction[18] eu1/instruction[19] eu1/instruction[1] eu1/instruction[20]
+ eu1/instruction[21] eu1/instruction[22] eu1/instruction[23] eu1/instruction[24]
+ eu1/instruction[25] eu1/instruction[26] eu1/instruction[27] eu1/instruction[28]
+ eu1/instruction[29] eu1/instruction[2] eu1/instruction[30] eu1/instruction[31] eu1/instruction[32]
+ eu1/instruction[33] eu1/instruction[34] eu1/instruction[35] eu1/instruction[36]
+ eu1/instruction[37] eu1/instruction[38] eu1/instruction[39] eu1/instruction[3] eu1/instruction[40]
+ eu1/instruction[41] eu1/instruction[4] eu1/instruction[5] eu1/instruction[6] eu1/instruction[7]
+ eu1/instruction[8] eu1/instruction[9] eu2/busy eu2/instruction[0] eu2/instruction[10]
+ eu2/instruction[11] eu2/instruction[12] eu2/instruction[13] eu2/instruction[14]
+ eu2/instruction[15] eu2/instruction[16] eu2/instruction[17] eu2/instruction[18]
+ eu2/instruction[19] eu2/instruction[1] eu2/instruction[20] eu2/instruction[21] eu2/instruction[22]
+ eu2/instruction[23] eu2/instruction[24] eu2/instruction[25] eu2/instruction[26]
+ eu2/instruction[27] eu2/instruction[28] eu2/instruction[29] eu2/instruction[2] eu2/instruction[30]
+ eu2/instruction[31] eu2/instruction[32] eu2/instruction[33] eu2/instruction[34]
+ eu2/instruction[35] eu2/instruction[36] eu2/instruction[37] eu2/instruction[38]
+ eu2/instruction[39] eu2/instruction[3] eu2/instruction[40] eu2/instruction[41] eu2/instruction[4]
+ eu2/instruction[5] eu2/instruction[6] eu2/instruction[7] eu2/instruction[8] eu2/instruction[9]
+ eu0/int_return eu1/int_return eu2/int_return io_in[1] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[2] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[30]
+ io_in[31] io_in[4] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] io_in[11] vliw/io_oeb[0] vliw/io_oeb[10]
+ vliw/io_oeb[11] vliw/io_oeb[12] vliw/io_oeb[13] vliw/io_oeb[14] vliw/io_oeb[15]
+ vliw/io_oeb[16] vliw/io_oeb[17] vliw/io_oeb[18] vliw/io_oeb[19] vliw/io_oeb[1] vliw/io_oeb[20]
+ vliw/io_oeb[21] vliw/io_oeb[22] vliw/io_oeb[23] vliw/io_oeb[24] vliw/io_oeb[25]
+ vliw/io_oeb[26] vliw/io_oeb[27] vliw/io_oeb[28] vliw/io_oeb[29] vliw/io_oeb[2] vliw/io_oeb[30]
+ vliw/io_oeb[31] vliw/io_oeb[32] vliw/io_oeb[33] vliw/io_oeb[34] vliw/io_oeb[35]
+ vliw/io_oeb[3] vliw/io_oeb[4] vliw/io_oeb[5] vliw/io_oeb[6] vliw/io_oeb[7] vliw/io_oeb[8]
+ vliw/io_oeb[9] vliw/io_out[0] vliw/io_out[10] vliw/io_out[11] vliw/io_out[12] vliw/io_out[13]
+ vliw/io_out[14] vliw/io_out[15] vliw/io_out[16] vliw/io_out[17] vliw/io_out[18]
+ vliw/io_out[19] vliw/io_out[1] vliw/io_out[20] vliw/io_out[21] vliw/io_out[22] vliw/io_out[23]
+ vliw/io_out[24] vliw/io_out[25] vliw/io_out[26] vliw/io_out[27] vliw/io_out[28]
+ vliw/io_out[29] vliw/io_out[2] vliw/io_out[30] vliw/io_out[31] vliw/io_out[32] vliw/io_out[33]
+ vliw/io_out[34] vliw/io_out[35] vliw/io_out[3] vliw/io_out[4] vliw/io_out[5] vliw/io_out[6]
+ vliw/io_out[7] vliw/io_out[8] vliw/io_out[9] eu0/is_load eu1/is_load eu2/is_load
+ eu0/is_store eu1/is_store eu2/is_store eu0/loadstore_address[0] eu0/loadstore_address[10]
+ eu0/loadstore_address[11] eu0/loadstore_address[12] eu0/loadstore_address[13] eu0/loadstore_address[14]
+ eu0/loadstore_address[15] eu0/loadstore_address[16] eu0/loadstore_address[17] eu0/loadstore_address[18]
+ eu0/loadstore_address[19] eu0/loadstore_address[1] eu0/loadstore_address[20] eu0/loadstore_address[21]
+ eu0/loadstore_address[22] eu0/loadstore_address[23] eu0/loadstore_address[24] eu0/loadstore_address[25]
+ eu0/loadstore_address[26] eu0/loadstore_address[27] eu0/loadstore_address[28] eu0/loadstore_address[29]
+ eu0/loadstore_address[2] eu0/loadstore_address[30] eu0/loadstore_address[31] eu0/loadstore_address[3]
+ eu0/loadstore_address[4] eu0/loadstore_address[5] eu0/loadstore_address[6] eu0/loadstore_address[7]
+ eu0/loadstore_address[8] eu0/loadstore_address[9] eu1/loadstore_address[0] eu1/loadstore_address[10]
+ eu1/loadstore_address[11] eu1/loadstore_address[12] eu1/loadstore_address[13] eu1/loadstore_address[14]
+ eu1/loadstore_address[15] eu1/loadstore_address[16] eu1/loadstore_address[17] eu1/loadstore_address[18]
+ eu1/loadstore_address[19] eu1/loadstore_address[1] eu1/loadstore_address[20] eu1/loadstore_address[21]
+ eu1/loadstore_address[22] eu1/loadstore_address[23] eu1/loadstore_address[24] eu1/loadstore_address[25]
+ eu1/loadstore_address[26] eu1/loadstore_address[27] eu1/loadstore_address[28] eu1/loadstore_address[29]
+ eu1/loadstore_address[2] eu1/loadstore_address[30] eu1/loadstore_address[31] eu1/loadstore_address[3]
+ eu1/loadstore_address[4] eu1/loadstore_address[5] eu1/loadstore_address[6] eu1/loadstore_address[7]
+ eu1/loadstore_address[8] eu1/loadstore_address[9] eu2/loadstore_address[0] eu2/loadstore_address[10]
+ eu2/loadstore_address[11] eu2/loadstore_address[12] eu2/loadstore_address[13] eu2/loadstore_address[14]
+ eu2/loadstore_address[15] eu2/loadstore_address[16] eu2/loadstore_address[17] eu2/loadstore_address[18]
+ eu2/loadstore_address[19] eu2/loadstore_address[1] eu2/loadstore_address[20] eu2/loadstore_address[21]
+ eu2/loadstore_address[22] eu2/loadstore_address[23] eu2/loadstore_address[24] eu2/loadstore_address[25]
+ eu2/loadstore_address[26] eu2/loadstore_address[27] eu2/loadstore_address[28] eu2/loadstore_address[29]
+ eu2/loadstore_address[2] eu2/loadstore_address[30] eu2/loadstore_address[31] eu2/loadstore_address[3]
+ eu2/loadstore_address[4] eu2/loadstore_address[5] eu2/loadstore_address[6] eu2/loadstore_address[7]
+ eu2/loadstore_address[8] eu2/loadstore_address[9] eu0/loadstore_dest[0] eu0/loadstore_dest[1]
+ eu0/loadstore_dest[2] eu0/loadstore_dest[3] eu0/loadstore_dest[4] eu0/loadstore_dest[5]
+ eu1/loadstore_dest[0] eu1/loadstore_dest[1] eu1/loadstore_dest[2] eu1/loadstore_dest[3]
+ eu1/loadstore_dest[4] eu1/loadstore_dest[5] eu2/loadstore_dest[0] eu2/loadstore_dest[1]
+ eu2/loadstore_dest[2] eu2/loadstore_dest[3] eu2/loadstore_dest[4] eu2/loadstore_dest[5]
+ eu0/loadstore_size[0] eu0/loadstore_size[1] eu1/loadstore_size[0] eu1/loadstore_size[1]
+ eu2/loadstore_size[0] eu2/loadstore_size[1] eu0/new_PC[0] eu0/new_PC[10] eu0/new_PC[11]
+ eu0/new_PC[12] eu0/new_PC[13] eu0/new_PC[14] eu0/new_PC[15] eu0/new_PC[16] eu0/new_PC[17]
+ eu0/new_PC[18] eu0/new_PC[19] eu0/new_PC[1] eu0/new_PC[20] eu0/new_PC[21] eu0/new_PC[22]
+ eu0/new_PC[23] eu0/new_PC[24] eu0/new_PC[25] eu0/new_PC[26] eu0/new_PC[27] eu0/new_PC[2]
+ eu0/new_PC[3] eu0/new_PC[4] eu0/new_PC[5] eu0/new_PC[6] eu0/new_PC[7] eu0/new_PC[8]
+ eu0/new_PC[9] eu1/new_PC[0] eu1/new_PC[10] eu1/new_PC[11] eu1/new_PC[12] eu1/new_PC[13]
+ eu1/new_PC[14] eu1/new_PC[15] eu1/new_PC[16] eu1/new_PC[17] eu1/new_PC[18] eu1/new_PC[19]
+ eu1/new_PC[1] eu1/new_PC[20] eu1/new_PC[21] eu1/new_PC[22] eu1/new_PC[23] eu1/new_PC[24]
+ eu1/new_PC[25] eu1/new_PC[26] eu1/new_PC[27] eu1/new_PC[2] eu1/new_PC[3] eu1/new_PC[4]
+ eu1/new_PC[5] eu1/new_PC[6] eu1/new_PC[7] eu1/new_PC[8] eu1/new_PC[9] eu2/new_PC[0]
+ eu2/new_PC[10] eu2/new_PC[11] eu2/new_PC[12] eu2/new_PC[13] eu2/new_PC[14] eu2/new_PC[15]
+ eu2/new_PC[16] eu2/new_PC[17] eu2/new_PC[18] eu2/new_PC[19] eu2/new_PC[1] eu2/new_PC[20]
+ eu2/new_PC[21] eu2/new_PC[22] eu2/new_PC[23] eu2/new_PC[24] eu2/new_PC[25] eu2/new_PC[26]
+ eu2/new_PC[27] eu2/new_PC[2] eu2/new_PC[3] eu2/new_PC[4] eu2/new_PC[5] eu2/new_PC[6]
+ eu2/new_PC[7] eu2/new_PC[8] eu2/new_PC[9] eu0/pred_idx[0] eu0/pred_idx[1] eu0/pred_idx[2]
+ eu1/pred_idx[0] eu1/pred_idx[1] eu1/pred_idx[2] eu2/pred_idx[0] eu2/pred_idx[1]
+ eu2/pred_idx[2] eu0/pred_val eu1/pred_val eu2/pred_val eu0/reg1_idx[0] eu0/reg1_idx[1]
+ eu0/reg1_idx[2] eu0/reg1_idx[3] eu0/reg1_idx[4] eu0/reg1_idx[5] eu1/reg1_idx[0]
+ eu1/reg1_idx[1] eu1/reg1_idx[2] eu1/reg1_idx[3] eu1/reg1_idx[4] eu1/reg1_idx[5]
+ eu2/reg1_idx[0] eu2/reg1_idx[1] eu2/reg1_idx[2] eu2/reg1_idx[3] eu2/reg1_idx[4]
+ eu2/reg1_idx[5] eu0/reg1_val[0] eu0/reg1_val[10] eu0/reg1_val[11] eu0/reg1_val[12]
+ eu0/reg1_val[13] eu0/reg1_val[14] eu0/reg1_val[15] eu0/reg1_val[16] eu0/reg1_val[17]
+ eu0/reg1_val[18] eu0/reg1_val[19] eu0/reg1_val[1] eu0/reg1_val[20] eu0/reg1_val[21]
+ eu0/reg1_val[22] eu0/reg1_val[23] eu0/reg1_val[24] eu0/reg1_val[25] eu0/reg1_val[26]
+ eu0/reg1_val[27] eu0/reg1_val[28] eu0/reg1_val[29] eu0/reg1_val[2] eu0/reg1_val[30]
+ eu0/reg1_val[31] eu0/reg1_val[3] eu0/reg1_val[4] eu0/reg1_val[5] eu0/reg1_val[6]
+ eu0/reg1_val[7] eu0/reg1_val[8] eu0/reg1_val[9] eu1/reg1_val[0] eu1/reg1_val[10]
+ eu1/reg1_val[11] eu1/reg1_val[12] eu1/reg1_val[13] eu1/reg1_val[14] eu1/reg1_val[15]
+ eu1/reg1_val[16] eu1/reg1_val[17] eu1/reg1_val[18] eu1/reg1_val[19] eu1/reg1_val[1]
+ eu1/reg1_val[20] eu1/reg1_val[21] eu1/reg1_val[22] eu1/reg1_val[23] eu1/reg1_val[24]
+ eu1/reg1_val[25] eu1/reg1_val[26] eu1/reg1_val[27] eu1/reg1_val[28] eu1/reg1_val[29]
+ eu1/reg1_val[2] eu1/reg1_val[30] eu1/reg1_val[31] eu1/reg1_val[3] eu1/reg1_val[4]
+ eu1/reg1_val[5] eu1/reg1_val[6] eu1/reg1_val[7] eu1/reg1_val[8] eu1/reg1_val[9]
+ eu2/reg1_val[0] eu2/reg1_val[10] eu2/reg1_val[11] eu2/reg1_val[12] eu2/reg1_val[13]
+ eu2/reg1_val[14] eu2/reg1_val[15] eu2/reg1_val[16] eu2/reg1_val[17] eu2/reg1_val[18]
+ eu2/reg1_val[19] eu2/reg1_val[1] eu2/reg1_val[20] eu2/reg1_val[21] eu2/reg1_val[22]
+ eu2/reg1_val[23] eu2/reg1_val[24] eu2/reg1_val[25] eu2/reg1_val[26] eu2/reg1_val[27]
+ eu2/reg1_val[28] eu2/reg1_val[29] eu2/reg1_val[2] eu2/reg1_val[30] eu2/reg1_val[31]
+ eu2/reg1_val[3] eu2/reg1_val[4] eu2/reg1_val[5] eu2/reg1_val[6] eu2/reg1_val[7]
+ eu2/reg1_val[8] eu2/reg1_val[9] eu0/reg2_idx[0] eu0/reg2_idx[1] eu0/reg2_idx[2]
+ eu0/reg2_idx[3] eu0/reg2_idx[4] eu0/reg2_idx[5] eu1/reg2_idx[0] eu1/reg2_idx[1]
+ eu1/reg2_idx[2] eu1/reg2_idx[3] eu1/reg2_idx[4] eu1/reg2_idx[5] eu2/reg2_idx[0]
+ eu2/reg2_idx[1] eu2/reg2_idx[2] eu2/reg2_idx[3] eu2/reg2_idx[4] eu2/reg2_idx[5]
+ eu0/reg2_val[0] eu0/reg2_val[10] eu0/reg2_val[11] eu0/reg2_val[12] eu0/reg2_val[13]
+ eu0/reg2_val[14] eu0/reg2_val[15] eu0/reg2_val[16] eu0/reg2_val[17] eu0/reg2_val[18]
+ eu0/reg2_val[19] eu0/reg2_val[1] eu0/reg2_val[20] eu0/reg2_val[21] eu0/reg2_val[22]
+ eu0/reg2_val[23] eu0/reg2_val[24] eu0/reg2_val[25] eu0/reg2_val[26] eu0/reg2_val[27]
+ eu0/reg2_val[28] eu0/reg2_val[29] eu0/reg2_val[2] eu0/reg2_val[30] eu0/reg2_val[31]
+ eu0/reg2_val[3] eu0/reg2_val[4] eu0/reg2_val[5] eu0/reg2_val[6] eu0/reg2_val[7]
+ eu0/reg2_val[8] eu0/reg2_val[9] eu1/reg2_val[0] eu1/reg2_val[10] eu1/reg2_val[11]
+ eu1/reg2_val[12] eu1/reg2_val[13] eu1/reg2_val[14] eu1/reg2_val[15] eu1/reg2_val[16]
+ eu1/reg2_val[17] eu1/reg2_val[18] eu1/reg2_val[19] eu1/reg2_val[1] eu1/reg2_val[20]
+ eu1/reg2_val[21] eu1/reg2_val[22] eu1/reg2_val[23] eu1/reg2_val[24] eu1/reg2_val[25]
+ eu1/reg2_val[26] eu1/reg2_val[27] eu1/reg2_val[28] eu1/reg2_val[29] eu1/reg2_val[2]
+ eu1/reg2_val[30] eu1/reg2_val[31] eu1/reg2_val[3] eu1/reg2_val[4] eu1/reg2_val[5]
+ eu1/reg2_val[6] eu1/reg2_val[7] eu1/reg2_val[8] eu1/reg2_val[9] eu2/reg2_val[0]
+ eu2/reg2_val[10] eu2/reg2_val[11] eu2/reg2_val[12] eu2/reg2_val[13] eu2/reg2_val[14]
+ eu2/reg2_val[15] eu2/reg2_val[16] eu2/reg2_val[17] eu2/reg2_val[18] eu2/reg2_val[19]
+ eu2/reg2_val[1] eu2/reg2_val[20] eu2/reg2_val[21] eu2/reg2_val[22] eu2/reg2_val[23]
+ eu2/reg2_val[24] eu2/reg2_val[25] eu2/reg2_val[26] eu2/reg2_val[27] eu2/reg2_val[28]
+ eu2/reg2_val[29] eu2/reg2_val[2] eu2/reg2_val[30] eu2/reg2_val[31] eu2/reg2_val[3]
+ eu2/reg2_val[4] eu2/reg2_val[5] eu2/reg2_val[6] eu2/reg2_val[7] eu2/reg2_val[8]
+ eu2/reg2_val[9] eu2/rst vliw/rst_n eu0/sign_extend eu1/sign_extend eu2/sign_extend
+ eu0/take_branch eu1/take_branch eu2/take_branch vccd1 vssd1 wb_clk_i vliw
Xwrapped_as1802 vliw/custom_settings[0] multiplexer/custom_settings[10] multiplexer/custom_settings[11]
+ multiplexer/custom_settings[12] multiplexer/custom_settings[13] multiplexer/custom_settings[14]
+ multiplexer/custom_settings[15] multiplexer/custom_settings[16] multiplexer/custom_settings[17]
+ multiplexer/custom_settings[18] multiplexer/custom_settings[19] vliw/custom_settings[1]
+ multiplexer/custom_settings[20] multiplexer/custom_settings[21] multiplexer/custom_settings[22]
+ multiplexer/custom_settings[23] multiplexer/custom_settings[24] multiplexer/custom_settings[25]
+ multiplexer/custom_settings[26] multiplexer/custom_settings[27] multiplexer/custom_settings[28]
+ multiplexer/custom_settings[29] vliw/custom_settings[2] vliw/custom_settings[3]
+ vliw/custom_settings[4] multiplexer/custom_settings[5] multiplexer/custom_settings[6]
+ multiplexer/custom_settings[7] multiplexer/custom_settings[8] multiplexer/custom_settings[9]
+ io_in[1] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[20] io_in[21] io_in[2] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[30] io_in[31] io_in[4] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[36] io_in[37] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] io_in[11]
+ wrapped_as1802/io_oeb wrapped_as1802/io_out[0] wrapped_as1802/io_out[10] wrapped_as1802/io_out[11]
+ wrapped_as1802/io_out[12] wrapped_as1802/io_out[13] wrapped_as1802/io_out[14] wrapped_as1802/io_out[15]
+ wrapped_as1802/io_out[16] wrapped_as1802/io_out[17] wrapped_as1802/io_out[18] wrapped_as1802/io_out[19]
+ wrapped_as1802/io_out[1] wrapped_as1802/io_out[20] wrapped_as1802/io_out[21] wrapped_as1802/io_out[22]
+ wrapped_as1802/io_out[23] wrapped_as1802/io_out[24] wrapped_as1802/io_out[25] wrapped_as1802/io_out[26]
+ wrapped_as1802/io_out[27] wrapped_as1802/io_out[28] wrapped_as1802/io_out[29] wrapped_as1802/io_out[2]
+ wrapped_as1802/io_out[30] wrapped_as1802/io_out[31] wrapped_as1802/io_out[32] wrapped_as1802/io_out[33]
+ wrapped_as1802/io_out[34] wrapped_as1802/io_out[35] wrapped_as1802/io_out[3] wrapped_as1802/io_out[4]
+ wrapped_as1802/io_out[5] wrapped_as1802/io_out[6] wrapped_as1802/io_out[7] wrapped_as1802/io_out[8]
+ wrapped_as1802/io_out[9] wrapped_as1802/rst_n vccd1 vssd1 wb_clk_i wrapped_as1802
Xwrapped_6502 vliw/custom_settings[0] vliw/custom_settings[1] io_in[1] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21]
+ io_in[2] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[30] io_in[31] io_in[4] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10] io_in[11] wrapped_6502/io_oeb
+ wrapped_6502/io_out[0] wrapped_6502/io_out[10] wrapped_6502/io_out[11] wrapped_6502/io_out[12]
+ wrapped_6502/io_out[13] wrapped_6502/io_out[14] wrapped_6502/io_out[15] wrapped_6502/io_out[16]
+ wrapped_6502/io_out[17] wrapped_6502/io_out[18] wrapped_6502/io_out[19] wrapped_6502/io_out[1]
+ wrapped_6502/io_out[20] wrapped_6502/io_out[21] wrapped_6502/io_out[22] wrapped_6502/io_out[23]
+ wrapped_6502/io_out[24] wrapped_6502/io_out[25] wrapped_6502/io_out[26] wrapped_6502/io_out[27]
+ wrapped_6502/io_out[28] wrapped_6502/io_out[29] wrapped_6502/io_out[2] wrapped_6502/io_out[30]
+ wrapped_6502/io_out[31] wrapped_6502/io_out[32] wrapped_6502/io_out[33] wrapped_6502/io_out[34]
+ wrapped_6502/io_out[35] wrapped_6502/io_out[3] wrapped_6502/io_out[4] wrapped_6502/io_out[5]
+ wrapped_6502/io_out[6] wrapped_6502/io_out[7] wrapped_6502/io_out[8] wrapped_6502/io_out[9]
+ wrapped_6502/rst_n vccd1 vssd1 wb_clk_i wrapped_6502
Xunused_tie user_irq[0] user_irq[1] user_irq[2] la_data_out[40] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[41] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65]
+ la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[42]
+ la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[43] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[44] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[45] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[46] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[47]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[48] la_data_out[49]
+ vccd1 vssd1 wb_clk_i wb_rst_i unused_tie
Xci2406_z80 io_in[1] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] io_in[21] io_in[2] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[27] io_in[28] io_in[29] io_in[30] io_in[31] io_in[4] io_in[32] io_in[33] io_in[34]
+ io_in[35] io_in[36] io_in[37] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in[10]
+ io_in[11] ci2406_z80/io_oeb[0] ci2406_z80/io_oeb[10] ci2406_z80/io_oeb[11] ci2406_z80/io_oeb[12]
+ ci2406_z80/io_oeb[13] ci2406_z80/io_oeb[14] ci2406_z80/io_oeb[15] ci2406_z80/io_oeb[16]
+ ci2406_z80/io_oeb[17] ci2406_z80/io_oeb[18] ci2406_z80/io_oeb[19] ci2406_z80/io_oeb[1]
+ ci2406_z80/io_oeb[20] ci2406_z80/io_oeb[21] ci2406_z80/io_oeb[22] ci2406_z80/io_oeb[23]
+ ci2406_z80/io_oeb[24] ci2406_z80/io_oeb[25] ci2406_z80/io_oeb[26] ci2406_z80/io_oeb[27]
+ ci2406_z80/io_oeb[28] ci2406_z80/io_oeb[29] ci2406_z80/io_oeb[2] ci2406_z80/io_oeb[30]
+ ci2406_z80/io_oeb[31] ci2406_z80/io_oeb[32] ci2406_z80/io_oeb[33] ci2406_z80/io_oeb[34]
+ ci2406_z80/io_oeb[35] ci2406_z80/io_oeb[3] ci2406_z80/io_oeb[4] ci2406_z80/io_oeb[5]
+ ci2406_z80/io_oeb[6] ci2406_z80/io_oeb[7] ci2406_z80/io_oeb[8] ci2406_z80/io_oeb[9]
+ ci2406_z80/io_out[0] ci2406_z80/io_out[10] ci2406_z80/io_out[11] ci2406_z80/io_out[12]
+ ci2406_z80/io_out[13] ci2406_z80/io_out[14] ci2406_z80/io_out[15] ci2406_z80/io_out[16]
+ ci2406_z80/io_out[17] ci2406_z80/io_out[18] ci2406_z80/io_out[19] ci2406_z80/io_out[1]
+ ci2406_z80/io_out[20] ci2406_z80/io_out[21] ci2406_z80/io_out[22] ci2406_z80/io_out[23]
+ ci2406_z80/io_out[24] ci2406_z80/io_out[25] ci2406_z80/io_out[26] ci2406_z80/io_out[27]
+ ci2406_z80/io_out[28] ci2406_z80/io_out[29] ci2406_z80/io_out[2] ci2406_z80/io_out[30]
+ ci2406_z80/io_out[31] ci2406_z80/io_out[32] ci2406_z80/io_out[33] ci2406_z80/io_out[34]
+ ci2406_z80/io_out[35] ci2406_z80/io_out[3] ci2406_z80/io_out[4] ci2406_z80/io_out[5]
+ ci2406_z80/io_out[6] ci2406_z80/io_out[7] ci2406_z80/io_out[8] ci2406_z80/io_out[9]
+ ci2406_z80/rst_n vccd1 vssd1 wb_clk_i ci2406_z80
.ends

