VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 500.000 ;
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END custom_settings[9]
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 7.450 496.000 7.730 500.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_oeb[9]
  PIN io_oeb_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END io_oeb_scrapcpu[0]
  PIN io_oeb_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_oeb_scrapcpu[10]
  PIN io_oeb_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END io_oeb_scrapcpu[11]
  PIN io_oeb_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END io_oeb_scrapcpu[12]
  PIN io_oeb_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END io_oeb_scrapcpu[13]
  PIN io_oeb_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END io_oeb_scrapcpu[14]
  PIN io_oeb_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END io_oeb_scrapcpu[15]
  PIN io_oeb_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END io_oeb_scrapcpu[16]
  PIN io_oeb_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END io_oeb_scrapcpu[17]
  PIN io_oeb_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_oeb_scrapcpu[18]
  PIN io_oeb_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END io_oeb_scrapcpu[19]
  PIN io_oeb_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END io_oeb_scrapcpu[1]
  PIN io_oeb_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END io_oeb_scrapcpu[20]
  PIN io_oeb_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_oeb_scrapcpu[21]
  PIN io_oeb_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END io_oeb_scrapcpu[22]
  PIN io_oeb_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END io_oeb_scrapcpu[23]
  PIN io_oeb_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_oeb_scrapcpu[24]
  PIN io_oeb_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END io_oeb_scrapcpu[25]
  PIN io_oeb_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END io_oeb_scrapcpu[26]
  PIN io_oeb_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END io_oeb_scrapcpu[27]
  PIN io_oeb_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END io_oeb_scrapcpu[28]
  PIN io_oeb_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_oeb_scrapcpu[29]
  PIN io_oeb_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_oeb_scrapcpu[2]
  PIN io_oeb_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END io_oeb_scrapcpu[30]
  PIN io_oeb_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END io_oeb_scrapcpu[31]
  PIN io_oeb_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END io_oeb_scrapcpu[32]
  PIN io_oeb_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END io_oeb_scrapcpu[33]
  PIN io_oeb_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END io_oeb_scrapcpu[34]
  PIN io_oeb_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END io_oeb_scrapcpu[35]
  PIN io_oeb_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END io_oeb_scrapcpu[3]
  PIN io_oeb_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END io_oeb_scrapcpu[4]
  PIN io_oeb_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END io_oeb_scrapcpu[5]
  PIN io_oeb_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END io_oeb_scrapcpu[6]
  PIN io_oeb_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END io_oeb_scrapcpu[7]
  PIN io_oeb_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END io_oeb_scrapcpu[8]
  PIN io_oeb_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END io_oeb_scrapcpu[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 496.000 17.850 500.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 118.770 496.000 119.050 500.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 496.000 129.170 500.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.010 496.000 139.290 500.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 149.130 496.000 149.410 500.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 496.000 159.530 500.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 496.000 169.650 500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 179.490 496.000 179.770 500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 189.610 496.000 189.890 500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 496.000 200.010 500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 496.000 210.130 500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 27.690 496.000 27.970 500.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.970 496.000 220.250 500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 230.090 496.000 230.370 500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 240.210 496.000 240.490 500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 250.330 496.000 250.610 500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 496.000 260.730 500.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 496.000 270.850 500.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 280.690 496.000 280.970 500.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 290.810 496.000 291.090 500.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 300.930 496.000 301.210 500.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 311.050 496.000 311.330 500.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 496.000 38.090 500.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 321.170 496.000 321.450 500.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 331.290 496.000 331.570 500.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 351.530 496.000 351.810 500.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 361.650 496.000 361.930 500.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 371.770 496.000 372.050 500.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 381.890 496.000 382.170 500.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.010 496.000 392.290 500.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.930 496.000 48.210 500.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 496.000 58.330 500.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 496.000 68.450 500.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 78.290 496.000 78.570 500.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 496.000 88.690 500.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 496.000 98.810 500.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 108.650 496.000 108.930 500.000 ;
    END
  END io_out[9]
  PIN io_out_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_out_scrapcpu[0]
  PIN io_out_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_out_scrapcpu[10]
  PIN io_out_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END io_out_scrapcpu[11]
  PIN io_out_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END io_out_scrapcpu[12]
  PIN io_out_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_out_scrapcpu[13]
  PIN io_out_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END io_out_scrapcpu[14]
  PIN io_out_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_out_scrapcpu[15]
  PIN io_out_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_out_scrapcpu[16]
  PIN io_out_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_out_scrapcpu[17]
  PIN io_out_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_out_scrapcpu[18]
  PIN io_out_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END io_out_scrapcpu[19]
  PIN io_out_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END io_out_scrapcpu[1]
  PIN io_out_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_out_scrapcpu[20]
  PIN io_out_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END io_out_scrapcpu[21]
  PIN io_out_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END io_out_scrapcpu[22]
  PIN io_out_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END io_out_scrapcpu[23]
  PIN io_out_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END io_out_scrapcpu[24]
  PIN io_out_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_out_scrapcpu[25]
  PIN io_out_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END io_out_scrapcpu[26]
  PIN io_out_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END io_out_scrapcpu[27]
  PIN io_out_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END io_out_scrapcpu[28]
  PIN io_out_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END io_out_scrapcpu[29]
  PIN io_out_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END io_out_scrapcpu[2]
  PIN io_out_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_out_scrapcpu[30]
  PIN io_out_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END io_out_scrapcpu[31]
  PIN io_out_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END io_out_scrapcpu[32]
  PIN io_out_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END io_out_scrapcpu[33]
  PIN io_out_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END io_out_scrapcpu[34]
  PIN io_out_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END io_out_scrapcpu[35]
  PIN io_out_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END io_out_scrapcpu[3]
  PIN io_out_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END io_out_scrapcpu[4]
  PIN io_out_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_out_scrapcpu[5]
  PIN io_out_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END io_out_scrapcpu[6]
  PIN io_out_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_out_scrapcpu[7]
  PIN io_out_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END io_out_scrapcpu[8]
  PIN io_out_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_out_scrapcpu[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.200 400.000 178.800 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.000 400.000 219.600 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.080 400.000 223.680 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.160 400.000 227.760 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.240 400.000 231.840 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 235.320 400.000 235.920 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 239.400 400.000 240.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 243.480 400.000 244.080 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 247.560 400.000 248.160 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.720 400.000 256.320 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.280 400.000 182.880 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.800 400.000 260.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.880 400.000 264.480 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.960 400.000 268.560 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.040 400.000 272.640 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.120 400.000 276.720 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.200 400.000 280.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.280 400.000 284.880 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 288.360 400.000 288.960 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 292.440 400.000 293.040 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 296.520 400.000 297.120 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 186.360 400.000 186.960 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 300.600 400.000 301.200 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.680 400.000 305.280 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.760 400.000 309.360 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.840 400.000 313.440 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.920 400.000 317.520 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.080 400.000 325.680 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.160 400.000 329.760 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.240 400.000 333.840 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 337.320 400.000 337.920 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 194.520 400.000 195.120 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 198.600 400.000 199.200 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.680 400.000 203.280 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.760 400.000 207.360 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.920 400.000 215.520 ;
    END
  END la_data_out[9]
  PIN rst_scrapcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END rst_scrapcpu
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 174.120 400.000 174.720 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.960 400.000 166.560 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 382.200 400.000 382.800 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 386.280 400.000 386.880 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 390.360 400.000 390.960 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 394.440 400.000 395.040 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 398.520 400.000 399.120 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 402.600 400.000 403.200 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 406.680 400.000 407.280 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 410.760 400.000 411.360 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 414.840 400.000 415.440 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 418.920 400.000 419.520 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 345.480 400.000 346.080 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 423.000 400.000 423.600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 427.080 400.000 427.680 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 431.160 400.000 431.760 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 435.240 400.000 435.840 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 439.320 400.000 439.920 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 443.400 400.000 444.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 447.480 400.000 448.080 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 451.560 400.000 452.160 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 455.640 400.000 456.240 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 459.720 400.000 460.320 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 349.560 400.000 350.160 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 463.800 400.000 464.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 467.880 400.000 468.480 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 353.640 400.000 354.240 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.720 400.000 358.320 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.800 400.000 362.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.880 400.000 366.480 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 369.960 400.000 370.560 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.040 400.000 374.640 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 378.120 400.000 378.720 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 31.320 400.000 31.920 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.280 400.000 80.880 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 84.360 400.000 84.960 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 92.520 400.000 93.120 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 96.600 400.000 97.200 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.680 400.000 101.280 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.760 400.000 105.360 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 35.400 400.000 36.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.920 400.000 113.520 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.000 400.000 117.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.080 400.000 121.680 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.160 400.000 125.760 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 133.320 400.000 133.920 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 137.400 400.000 138.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 141.480 400.000 142.080 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 145.560 400.000 146.160 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 39.480 400.000 40.080 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.720 400.000 154.320 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.800 400.000 158.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 43.560 400.000 44.160 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 47.640 400.000 48.240 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.720 400.000 52.320 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.800 400.000 56.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.880 400.000 60.480 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.960 400.000 64.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.880 400.000 162.480 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 486.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 395.530 487.120 ;
      LAYER met2 ;
        RECT 0.100 495.720 7.170 496.810 ;
        RECT 8.010 495.720 17.290 496.810 ;
        RECT 18.130 495.720 27.410 496.810 ;
        RECT 28.250 495.720 37.530 496.810 ;
        RECT 38.370 495.720 47.650 496.810 ;
        RECT 48.490 495.720 57.770 496.810 ;
        RECT 58.610 495.720 67.890 496.810 ;
        RECT 68.730 495.720 78.010 496.810 ;
        RECT 78.850 495.720 88.130 496.810 ;
        RECT 88.970 495.720 98.250 496.810 ;
        RECT 99.090 495.720 108.370 496.810 ;
        RECT 109.210 495.720 118.490 496.810 ;
        RECT 119.330 495.720 128.610 496.810 ;
        RECT 129.450 495.720 138.730 496.810 ;
        RECT 139.570 495.720 148.850 496.810 ;
        RECT 149.690 495.720 158.970 496.810 ;
        RECT 159.810 495.720 169.090 496.810 ;
        RECT 169.930 495.720 179.210 496.810 ;
        RECT 180.050 495.720 189.330 496.810 ;
        RECT 190.170 495.720 199.450 496.810 ;
        RECT 200.290 495.720 209.570 496.810 ;
        RECT 210.410 495.720 219.690 496.810 ;
        RECT 220.530 495.720 229.810 496.810 ;
        RECT 230.650 495.720 239.930 496.810 ;
        RECT 240.770 495.720 250.050 496.810 ;
        RECT 250.890 495.720 260.170 496.810 ;
        RECT 261.010 495.720 270.290 496.810 ;
        RECT 271.130 495.720 280.410 496.810 ;
        RECT 281.250 495.720 290.530 496.810 ;
        RECT 291.370 495.720 300.650 496.810 ;
        RECT 301.490 495.720 310.770 496.810 ;
        RECT 311.610 495.720 320.890 496.810 ;
        RECT 321.730 495.720 331.010 496.810 ;
        RECT 331.850 495.720 341.130 496.810 ;
        RECT 341.970 495.720 351.250 496.810 ;
        RECT 352.090 495.720 361.370 496.810 ;
        RECT 362.210 495.720 371.490 496.810 ;
        RECT 372.330 495.720 381.610 496.810 ;
        RECT 382.450 495.720 391.730 496.810 ;
        RECT 392.570 495.720 395.510 496.810 ;
        RECT 0.100 4.280 395.510 495.720 ;
        RECT 0.100 3.670 4.870 4.280 ;
        RECT 5.710 3.670 10.850 4.280 ;
        RECT 11.690 3.670 16.830 4.280 ;
        RECT 17.670 3.670 22.810 4.280 ;
        RECT 23.650 3.670 28.790 4.280 ;
        RECT 29.630 3.670 34.770 4.280 ;
        RECT 35.610 3.670 40.750 4.280 ;
        RECT 41.590 3.670 46.730 4.280 ;
        RECT 47.570 3.670 52.710 4.280 ;
        RECT 53.550 3.670 58.690 4.280 ;
        RECT 59.530 3.670 64.670 4.280 ;
        RECT 65.510 3.670 70.650 4.280 ;
        RECT 71.490 3.670 76.630 4.280 ;
        RECT 77.470 3.670 82.610 4.280 ;
        RECT 83.450 3.670 88.590 4.280 ;
        RECT 89.430 3.670 94.570 4.280 ;
        RECT 95.410 3.670 100.550 4.280 ;
        RECT 101.390 3.670 106.530 4.280 ;
        RECT 107.370 3.670 112.510 4.280 ;
        RECT 113.350 3.670 118.490 4.280 ;
        RECT 119.330 3.670 124.470 4.280 ;
        RECT 125.310 3.670 130.450 4.280 ;
        RECT 131.290 3.670 136.430 4.280 ;
        RECT 137.270 3.670 142.410 4.280 ;
        RECT 143.250 3.670 148.390 4.280 ;
        RECT 149.230 3.670 154.370 4.280 ;
        RECT 155.210 3.670 160.350 4.280 ;
        RECT 161.190 3.670 166.330 4.280 ;
        RECT 167.170 3.670 172.310 4.280 ;
        RECT 173.150 3.670 178.290 4.280 ;
        RECT 179.130 3.670 184.270 4.280 ;
        RECT 185.110 3.670 190.250 4.280 ;
        RECT 191.090 3.670 196.230 4.280 ;
        RECT 197.070 3.670 202.210 4.280 ;
        RECT 203.050 3.670 208.190 4.280 ;
        RECT 209.030 3.670 214.170 4.280 ;
        RECT 215.010 3.670 220.150 4.280 ;
        RECT 220.990 3.670 226.130 4.280 ;
        RECT 226.970 3.670 232.110 4.280 ;
        RECT 232.950 3.670 238.090 4.280 ;
        RECT 238.930 3.670 244.070 4.280 ;
        RECT 244.910 3.670 250.050 4.280 ;
        RECT 250.890 3.670 256.030 4.280 ;
        RECT 256.870 3.670 262.010 4.280 ;
        RECT 262.850 3.670 267.990 4.280 ;
        RECT 268.830 3.670 273.970 4.280 ;
        RECT 274.810 3.670 279.950 4.280 ;
        RECT 280.790 3.670 285.930 4.280 ;
        RECT 286.770 3.670 291.910 4.280 ;
        RECT 292.750 3.670 297.890 4.280 ;
        RECT 298.730 3.670 303.870 4.280 ;
        RECT 304.710 3.670 309.850 4.280 ;
        RECT 310.690 3.670 315.830 4.280 ;
        RECT 316.670 3.670 321.810 4.280 ;
        RECT 322.650 3.670 327.790 4.280 ;
        RECT 328.630 3.670 333.770 4.280 ;
        RECT 334.610 3.670 339.750 4.280 ;
        RECT 340.590 3.670 345.730 4.280 ;
        RECT 346.570 3.670 351.710 4.280 ;
        RECT 352.550 3.670 357.690 4.280 ;
        RECT 358.530 3.670 363.670 4.280 ;
        RECT 364.510 3.670 369.650 4.280 ;
        RECT 370.490 3.670 375.630 4.280 ;
        RECT 376.470 3.670 381.610 4.280 ;
        RECT 382.450 3.670 387.590 4.280 ;
        RECT 388.430 3.670 393.570 4.280 ;
        RECT 394.410 3.670 395.510 4.280 ;
      LAYER met3 ;
        RECT 3.990 474.320 396.000 487.045 ;
        RECT 4.400 472.920 396.000 474.320 ;
        RECT 3.990 470.240 396.000 472.920 ;
        RECT 4.400 468.880 396.000 470.240 ;
        RECT 4.400 468.840 395.600 468.880 ;
        RECT 3.990 467.480 395.600 468.840 ;
        RECT 3.990 466.160 396.000 467.480 ;
        RECT 4.400 464.800 396.000 466.160 ;
        RECT 4.400 464.760 395.600 464.800 ;
        RECT 3.990 463.400 395.600 464.760 ;
        RECT 3.990 462.080 396.000 463.400 ;
        RECT 4.400 460.720 396.000 462.080 ;
        RECT 4.400 460.680 395.600 460.720 ;
        RECT 3.990 459.320 395.600 460.680 ;
        RECT 3.990 458.000 396.000 459.320 ;
        RECT 4.400 456.640 396.000 458.000 ;
        RECT 4.400 456.600 395.600 456.640 ;
        RECT 3.990 455.240 395.600 456.600 ;
        RECT 3.990 453.920 396.000 455.240 ;
        RECT 4.400 452.560 396.000 453.920 ;
        RECT 4.400 452.520 395.600 452.560 ;
        RECT 3.990 451.160 395.600 452.520 ;
        RECT 3.990 449.840 396.000 451.160 ;
        RECT 4.400 448.480 396.000 449.840 ;
        RECT 4.400 448.440 395.600 448.480 ;
        RECT 3.990 447.080 395.600 448.440 ;
        RECT 3.990 445.760 396.000 447.080 ;
        RECT 4.400 444.400 396.000 445.760 ;
        RECT 4.400 444.360 395.600 444.400 ;
        RECT 3.990 443.000 395.600 444.360 ;
        RECT 3.990 441.680 396.000 443.000 ;
        RECT 4.400 440.320 396.000 441.680 ;
        RECT 4.400 440.280 395.600 440.320 ;
        RECT 3.990 438.920 395.600 440.280 ;
        RECT 3.990 437.600 396.000 438.920 ;
        RECT 4.400 436.240 396.000 437.600 ;
        RECT 4.400 436.200 395.600 436.240 ;
        RECT 3.990 434.840 395.600 436.200 ;
        RECT 3.990 433.520 396.000 434.840 ;
        RECT 4.400 432.160 396.000 433.520 ;
        RECT 4.400 432.120 395.600 432.160 ;
        RECT 3.990 430.760 395.600 432.120 ;
        RECT 3.990 429.440 396.000 430.760 ;
        RECT 4.400 428.080 396.000 429.440 ;
        RECT 4.400 428.040 395.600 428.080 ;
        RECT 3.990 426.680 395.600 428.040 ;
        RECT 3.990 425.360 396.000 426.680 ;
        RECT 4.400 424.000 396.000 425.360 ;
        RECT 4.400 423.960 395.600 424.000 ;
        RECT 3.990 422.600 395.600 423.960 ;
        RECT 3.990 421.280 396.000 422.600 ;
        RECT 4.400 419.920 396.000 421.280 ;
        RECT 4.400 419.880 395.600 419.920 ;
        RECT 3.990 418.520 395.600 419.880 ;
        RECT 3.990 417.200 396.000 418.520 ;
        RECT 4.400 415.840 396.000 417.200 ;
        RECT 4.400 415.800 395.600 415.840 ;
        RECT 3.990 414.440 395.600 415.800 ;
        RECT 3.990 413.120 396.000 414.440 ;
        RECT 4.400 411.760 396.000 413.120 ;
        RECT 4.400 411.720 395.600 411.760 ;
        RECT 3.990 410.360 395.600 411.720 ;
        RECT 3.990 409.040 396.000 410.360 ;
        RECT 4.400 407.680 396.000 409.040 ;
        RECT 4.400 407.640 395.600 407.680 ;
        RECT 3.990 406.280 395.600 407.640 ;
        RECT 3.990 404.960 396.000 406.280 ;
        RECT 4.400 403.600 396.000 404.960 ;
        RECT 4.400 403.560 395.600 403.600 ;
        RECT 3.990 402.200 395.600 403.560 ;
        RECT 3.990 400.880 396.000 402.200 ;
        RECT 4.400 399.520 396.000 400.880 ;
        RECT 4.400 399.480 395.600 399.520 ;
        RECT 3.990 398.120 395.600 399.480 ;
        RECT 3.990 396.800 396.000 398.120 ;
        RECT 4.400 395.440 396.000 396.800 ;
        RECT 4.400 395.400 395.600 395.440 ;
        RECT 3.990 394.040 395.600 395.400 ;
        RECT 3.990 392.720 396.000 394.040 ;
        RECT 4.400 391.360 396.000 392.720 ;
        RECT 4.400 391.320 395.600 391.360 ;
        RECT 3.990 389.960 395.600 391.320 ;
        RECT 3.990 388.640 396.000 389.960 ;
        RECT 4.400 387.280 396.000 388.640 ;
        RECT 4.400 387.240 395.600 387.280 ;
        RECT 3.990 385.880 395.600 387.240 ;
        RECT 3.990 384.560 396.000 385.880 ;
        RECT 4.400 383.200 396.000 384.560 ;
        RECT 4.400 383.160 395.600 383.200 ;
        RECT 3.990 381.800 395.600 383.160 ;
        RECT 3.990 380.480 396.000 381.800 ;
        RECT 4.400 379.120 396.000 380.480 ;
        RECT 4.400 379.080 395.600 379.120 ;
        RECT 3.990 377.720 395.600 379.080 ;
        RECT 3.990 376.400 396.000 377.720 ;
        RECT 4.400 375.040 396.000 376.400 ;
        RECT 4.400 375.000 395.600 375.040 ;
        RECT 3.990 373.640 395.600 375.000 ;
        RECT 3.990 372.320 396.000 373.640 ;
        RECT 4.400 370.960 396.000 372.320 ;
        RECT 4.400 370.920 395.600 370.960 ;
        RECT 3.990 369.560 395.600 370.920 ;
        RECT 3.990 368.240 396.000 369.560 ;
        RECT 4.400 366.880 396.000 368.240 ;
        RECT 4.400 366.840 395.600 366.880 ;
        RECT 3.990 365.480 395.600 366.840 ;
        RECT 3.990 364.160 396.000 365.480 ;
        RECT 4.400 362.800 396.000 364.160 ;
        RECT 4.400 362.760 395.600 362.800 ;
        RECT 3.990 361.400 395.600 362.760 ;
        RECT 3.990 360.080 396.000 361.400 ;
        RECT 4.400 358.720 396.000 360.080 ;
        RECT 4.400 358.680 395.600 358.720 ;
        RECT 3.990 357.320 395.600 358.680 ;
        RECT 3.990 356.000 396.000 357.320 ;
        RECT 4.400 354.640 396.000 356.000 ;
        RECT 4.400 354.600 395.600 354.640 ;
        RECT 3.990 353.240 395.600 354.600 ;
        RECT 3.990 351.920 396.000 353.240 ;
        RECT 4.400 350.560 396.000 351.920 ;
        RECT 4.400 350.520 395.600 350.560 ;
        RECT 3.990 349.160 395.600 350.520 ;
        RECT 3.990 347.840 396.000 349.160 ;
        RECT 4.400 346.480 396.000 347.840 ;
        RECT 4.400 346.440 395.600 346.480 ;
        RECT 3.990 345.080 395.600 346.440 ;
        RECT 3.990 343.760 396.000 345.080 ;
        RECT 4.400 342.400 396.000 343.760 ;
        RECT 4.400 342.360 395.600 342.400 ;
        RECT 3.990 341.000 395.600 342.360 ;
        RECT 3.990 339.680 396.000 341.000 ;
        RECT 4.400 338.320 396.000 339.680 ;
        RECT 4.400 338.280 395.600 338.320 ;
        RECT 3.990 336.920 395.600 338.280 ;
        RECT 3.990 335.600 396.000 336.920 ;
        RECT 4.400 334.240 396.000 335.600 ;
        RECT 4.400 334.200 395.600 334.240 ;
        RECT 3.990 332.840 395.600 334.200 ;
        RECT 3.990 331.520 396.000 332.840 ;
        RECT 4.400 330.160 396.000 331.520 ;
        RECT 4.400 330.120 395.600 330.160 ;
        RECT 3.990 328.760 395.600 330.120 ;
        RECT 3.990 327.440 396.000 328.760 ;
        RECT 4.400 326.080 396.000 327.440 ;
        RECT 4.400 326.040 395.600 326.080 ;
        RECT 3.990 324.680 395.600 326.040 ;
        RECT 3.990 323.360 396.000 324.680 ;
        RECT 4.400 322.000 396.000 323.360 ;
        RECT 4.400 321.960 395.600 322.000 ;
        RECT 3.990 320.600 395.600 321.960 ;
        RECT 3.990 319.280 396.000 320.600 ;
        RECT 4.400 317.920 396.000 319.280 ;
        RECT 4.400 317.880 395.600 317.920 ;
        RECT 3.990 316.520 395.600 317.880 ;
        RECT 3.990 315.200 396.000 316.520 ;
        RECT 4.400 313.840 396.000 315.200 ;
        RECT 4.400 313.800 395.600 313.840 ;
        RECT 3.990 312.440 395.600 313.800 ;
        RECT 3.990 311.120 396.000 312.440 ;
        RECT 4.400 309.760 396.000 311.120 ;
        RECT 4.400 309.720 395.600 309.760 ;
        RECT 3.990 308.360 395.600 309.720 ;
        RECT 3.990 307.040 396.000 308.360 ;
        RECT 4.400 305.680 396.000 307.040 ;
        RECT 4.400 305.640 395.600 305.680 ;
        RECT 3.990 304.280 395.600 305.640 ;
        RECT 3.990 302.960 396.000 304.280 ;
        RECT 4.400 301.600 396.000 302.960 ;
        RECT 4.400 301.560 395.600 301.600 ;
        RECT 3.990 300.200 395.600 301.560 ;
        RECT 3.990 298.880 396.000 300.200 ;
        RECT 4.400 297.520 396.000 298.880 ;
        RECT 4.400 297.480 395.600 297.520 ;
        RECT 3.990 296.120 395.600 297.480 ;
        RECT 3.990 294.800 396.000 296.120 ;
        RECT 4.400 293.440 396.000 294.800 ;
        RECT 4.400 293.400 395.600 293.440 ;
        RECT 3.990 292.040 395.600 293.400 ;
        RECT 3.990 290.720 396.000 292.040 ;
        RECT 4.400 289.360 396.000 290.720 ;
        RECT 4.400 289.320 395.600 289.360 ;
        RECT 3.990 287.960 395.600 289.320 ;
        RECT 3.990 286.640 396.000 287.960 ;
        RECT 4.400 285.280 396.000 286.640 ;
        RECT 4.400 285.240 395.600 285.280 ;
        RECT 3.990 283.880 395.600 285.240 ;
        RECT 3.990 282.560 396.000 283.880 ;
        RECT 4.400 281.200 396.000 282.560 ;
        RECT 4.400 281.160 395.600 281.200 ;
        RECT 3.990 279.800 395.600 281.160 ;
        RECT 3.990 278.480 396.000 279.800 ;
        RECT 4.400 277.120 396.000 278.480 ;
        RECT 4.400 277.080 395.600 277.120 ;
        RECT 3.990 275.720 395.600 277.080 ;
        RECT 3.990 274.400 396.000 275.720 ;
        RECT 4.400 273.040 396.000 274.400 ;
        RECT 4.400 273.000 395.600 273.040 ;
        RECT 3.990 271.640 395.600 273.000 ;
        RECT 3.990 270.320 396.000 271.640 ;
        RECT 4.400 268.960 396.000 270.320 ;
        RECT 4.400 268.920 395.600 268.960 ;
        RECT 3.990 267.560 395.600 268.920 ;
        RECT 3.990 266.240 396.000 267.560 ;
        RECT 4.400 264.880 396.000 266.240 ;
        RECT 4.400 264.840 395.600 264.880 ;
        RECT 3.990 263.480 395.600 264.840 ;
        RECT 3.990 262.160 396.000 263.480 ;
        RECT 4.400 260.800 396.000 262.160 ;
        RECT 4.400 260.760 395.600 260.800 ;
        RECT 3.990 259.400 395.600 260.760 ;
        RECT 3.990 258.080 396.000 259.400 ;
        RECT 4.400 256.720 396.000 258.080 ;
        RECT 4.400 256.680 395.600 256.720 ;
        RECT 3.990 255.320 395.600 256.680 ;
        RECT 3.990 254.000 396.000 255.320 ;
        RECT 4.400 252.640 396.000 254.000 ;
        RECT 4.400 252.600 395.600 252.640 ;
        RECT 3.990 251.240 395.600 252.600 ;
        RECT 3.990 249.920 396.000 251.240 ;
        RECT 4.400 248.560 396.000 249.920 ;
        RECT 4.400 248.520 395.600 248.560 ;
        RECT 3.990 247.160 395.600 248.520 ;
        RECT 3.990 245.840 396.000 247.160 ;
        RECT 4.400 244.480 396.000 245.840 ;
        RECT 4.400 244.440 395.600 244.480 ;
        RECT 3.990 243.080 395.600 244.440 ;
        RECT 3.990 241.760 396.000 243.080 ;
        RECT 4.400 240.400 396.000 241.760 ;
        RECT 4.400 240.360 395.600 240.400 ;
        RECT 3.990 239.000 395.600 240.360 ;
        RECT 3.990 237.680 396.000 239.000 ;
        RECT 4.400 236.320 396.000 237.680 ;
        RECT 4.400 236.280 395.600 236.320 ;
        RECT 3.990 234.920 395.600 236.280 ;
        RECT 3.990 233.600 396.000 234.920 ;
        RECT 4.400 232.240 396.000 233.600 ;
        RECT 4.400 232.200 395.600 232.240 ;
        RECT 3.990 230.840 395.600 232.200 ;
        RECT 3.990 229.520 396.000 230.840 ;
        RECT 4.400 228.160 396.000 229.520 ;
        RECT 4.400 228.120 395.600 228.160 ;
        RECT 3.990 226.760 395.600 228.120 ;
        RECT 3.990 225.440 396.000 226.760 ;
        RECT 4.400 224.080 396.000 225.440 ;
        RECT 4.400 224.040 395.600 224.080 ;
        RECT 3.990 222.680 395.600 224.040 ;
        RECT 3.990 221.360 396.000 222.680 ;
        RECT 4.400 220.000 396.000 221.360 ;
        RECT 4.400 219.960 395.600 220.000 ;
        RECT 3.990 218.600 395.600 219.960 ;
        RECT 3.990 217.280 396.000 218.600 ;
        RECT 4.400 215.920 396.000 217.280 ;
        RECT 4.400 215.880 395.600 215.920 ;
        RECT 3.990 214.520 395.600 215.880 ;
        RECT 3.990 213.200 396.000 214.520 ;
        RECT 4.400 211.840 396.000 213.200 ;
        RECT 4.400 211.800 395.600 211.840 ;
        RECT 3.990 210.440 395.600 211.800 ;
        RECT 3.990 209.120 396.000 210.440 ;
        RECT 4.400 207.760 396.000 209.120 ;
        RECT 4.400 207.720 395.600 207.760 ;
        RECT 3.990 206.360 395.600 207.720 ;
        RECT 3.990 205.040 396.000 206.360 ;
        RECT 4.400 203.680 396.000 205.040 ;
        RECT 4.400 203.640 395.600 203.680 ;
        RECT 3.990 202.280 395.600 203.640 ;
        RECT 3.990 200.960 396.000 202.280 ;
        RECT 4.400 199.600 396.000 200.960 ;
        RECT 4.400 199.560 395.600 199.600 ;
        RECT 3.990 198.200 395.600 199.560 ;
        RECT 3.990 196.880 396.000 198.200 ;
        RECT 4.400 195.520 396.000 196.880 ;
        RECT 4.400 195.480 395.600 195.520 ;
        RECT 3.990 194.120 395.600 195.480 ;
        RECT 3.990 192.800 396.000 194.120 ;
        RECT 4.400 191.440 396.000 192.800 ;
        RECT 4.400 191.400 395.600 191.440 ;
        RECT 3.990 190.040 395.600 191.400 ;
        RECT 3.990 188.720 396.000 190.040 ;
        RECT 4.400 187.360 396.000 188.720 ;
        RECT 4.400 187.320 395.600 187.360 ;
        RECT 3.990 185.960 395.600 187.320 ;
        RECT 3.990 184.640 396.000 185.960 ;
        RECT 4.400 183.280 396.000 184.640 ;
        RECT 4.400 183.240 395.600 183.280 ;
        RECT 3.990 181.880 395.600 183.240 ;
        RECT 3.990 180.560 396.000 181.880 ;
        RECT 4.400 179.200 396.000 180.560 ;
        RECT 4.400 179.160 395.600 179.200 ;
        RECT 3.990 177.800 395.600 179.160 ;
        RECT 3.990 176.480 396.000 177.800 ;
        RECT 4.400 175.120 396.000 176.480 ;
        RECT 4.400 175.080 395.600 175.120 ;
        RECT 3.990 173.720 395.600 175.080 ;
        RECT 3.990 172.400 396.000 173.720 ;
        RECT 4.400 171.040 396.000 172.400 ;
        RECT 4.400 171.000 395.600 171.040 ;
        RECT 3.990 169.640 395.600 171.000 ;
        RECT 3.990 168.320 396.000 169.640 ;
        RECT 4.400 166.960 396.000 168.320 ;
        RECT 4.400 166.920 395.600 166.960 ;
        RECT 3.990 165.560 395.600 166.920 ;
        RECT 3.990 164.240 396.000 165.560 ;
        RECT 4.400 162.880 396.000 164.240 ;
        RECT 4.400 162.840 395.600 162.880 ;
        RECT 3.990 161.480 395.600 162.840 ;
        RECT 3.990 160.160 396.000 161.480 ;
        RECT 4.400 158.800 396.000 160.160 ;
        RECT 4.400 158.760 395.600 158.800 ;
        RECT 3.990 157.400 395.600 158.760 ;
        RECT 3.990 156.080 396.000 157.400 ;
        RECT 4.400 154.720 396.000 156.080 ;
        RECT 4.400 154.680 395.600 154.720 ;
        RECT 3.990 153.320 395.600 154.680 ;
        RECT 3.990 152.000 396.000 153.320 ;
        RECT 4.400 150.640 396.000 152.000 ;
        RECT 4.400 150.600 395.600 150.640 ;
        RECT 3.990 149.240 395.600 150.600 ;
        RECT 3.990 147.920 396.000 149.240 ;
        RECT 4.400 146.560 396.000 147.920 ;
        RECT 4.400 146.520 395.600 146.560 ;
        RECT 3.990 145.160 395.600 146.520 ;
        RECT 3.990 143.840 396.000 145.160 ;
        RECT 4.400 142.480 396.000 143.840 ;
        RECT 4.400 142.440 395.600 142.480 ;
        RECT 3.990 141.080 395.600 142.440 ;
        RECT 3.990 139.760 396.000 141.080 ;
        RECT 4.400 138.400 396.000 139.760 ;
        RECT 4.400 138.360 395.600 138.400 ;
        RECT 3.990 137.000 395.600 138.360 ;
        RECT 3.990 135.680 396.000 137.000 ;
        RECT 4.400 134.320 396.000 135.680 ;
        RECT 4.400 134.280 395.600 134.320 ;
        RECT 3.990 132.920 395.600 134.280 ;
        RECT 3.990 131.600 396.000 132.920 ;
        RECT 4.400 130.240 396.000 131.600 ;
        RECT 4.400 130.200 395.600 130.240 ;
        RECT 3.990 128.840 395.600 130.200 ;
        RECT 3.990 127.520 396.000 128.840 ;
        RECT 4.400 126.160 396.000 127.520 ;
        RECT 4.400 126.120 395.600 126.160 ;
        RECT 3.990 124.760 395.600 126.120 ;
        RECT 3.990 123.440 396.000 124.760 ;
        RECT 4.400 122.080 396.000 123.440 ;
        RECT 4.400 122.040 395.600 122.080 ;
        RECT 3.990 120.680 395.600 122.040 ;
        RECT 3.990 119.360 396.000 120.680 ;
        RECT 4.400 118.000 396.000 119.360 ;
        RECT 4.400 117.960 395.600 118.000 ;
        RECT 3.990 116.600 395.600 117.960 ;
        RECT 3.990 115.280 396.000 116.600 ;
        RECT 4.400 113.920 396.000 115.280 ;
        RECT 4.400 113.880 395.600 113.920 ;
        RECT 3.990 112.520 395.600 113.880 ;
        RECT 3.990 111.200 396.000 112.520 ;
        RECT 4.400 109.840 396.000 111.200 ;
        RECT 4.400 109.800 395.600 109.840 ;
        RECT 3.990 108.440 395.600 109.800 ;
        RECT 3.990 107.120 396.000 108.440 ;
        RECT 4.400 105.760 396.000 107.120 ;
        RECT 4.400 105.720 395.600 105.760 ;
        RECT 3.990 104.360 395.600 105.720 ;
        RECT 3.990 103.040 396.000 104.360 ;
        RECT 4.400 101.680 396.000 103.040 ;
        RECT 4.400 101.640 395.600 101.680 ;
        RECT 3.990 100.280 395.600 101.640 ;
        RECT 3.990 98.960 396.000 100.280 ;
        RECT 4.400 97.600 396.000 98.960 ;
        RECT 4.400 97.560 395.600 97.600 ;
        RECT 3.990 96.200 395.600 97.560 ;
        RECT 3.990 94.880 396.000 96.200 ;
        RECT 4.400 93.520 396.000 94.880 ;
        RECT 4.400 93.480 395.600 93.520 ;
        RECT 3.990 92.120 395.600 93.480 ;
        RECT 3.990 90.800 396.000 92.120 ;
        RECT 4.400 89.440 396.000 90.800 ;
        RECT 4.400 89.400 395.600 89.440 ;
        RECT 3.990 88.040 395.600 89.400 ;
        RECT 3.990 86.720 396.000 88.040 ;
        RECT 4.400 85.360 396.000 86.720 ;
        RECT 4.400 85.320 395.600 85.360 ;
        RECT 3.990 83.960 395.600 85.320 ;
        RECT 3.990 82.640 396.000 83.960 ;
        RECT 4.400 81.280 396.000 82.640 ;
        RECT 4.400 81.240 395.600 81.280 ;
        RECT 3.990 79.880 395.600 81.240 ;
        RECT 3.990 78.560 396.000 79.880 ;
        RECT 4.400 77.200 396.000 78.560 ;
        RECT 4.400 77.160 395.600 77.200 ;
        RECT 3.990 75.800 395.600 77.160 ;
        RECT 3.990 74.480 396.000 75.800 ;
        RECT 4.400 73.120 396.000 74.480 ;
        RECT 4.400 73.080 395.600 73.120 ;
        RECT 3.990 71.720 395.600 73.080 ;
        RECT 3.990 70.400 396.000 71.720 ;
        RECT 4.400 69.040 396.000 70.400 ;
        RECT 4.400 69.000 395.600 69.040 ;
        RECT 3.990 67.640 395.600 69.000 ;
        RECT 3.990 66.320 396.000 67.640 ;
        RECT 4.400 64.960 396.000 66.320 ;
        RECT 4.400 64.920 395.600 64.960 ;
        RECT 3.990 63.560 395.600 64.920 ;
        RECT 3.990 62.240 396.000 63.560 ;
        RECT 4.400 60.880 396.000 62.240 ;
        RECT 4.400 60.840 395.600 60.880 ;
        RECT 3.990 59.480 395.600 60.840 ;
        RECT 3.990 58.160 396.000 59.480 ;
        RECT 4.400 56.800 396.000 58.160 ;
        RECT 4.400 56.760 395.600 56.800 ;
        RECT 3.990 55.400 395.600 56.760 ;
        RECT 3.990 54.080 396.000 55.400 ;
        RECT 4.400 52.720 396.000 54.080 ;
        RECT 4.400 52.680 395.600 52.720 ;
        RECT 3.990 51.320 395.600 52.680 ;
        RECT 3.990 50.000 396.000 51.320 ;
        RECT 4.400 48.640 396.000 50.000 ;
        RECT 4.400 48.600 395.600 48.640 ;
        RECT 3.990 47.240 395.600 48.600 ;
        RECT 3.990 45.920 396.000 47.240 ;
        RECT 4.400 44.560 396.000 45.920 ;
        RECT 4.400 44.520 395.600 44.560 ;
        RECT 3.990 43.160 395.600 44.520 ;
        RECT 3.990 41.840 396.000 43.160 ;
        RECT 4.400 40.480 396.000 41.840 ;
        RECT 4.400 40.440 395.600 40.480 ;
        RECT 3.990 39.080 395.600 40.440 ;
        RECT 3.990 37.760 396.000 39.080 ;
        RECT 4.400 36.400 396.000 37.760 ;
        RECT 4.400 36.360 395.600 36.400 ;
        RECT 3.990 35.000 395.600 36.360 ;
        RECT 3.990 33.680 396.000 35.000 ;
        RECT 4.400 32.320 396.000 33.680 ;
        RECT 4.400 32.280 395.600 32.320 ;
        RECT 3.990 30.920 395.600 32.280 ;
        RECT 3.990 29.600 396.000 30.920 ;
        RECT 4.400 28.200 396.000 29.600 ;
        RECT 3.990 25.520 396.000 28.200 ;
        RECT 4.400 24.120 396.000 25.520 ;
        RECT 3.990 10.715 396.000 24.120 ;
      LAYER met4 ;
        RECT 5.815 26.015 20.640 401.025 ;
        RECT 23.040 26.015 97.440 401.025 ;
        RECT 99.840 26.015 174.240 401.025 ;
        RECT 176.640 26.015 251.040 401.025 ;
        RECT 253.440 26.015 327.840 401.025 ;
        RECT 330.240 26.015 383.345 401.025 ;
  END
END multiplexer
END LIBRARY

