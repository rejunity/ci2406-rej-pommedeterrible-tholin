* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_mask[0]
+ dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0] dest_val[10]
+ dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16] dest_val[17]
+ dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22] dest_val[23]
+ dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29] dest_val[2]
+ dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6] dest_val[7]
+ dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11] instruction[12]
+ instruction[13] instruction[14] instruction[15] instruction[16] instruction[17]
+ instruction[18] instruction[19] instruction[1] instruction[20] instruction[21] instruction[22]
+ instruction[23] instruction[24] instruction[25] instruction[26] instruction[27]
+ instruction[28] instruction[29] instruction[2] instruction[30] instruction[31] instruction[32]
+ instruction[33] instruction[34] instruction[35] instruction[36] instruction[37]
+ instruction[38] instruction[39] instruction[3] instruction[40] instruction[41] instruction[4]
+ instruction[5] instruction[6] instruction[7] instruction[8] instruction[9] is_load
+ is_store loadstore_address[0] loadstore_address[10] loadstore_address[11] loadstore_address[12]
+ loadstore_address[13] loadstore_address[14] loadstore_address[15] loadstore_address[16]
+ loadstore_address[17] loadstore_address[18] loadstore_address[19] loadstore_address[1]
+ loadstore_address[20] loadstore_address[21] loadstore_address[22] loadstore_address[23]
+ loadstore_address[24] loadstore_address[25] loadstore_address[26] loadstore_address[27]
+ loadstore_address[28] loadstore_address[29] loadstore_address[2] loadstore_address[30]
+ loadstore_address[31] loadstore_address[3] loadstore_address[4] loadstore_address[5]
+ loadstore_address[6] loadstore_address[7] loadstore_address[8] loadstore_address[9]
+ loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3] loadstore_dest[4]
+ loadstore_size[0] loadstore_size[1] new_PC[0] new_PC[10] new_PC[11] new_PC[12] new_PC[13]
+ new_PC[14] new_PC[15] new_PC[16] new_PC[17] new_PC[18] new_PC[19] new_PC[1] new_PC[20]
+ new_PC[21] new_PC[22] new_PC[23] new_PC[24] new_PC[25] new_PC[26] new_PC[27] new_PC[2]
+ new_PC[3] new_PC[4] new_PC[5] new_PC[6] new_PC[7] new_PC[8] new_PC[9] pred_idx[0]
+ pred_idx[1] pred_idx[2] pred_val reg1_idx[0] reg1_idx[1] reg1_idx[2] reg1_idx[3]
+ reg1_idx[4] reg1_val[0] reg1_val[10] reg1_val[11] reg1_val[12] reg1_val[13] reg1_val[14]
+ reg1_val[15] reg1_val[16] reg1_val[17] reg1_val[18] reg1_val[19] reg1_val[1] reg1_val[20]
+ reg1_val[21] reg1_val[22] reg1_val[23] reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27]
+ reg1_val[28] reg1_val[29] reg1_val[2] reg1_val[30] reg1_val[31] reg1_val[3] reg1_val[4]
+ reg1_val[5] reg1_val[6] reg1_val[7] reg1_val[8] reg1_val[9] reg2_idx[0] reg2_idx[1]
+ reg2_idx[2] reg2_idx[3] reg2_idx[4] reg2_val[0] reg2_val[10] reg2_val[11] reg2_val[12]
+ reg2_val[13] reg2_val[14] reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18] reg2_val[19]
+ reg2_val[1] reg2_val[20] reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24] reg2_val[25]
+ reg2_val[26] reg2_val[27] reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30] reg2_val[31]
+ reg2_val[3] reg2_val[4] reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8] reg2_val[9]
+ rst sign_extend take_branch vccd1 vssd1 wb_clk_i
X_06883_ instruction[27] _06887_/B vssd1 vssd1 vccd1 vccd1 _06883_/X sky130_fd_sc_hd__or2_1
X_09671_ _11153_/A _09667_/X _09668_/X _09670_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a22o_4
X_08622_ _08622_/A _08624_/A _08622_/C vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__or3_1
XANTENNA__09304__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09287__A1 _09617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _08553_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08843_/B sky130_fd_sc_hd__nor2_1
X_07504_ _07504_/A _07504_/B vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout162_A _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ _08801_/A _08484_/B vssd1 vssd1 vccd1 vccd1 _08490_/A sky130_fd_sc_hd__xnor2_1
X_07435_ _07541_/B _07541_/A vssd1 vssd1 vccd1 vccd1 _07435_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_92_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__B2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ _07366_/A _07366_/B vssd1 vssd1 vccd1 vccd1 _07368_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08444__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09105_ _10920_/A reg1_val[18] _09120_/S vssd1 vssd1 vccd1 vccd1 _09105_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07297_ reg1_val[13] _07091_/B _07091_/C _07087_/B _07128_/A vssd1 vssd1 vccd1 vccd1
+ _07298_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_5_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09036_ _09001_/A _09001_/B _08842_/A vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06899__A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07222__B1 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _10201_/S _09311_/X _09937_/Y vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07773__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09869_ _10156_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__xor2_1
X_12880_ _13071_/A hold192/X vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__and2_1
X_11900_ _11973_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11902_/C sky130_fd_sc_hd__and2_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11831_ _11871_/B _11869_/C vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__nand2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ _11834_/D _11761_/B _12113_/A vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _11691_/Y _11693_/B vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__and2b_1
X_10713_ _10203_/S _09793_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10713_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _10644_/A _10644_/B vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__nor2_1
X_10575_ _10461_/A _10458_/Y _10460_/B vssd1 vssd1 vccd1 vccd1 _10577_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07461__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _12299_/X _12300_/Y _12303_/X _12313_/X vssd1 vssd1 vccd1 vccd1 _12314_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10596__B1 _10595_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12245_ _12245_/A _12245_/B fanout4/A vssd1 vssd1 vccd1 vccd1 _12248_/C sky130_fd_sc_hd__or3_1
X_12176_ _12175_/A _12175_/B _12175_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12195_/A
+ sky130_fd_sc_hd__o211a_1
X_11127_ _06831_/A _11126_/X _09498_/A vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09505__A2 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10009_/A fanout4/X vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07152__B _07152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07220_ _10009_/A _12714_/A _12716_/A _09725_/B2 vssd1 vssd1 vccd1 vccd1 _07221_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _07149_/A _07149_/B _07152_/B vssd1 vssd1 vccd1 vccd1 _07156_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__B1 _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ _07082_/A _07082_/B vssd1 vssd1 vccd1 vccd1 _07339_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09992__A2 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11536__C1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 _08606_/A2 vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__buf_6
Xfanout127 _06960_/Y vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__buf_6
Xfanout138 _11072_/A vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__clkbuf_16
Xfanout105 _07916_/A vssd1 vssd1 vccd1 vccd1 _11656_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout149 _07111_/X vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__buf_8
X_07984_ _07984_/A _07984_/B _07984_/C vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06935_ _06963_/B _06936_/C _06936_/A vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__o21ai_4
X_09723_ _09724_/A _09724_/B vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__nand2_1
X_06866_ instruction[13] _06868_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
X_09654_ _06834_/B _09652_/X _09653_/Y vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08605_ _08605_/A _08605_/B vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08439__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06797_ _06796_/A _06796_/B _06837_/A vssd1 vssd1 vccd1 vccd1 _06798_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ _10490_/B2 _11564_/A fanout38/X fanout80/X vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11067__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _08563_/A _08563_/B _08532_/X vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11067__B2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ _08427_/B _08427_/C _08427_/D _08427_/A vssd1 vssd1 vccd1 vccd1 _08467_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__08483__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07418_ _09880_/B2 _11564_/A fanout38/X _10117_/A vssd1 vssd1 vccd1 vccd1 _07419_/B
+ sky130_fd_sc_hd__o22a_1
X_08398_ _08741_/A _08398_/B vssd1 vssd1 vccd1 vccd1 _08401_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07438_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08174__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__C1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _11799_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__xnor2_1
X_09019_ _09019_/A _09019_/B vssd1 vssd1 vccd1 vccd1 _10187_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07994__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__B2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ _10165_/A _10164_/B _10164_/A vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ _12030_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__xor2_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10750__B1 _07277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ _11184_/B _12962_/B2 hold89/X vssd1 vssd1 vccd1 vccd1 _13207_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07253__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__B2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__A1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ hold205/X _13070_/B2 _13070_/A2 hold171/X vssd1 vssd1 vccd1 vccd1 hold206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12794_ _12971_/B _12972_/A _12787_/X vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__a21o_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11814_ _11895_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11816_/B sky130_fd_sc_hd__or2_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09671__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07682__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06522__C_N _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11676_ _11677_/A _11677_/B _11677_/C vssd1 vssd1 vccd1 vccd1 _11757_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08084__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ _10793_/B _10558_/B vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_12_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _12269_/B _12227_/Y _12271_/S vssd1 vssd1 vccd1 vccd1 _12228_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07428__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _10663_/B _10489_/B vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _12159_/A vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__inv_2
XANTENNA__10741__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ reg2_val[6] _06748_/B vssd1 vssd1 vccd1 vccd1 _06720_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06651_ reg1_val[17] _06978_/A vssd1 vssd1 vccd1 vccd1 _06653_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06582_ reg2_val[29] _06700_/B _06657_/B1 _06581_/X vssd1 vssd1 vccd1 vccd1 _06801_/B
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__11049__B2 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11049__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__B1 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ _09370_/A _09370_/B _09370_/C vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08321_ _08244_/A _08244_/C _08244_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08996_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _07203_/A _07203_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08217__A2 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout125_A _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _08189_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__B1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ _07132_/A _07132_/B _07132_/C _07132_/D vssd1 vssd1 vccd1 vccd1 _11727_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09965__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07065_ _07065_/A _07065_/B _07065_/C _07065_/D vssd1 vssd1 vccd1 vccd1 _07068_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09178__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07967_ _07967_/A _07967_/B vssd1 vssd1 vccd1 vccd1 _07976_/B sky130_fd_sc_hd__xor2_1
X_06918_ reg1_val[10] reg1_val[11] _06993_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _06919_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__11288__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _10607_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__xnor2_2
X_07898_ _07898_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _07899_/B sky130_fd_sc_hd__and2_1
XANTENNA__09350__B1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ instruction[1] _06850_/B instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06887_/B sky130_fd_sc_hd__and4b_4
X_09637_ _09629_/X _09636_/X _10809_/A vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12237__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09568_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07801__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout38_A _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ _08519_/A _08519_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__nor2_1
X_11530_ _11620_/B _11619_/B hold168/A vssd1 vssd1 vccd1 vccd1 _11530_/Y sky130_fd_sc_hd__a21oi_1
X_09499_ _13160_/Q hold189/A _12190_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout4_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08208__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ _11579_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11462_/C sky130_fd_sc_hd__or2_1
X_13200_ _13222_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07416__B1 _07304_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11392_ _11393_/A _11393_/B vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10015__A2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09728__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ fanout78/X _12095_/A fanout60/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10413_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12960__A1 _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _13253_/CLK _13131_/D vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
X_10343_ hold200/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ _13062_/A hold264/X vssd1 vssd1 vccd1 vccd1 _13243_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _10272_/Y _10274_/B vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__and2b_1
X_12013_ _12080_/A _12010_/X _12011_/X _12012_/Y vssd1 vssd1 vccd1 vccd1 dest_val[25]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09341__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ hold119/X _12662_/A _13112_/B _13199_/Q _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold120/A sky130_fd_sc_hd__o221a_1
XFILLER_0_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ _13071_/A hold223/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__and2_1
XANTENNA__12228__B1 _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ hold68/X hold285/X vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__and2b_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12329__A _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08447__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _07133_/Y _11385_/B _11727_/X _11796_/A vssd1 vssd1 vccd1 vccd1 _11730_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11660_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07158__A _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10962__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ _08870_/A _08870_/B vssd1 vssd1 vccd1 vccd1 _08870_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08907__B1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _07821_/A _07821_/B vssd1 vssd1 vccd1 vccd1 _07823_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06933__A2 _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__B _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _07811_/B _07752_/B _07750_/X vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__or3b_1
X_06703_ reg1_val[9] _07289_/A vssd1 vssd1 vccd1 vccd1 _06777_/A sky130_fd_sc_hd__nand2_1
X_07683_ _08916_/A _07683_/B vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__xnor2_1
X_06634_ reg1_val[19] _06980_/A vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _09422_/A fanout4/X vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09312__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _11636_/S _09351_/X _09352_/Y _09350_/X vssd1 vssd1 vccd1 vccd1 dest_val[1]
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06565_ reg1_val[25] _07059_/A vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08304_ _08304_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08438__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _08982_/A _09461_/A _08980_/Y vssd1 vssd1 vccd1 vccd1 _09285_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_90_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08235_ _11068_/A _08309_/A _08233_/X vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ _08166_/A _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__and2_1
XANTENNA__12942__A1 _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ _07284_/B _07118_/C reg1_val[23] vssd1 vssd1 vccd1 vccd1 _07149_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08097_ _08242_/A _08096_/Y _08092_/Y vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08071__B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _07065_/A _07065_/B _06578_/B _07058_/B1 vssd1 vssd1 vccd1 vccd1 _07048_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12702__A _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _09001_/A _09001_/B _09037_/A _08555_/Y vssd1 vssd1 vccd1 vccd1 _09000_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08126__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ _10961_/A _10961_/B vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07234__C _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ hold66/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ _12656_/A _07176_/C _12640_/B vssd1 vssd1 vccd1 vccd1 _12632_/B sky130_fd_sc_hd__a21bo_2
X_10892_ _10892_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10894_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ _12562_/A _12562_/B _12562_/C vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ _12493_/A _12493_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11513_ _12110_/A _11603_/C vssd1 vssd1 vccd1 vccd1 _11514_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11444_ hold287/A _11623_/B _11532_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11197__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ fanout17/X _11564_/A fanout38/X fanout9/A vssd1 vssd1 vccd1 vccd1 _11376_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08062__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ hold164/X _12663_/B _12657_/Y _12664_/A vssd1 vssd1 vccd1 vccd1 _13114_/X
+ sky130_fd_sc_hd__a22o_1
X_10326_ _10449_/A _09021_/A _09021_/B _12179_/A vssd1 vssd1 vccd1 vccd1 _10327_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13045_/A _13045_/B vssd1 vssd1 vccd1 vccd1 _13045_/Y sky130_fd_sc_hd__xnor2_1
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__xor2_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07168__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10188_ _10449_/A _10187_/C _10187_/B vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07441__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ _13095_/A _12828_/B _12828_/A vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07628__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _08167_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12924__A1 _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__B _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout7 fanout8/X vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _11796_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__xnor2_2
X_08922_ _11184_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08924_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07159__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _07689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _08853_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07828_/B sky130_fd_sc_hd__xnor2_2
X_08784_ _08784_/A _08784_/B _08784_/C vssd1 vssd1 vccd1 vccd1 _08792_/A sky130_fd_sc_hd__and3_1
X_07735_ _07735_/A _07735_/B _07735_/C vssd1 vssd1 vccd1 vccd1 _07736_/B sky130_fd_sc_hd__nand3_1
X_07666_ _07666_/A _07759_/A vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07351__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _09405_/A _09405_/B vssd1 vssd1 vccd1 vccd1 _09406_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06617_ reg1_val[21] _06987_/A vssd1 vssd1 vccd1 vccd1 _11704_/S sky130_fd_sc_hd__and2_1
X_07597_ _09422_/A _07070_/Y _12201_/A _09222_/B2 vssd1 vssd1 vccd1 vccd1 _07598_/B
+ sky130_fd_sc_hd__o22a_2
X_06548_ _06613_/A _12553_/B vssd1 vssd1 vccd1 vccd1 _06548_/X sky130_fd_sc_hd__or2_1
X_09336_ _12499_/A _09336_/B _12668_/A vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__or3_1
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07070__B _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _09267_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _09268_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_90_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ _08276_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08223_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _09198_/A _09198_/B vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ _08149_/A _08149_/B _08149_/C vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__and3_1
XFILLER_0_15_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _11160_/A _11160_/B _11160_/C vssd1 vssd1 vccd1 vccd1 _11160_/X sky130_fd_sc_hd__and3_1
X_10111_ _10111_/A _10111_/B vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__xnor2_4
X_11091_ _11091_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12143__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _10043_/B _10043_/A vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09544__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _11991_/Y _11993_/B vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_98_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _11636_/S _10941_/X _10943_/Y vssd1 vssd1 vccd1 vccd1 dest_val[13] sky130_fd_sc_hd__o21ai_4
XFILLER_0_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10875_ _10876_/A1 _12029_/B _10875_/C vssd1 vssd1 vccd1 vccd1 _10997_/B sky130_fd_sc_hd__and3b_1
X_12614_ _12611_/A _12613_/B _12611_/B vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ reg1_val[10] _12546_/B vssd1 vssd1 vccd1 vccd1 _12547_/A sky130_fd_sc_hd__or2_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12906__A1 _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ reg1_val[24] curr_PC[24] _12495_/S vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 curr_PC[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _11838_/A _11426_/C _11426_/B vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _09293_/A _11035_/Y _11353_/X _11357_/X vssd1 vssd1 vccd1 vccd1 _11358_/X
+ sky130_fd_sc_hd__o211a_1
X_10309_ _10309_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__nand2_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11289_ _11799_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11291_/B sky130_fd_sc_hd__xnor2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _13103_/A _13028_/B vssd1 vssd1 vccd1 vccd1 _13236_/D sky130_fd_sc_hd__and2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07561__A2 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _07670_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__or2_1
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ _09862_/B _07451_/B vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__xnor2_2
X_07382_ _06828_/A _12094_/A _08765_/A _12720_/A vssd1 vssd1 vccd1 vccd1 _07383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ reg1_val[5] reg1_val[26] _09124_/S vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08813__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09052_ _11838_/B _09052_/B _09052_/C _09052_/D vssd1 vssd1 vccd1 vccd1 _09056_/C
+ sky130_fd_sc_hd__or4_2
X_08003_ _08607_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08010_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap230 _07186_/A vssd1 vssd1 vccd1 vccd1 _09630_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09826__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09954_ _09498_/A _09926_/Y _09942_/X _09953_/X vssd1 vssd1 vccd1 vccd1 _09954_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08329__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ _06977_/A fanout65/X fanout58/X _06985_/A vssd1 vssd1 vccd1 vccd1 _08906_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11333__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10136__B2 _11091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A1 _08384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _09885_/A _11885_/A _09886_/A vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__or3_1
XANTENNA__07001__A1 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _09004_/A _09004_/B _09025_/A _08834_/Y vssd1 vssd1 vccd1 vccd1 _09003_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11884__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08767_ _08768_/B _08768_/C _09420_/A vssd1 vssd1 vccd1 vccd1 _08771_/C sky130_fd_sc_hd__a21o_1
X_07718_ _07830_/A _07830_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07722_/A sky130_fd_sc_hd__nand3_1
X_08698_ _08698_/A _08698_/B vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__xnor2_2
X_09319_ _09121_/X _09123_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09319_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _07296_/A _12238_/C1 _10589_/Y _10590_/X vssd1 vssd1 vccd1 vccd1 _10591_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_105_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ _12507_/B _12330_/B vssd1 vssd1 vccd1 vccd1 _12331_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__and2_1
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08568__A1 _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _11212_/A _11212_/B _11212_/C vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__and3_1
X_12192_ _06591_/X _09147_/X _12191_/Y _06593_/B _12280_/A vssd1 vssd1 vccd1 vccd1
+ _12192_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_101_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11143_ _09147_/X _09141_/Y _11143_/S vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07240__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A1_N _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ _11075_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__or2_1
XANTENNA__11875__A1 _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _10159_/B _10025_/B vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__or2_1
XANTENNA__08740__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11976_ _11976_/A _11976_/B _11976_/C vssd1 vssd1 vccd1 vccd1 _11978_/A sky130_fd_sc_hd__nand3_1
X_10927_ hold207/A _10927_/B vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08815__A _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10858_ _11739_/A fanout50/X _07988_/B fanout64/X vssd1 vssd1 vccd1 vccd1 _10859_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12337__A _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ _10790_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10791_/A sky130_fd_sc_hd__nor2_1
X_12528_ _12526_/Y _12528_/B vssd1 vssd1 vccd1 vccd1 _12529_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12459_ reg1_val[21] curr_PC[21] _12495_/S vssd1 vssd1 vccd1 vccd1 _12460_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06951_ _10920_/A reg1_val[14] _07091_/B _07128_/A vssd1 vssd1 vccd1 vccd1 _06952_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ _11153_/A _09957_/C vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__nor2_1
X_06882_ instruction[19] _06850_/Y _06881_/X _06637_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09381__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _08622_/A _08624_/A _08622_/C vssd1 vssd1 vccd1 vccd1 _08621_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08552_ _08841_/B _08841_/C _08841_/A vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__a21oi_1
X_07503_ _07503_/A _07503_/B vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _08782_/A2 _08689_/B1 _09180_/B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08484_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11850__S _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _07434_/A _07434_/B vssd1 vssd1 vccd1 vccd1 _07541_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07365_ _07364_/B _07364_/C _07364_/A vssd1 vssd1 vccd1 vccd1 _07366_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ _07296_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _07296_/Y sky130_fd_sc_hd__xnor2_1
X_09104_ reg1_val[12] reg1_val[19] _09120_/S vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10054__B1 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__B1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _11236_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07222__B2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09320_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09937_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07773__A2 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12710__A _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ fanout78/X fanout68/X fanout65/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _09869_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09799_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__or2_1
X_08819_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__xnor2_1
X_11830_ _11830_/A vssd1 vssd1 vccd1 vccd1 _11869_/C sky130_fd_sc_hd__inv_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11761_ _11834_/D _11761_/B vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__nand2_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10704_/Y _10705_/X _10710_/X _10711_/Y vssd1 vssd1 vccd1 vccd1 _10712_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10644_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_118_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10574_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11061__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _12313_/A1 _12305_/Y _12308_/X _12312_/X vssd1 vssd1 vccd1 vccd1 _12313_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07461__A1 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__B1 _07112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07461__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ _12203_/A _12203_/B _12202_/B vssd1 vssd1 vccd1 vccd1 _12250_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11545__B1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ _11238_/A _11125_/X _11124_/X vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06972__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _11654_/A _11057_/B vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__xnor2_1
X_10008_ _10252_/A _10008_/B vssd1 vssd1 vccd1 vccd1 _10011_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12273__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _12085_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _07916_/A _07152_/B vssd1 vssd1 vccd1 vccd1 _07150_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10587__A1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07452__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07081_ _07081_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07082_/B sky130_fd_sc_hd__or2_1
XFILLER_0_54_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__B2 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout117 _06997_/X vssd1 vssd1 vccd1 vccd1 _08606_/A2 sky130_fd_sc_hd__buf_8
Xfanout128 _11169_/A vssd1 vssd1 vccd1 vccd1 _10099_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout106 _07916_/A vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__clkbuf_8
Xfanout139 _07232_/X vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__buf_8
X_07983_ _07913_/A _07913_/C _07913_/B vssd1 vssd1 vccd1 vccd1 _07984_/C sky130_fd_sc_hd__a21o_1
X_09722_ _09979_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09724_/B sky130_fd_sc_hd__xnor2_1
X_06934_ _12115_/A _07184_/B _06963_/A vssd1 vssd1 vccd1 vccd1 _06936_/C sky130_fd_sc_hd__and3_1
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout272_A _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06865_ instruction[12] _06868_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
X_09653_ _06834_/B _09652_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _09653_/Y sky130_fd_sc_hd__o21ai_1
X_08604_ _08616_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08617_/A sky130_fd_sc_hd__o21a_1
X_09584_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__xor2_1
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06796_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08535_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08563_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11067__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08466_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ _09979_/A _07417_/B vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__xnor2_1
X_08397_ _08740_/A2 _08689_/B1 _09180_/B2 _08755_/B vssd1 vssd1 vccd1 vccd1 _08398_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07348_ _07875_/A _07348_/B vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07279_ _12694_/A _08333_/B fanout92/X fanout42/X vssd1 vssd1 vccd1 vccd1 _07280_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10924__S _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07994__A2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__xnor2_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12931_ hold85/X _12665_/A _12955_/B1 hold83/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold89/A sky130_fd_sc_hd__o221a_1
XANTENNA__10502__A1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12862_ _13062_/A hold217/X vssd1 vssd1 vccd1 vccd1 _13172_/D sky130_fd_sc_hd__and2_1
XANTENNA__08171__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A3 _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ fanout65/X _11885_/A _11812_/C vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12793_ _12967_/A _12967_/B _12791_/A vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__a21o_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11744_ _11745_/B _11745_/A vssd1 vssd1 vccd1 vccd1 _11744_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12007__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__A1 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11677_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09671__A2 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ _11656_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__xor2_1
X_10557_ _10557_/A _10557_/B _10557_/C vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__nor3_1
XANTENNA__08631__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _10488_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__and2_1
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ reg1_val[28] _12226_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12227_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12191__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _12214_/A _12158_/B vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10741__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10741__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13251_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__12350__A _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12090_/A sky130_fd_sc_hd__xnor2_1
X_11109_ _11110_/A _11110_/B vssd1 vssd1 vccd1 vccd1 _11226_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06650_ reg1_val[17] _06978_/A vssd1 vssd1 vccd1 vccd1 _06653_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07370__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ _06646_/A _12571_/B vssd1 vssd1 vccd1 vccd1 _06581_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08251_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _07202_/A _07336_/A vssd1 vssd1 vccd1 vccd1 _07203_/B sky130_fd_sc_hd__or2_1
XFILLER_0_7_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08182_ _08193_/B _08182_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07425__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07425__B2 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07133_ _11796_/A _07138_/A vssd1 vssd1 vccd1 vccd1 _07133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07064_ _07064_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07065_/D sky130_fd_sc_hd__or2_1
XANTENNA_fanout118_A _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09178__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__A1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07966_ _07965_/B _07965_/C _07965_/A vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__a21bo_1
X_06917_ reg1_val[11] _06917_/B vssd1 vssd1 vccd1 vccd1 _06917_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__06951__A3 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08689__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _07000_/A fanout63/X fanout55/X _10481_/A vssd1 vssd1 vccd1 vccd1 _09706_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11288__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ _08986_/A vssd1 vssd1 vccd1 vccd1 _07897_/Y sky130_fd_sc_hd__inv_2
X_09636_ _09632_/X _09635_/Y _11134_/S vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__mux2_1
X_06848_ _06850_/B _06863_/A vssd1 vssd1 vccd1 vccd1 _06848_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_93_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06779_ _10689_/B _10689_/C _10692_/A vssd1 vssd1 vccd1 vccd1 _06779_/X sky130_fd_sc_hd__a21bo_1
X_09567_ _09567_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__xnor2_1
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07113__B1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ _08518_/A _08518_/B _08518_/C vssd1 vssd1 vccd1 vccd1 _08519_/B sky130_fd_sc_hd__and3_1
XANTENNA__11996__B1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06872__C1 _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11459_/B _11460_/B vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07416__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07416__B2 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ _11391_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11393_/B sky130_fd_sc_hd__and2_1
X_10411_ _11068_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ hold241/A _10465_/C _10208_/B vssd1 vssd1 vccd1 vccd1 _10343_/B sky130_fd_sc_hd__o21a_1
X_13130_ _13208_/CLK _13130_/D vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07529__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ hold263/X _13070_/A2 _13060_/X _13070_/B2 vssd1 vssd1 vccd1 vccd1 hold264/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__B2 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ curr_PC[25] _12079_/C _12080_/A vssd1 vssd1 vccd1 vccd1 _12012_/Y sky130_fd_sc_hd__a21oi_1
X_10273_ _10273_/A _10273_/B vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__nand2_1
X_12914_ _08698_/A _12692_/B hold145/X vssd1 vssd1 vccd1 vccd1 _13198_/D sky130_fd_sc_hd__a21boi_1
X_12845_ hold239/A _12885_/A2 _12885_/B1 hold222/X vssd1 vssd1 vccd1 vccd1 hold223/A
+ sky130_fd_sc_hd__a22o_1
X_12776_ hold289/X hold74/X vssd1 vssd1 vccd1 vccd1 _12994_/B sky130_fd_sc_hd__nand2b_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11727_ _11727_/A fanout3/X vssd1 vssd1 vccd1 vccd1 _11727_/X sky130_fd_sc_hd__or2_1
XANTENNA__08095__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11660_/A sky130_fd_sc_hd__or2_1
XFILLER_0_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11677_/A sky130_fd_sc_hd__and2_1
X_10609_ _10850_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10962__B2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10962__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ _13260_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12703__A2 _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__B2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _07824_/B _07824_/A vssd1 vssd1 vccd1 vccd1 _07823_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12080__A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ _07722_/A _07722_/B _07722_/C vssd1 vssd1 vccd1 vccd1 _07752_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06933__A3 _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__B1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _06763_/B _06646_/A _12546_/B _06700_/X vssd1 vssd1 vccd1 vccd1 _07289_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09332__A1 _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07682_ _06940_/A _12694_/A fanout92/X fanout82/X vssd1 vssd1 vccd1 vccd1 _07683_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06633_ reg1_val[19] _07002_/A vssd1 vssd1 vccd1 vccd1 _06790_/A sky130_fd_sc_hd__nand2_1
X_09421_ _09563_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__xnor2_2
X_06564_ _07059_/A reg1_val[25] vssd1 vssd1 vccd1 vccd1 _06566_/A sky130_fd_sc_hd__nand2b_1
X_09352_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _08299_/A _08299_/B _08355_/A vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout235_A _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09461_/B sky130_fd_sc_hd__xor2_4
X_08234_ _11068_/A _08309_/A _08233_/X vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10982__B fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07116_ reg1_val[22] _07128_/B _07128_/A vssd1 vssd1 vccd1 vccd1 _07118_/C sky130_fd_sc_hd__o21a_1
XANTENNA__08071__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ _08242_/B vssd1 vssd1 vccd1 vccd1 _08096_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08071__B2 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10953__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ _07065_/A _07065_/B _07058_/B1 vssd1 vssd1 vccd1 vccd1 _07047_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12702__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10503__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _11068_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07982_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08126__A2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08908__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10961_/A _10961_/B vssd1 vssd1 vccd1 vccd1 _11102_/B sky130_fd_sc_hd__nand2b_1
X_09619_ _11983_/A _09917_/B _10321_/A vssd1 vssd1 vccd1 vccd1 _09619_/Y sky130_fd_sc_hd__a21oi_1
X_10891_ _10890_/A _10890_/B _10892_/A vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__o21ai_1
X_12630_ _12630_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__or2_1
X_12561_ _12562_/A _12562_/B _12562_/C vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _12485_/B _12487_/B _12485_/A vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11509_/B _11422_/B _11233_/A _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1
+ _11603_/C sky130_fd_sc_hd__o2111a_1
X_11443_ _11623_/B _11532_/B hold287/A vssd1 vssd1 vccd1 vccd1 _11443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08062__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11197__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ hold100/X _12664_/A _13013_/A hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A
+ sky130_fd_sc_hd__o211a_1
X_11374_ _11799_/A _11374_/B vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08062__B2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ _10449_/A _09021_/B _09021_/A vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12697__A1 _08384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ _12755_/X _13044_/B vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__nand2b_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _10256_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06610__B _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _10449_/A _10187_/B _10187_/C vssd1 vssd1 vccd1 vccd1 _10187_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__10413__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__A2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _12828_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _13095_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ hold47/X hold273/A vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07628__B2 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06851__A2 _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07169__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10935__A1 _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout8 fanout8/A vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__buf_6
XANTENNA__09250__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07800__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09970_ fanout80/X fanout50/X fanout49/X _10099_/A1 vssd1 vssd1 vccd1 vccd1 _09971_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08921_ _10852_/B2 _11387_/A _10359_/B2 fanout79/X vssd1 vssd1 vccd1 vccd1 _08922_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__B _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _08996_/A _08995_/A _08849_/X _08851_/Y vssd1 vssd1 vccd1 vccd1 _09048_/C
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09553__A1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _07885_/A _07885_/B _07798_/A vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout185_A _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ _08801_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08784_/C sky130_fd_sc_hd__xor2_1
X_07734_ _07732_/A _07732_/B _07826_/A vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__xnor2_1
X_06616_ reg1_val[21] _07012_/A vssd1 vssd1 vccd1 vccd1 _06794_/A sky130_fd_sc_hd__nand2_1
X_09404_ _09405_/A _09405_/B vssd1 vssd1 vccd1 vccd1 _09404_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07596_ _07596_/A vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__inv_2
X_06547_ instruction[36] _06637_/B vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__and2_4
X_09335_ _13160_/Q hold189/A _12190_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _09335_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06827__C1 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _09266_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09267_/B sky130_fd_sc_hd__or2_1
XANTENNA__10623__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08217_ _11169_/A _08813_/A1 _12702_/A _06828_/A vssd1 vssd1 vccd1 vccd1 _08218_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09197_ _09198_/A _09198_/B vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__or2_2
XFILLER_0_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12679__A1 _07147_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10111_/B sky130_fd_sc_hd__xor2_4
X_11090_ _10971_/A _10971_/B _10968_/A vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__a21oi_1
X_10041_ _10041_/A _10041_/B vssd1 vssd1 vccd1 vccd1 _10043_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09544__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__nand2_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12300__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ curr_PC[13] _11051_/C _10942_/Y vssd1 vssd1 vccd1 vccd1 _10943_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10874_ _10997_/A _10874_/B vssd1 vssd1 vccd1 vccd1 _10875_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08807__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12613_ _12620_/C _12613_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ _12544_/A _12544_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
XFILLER_0_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10090__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12475_ _12478_/D _12475_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12906__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 curr_PC[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _11838_/A _11426_/B _11426_/C vssd1 vssd1 vccd1 vccd1 _11428_/A sky130_fd_sc_hd__and3_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ _12073_/B2 _11047_/Y _11355_/Y _11356_/X vssd1 vssd1 vccd1 vccd1 _11357_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12119__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10308_ _10308_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__xnor2_2
X_13027_ hold297/X _06858_/B _13026_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 _13028_/B
+ sky130_fd_sc_hd__a22o_1
X_11288_ _11876_/A fanout13/X fanout47/X _11950_/A vssd1 vssd1 vccd1 vccd1 _11289_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _12684_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07450_ _12710_/A _09727_/A _08798_/B _12712_/A vssd1 vssd1 vccd1 vccd1 _07451_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07381_ _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07393_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ reg1_val[4] reg1_val[27] _09120_/S vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12070__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12517__B _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ _08992_/A _08992_/B _11914_/C vssd1 vssd1 vccd1 vccd1 _09052_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08002_ _08606_/A2 _10506_/A _10647_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08003_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout100_A _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ _12073_/B2 _09940_/X _09952_/X _09293_/A _09950_/Y vssd1 vssd1 vccd1 vccd1
+ _09953_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08329__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10053__A _10321_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10136__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _09885_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11884__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08706_/X _08835_/B vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__and2b_1
X_08766_ _07147_/A _07147_/B _06828_/A vssd1 vssd1 vccd1 vccd1 _08768_/C sky130_fd_sc_hd__a21o_1
X_07717_ _07830_/A _07830_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__and3_1
XFILLER_0_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12294__C1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _08740_/A2 _08782_/B2 _08813_/B1 _08755_/B vssd1 vssd1 vccd1 vccd1 _08698_/B
+ sky130_fd_sc_hd__o22a_1
X_07648_ _07565_/B _07217_/B _07276_/B _07275_/B _07275_/A vssd1 vssd1 vccd1 vccd1
+ _07651_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07579_ _12095_/B _07579_/B vssd1 vssd1 vccd1 vccd1 _07585_/A sky130_fd_sc_hd__xnor2_2
X_09318_ _09117_/X _09120_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09318_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ hold277/A _09808_/B _10708_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _10590_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout13_A _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _08887_/Y _08890_/B _08895_/A vssd1 vssd1 vccd1 vccd1 _09264_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _12112_/A _12257_/Y _12258_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _12261_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09214__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ _06591_/X _09501_/B _09138_/X vssd1 vssd1 vccd1 vccd1 _12191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _11212_/A _11212_/B _11212_/C vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11021__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ hold218/A _11620_/B _11249_/B _11141_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1
+ _11142_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07240__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07528__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11073_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__xnor2_1
X_10024_ _10024_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__and2_1
XANTENNA__08740__A2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11627__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__C1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ _11976_/C vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10926_ _10923_/Y _10925_/X _11696_/A vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10835__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _10948_/B _10856_/C _10856_/A vssd1 vssd1 vccd1 vccd1 _10868_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08815__B _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10788_ _10674_/A _10674_/B _10672_/X vssd1 vssd1 vccd1 vccd1 _10790_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ reg1_val[6] _12527_/B vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ _12468_/A _12458_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XANTENNA__09205__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12389_ _12389_/A _12389_/B _12389_/C vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06950_ _10920_/A _07091_/B _07128_/A vssd1 vssd1 vccd1 vccd1 _06953_/B sky130_fd_sc_hd__o21a_1
X_06881_ instruction[26] _06887_/B vssd1 vssd1 vccd1 vccd1 _06881_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08622_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08278__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__B _10320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08841_/C sky130_fd_sc_hd__or2_1
X_07502_ _07675_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07508_/A sky130_fd_sc_hd__xnor2_1
X_08482_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08539_/A sky130_fd_sc_hd__nor2_1
X_07433_ _07429_/A _07429_/B _07522_/A vssd1 vssd1 vccd1 vccd1 _07541_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout148_A _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07364_ _07364_/A _07364_/B _07364_/C vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__and3_1
X_09103_ _09099_/X _09102_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09103_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07295_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/B sky130_fd_sc_hd__or2_1
XFILLER_0_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ _11122_/B _11122_/C vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__and2_1
XFILLER_0_103_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08741__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07222__A2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ _10924_/S _09934_/Y _09935_/Y _10809_/A vssd1 vssd1 vccd1 vccd1 _09936_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09867_ _10607_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__xnor2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09798_/Y sky130_fd_sc_hd__nor2_1
X_08818_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10511__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08749_ _08749_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08762_/A sky130_fd_sc_hd__xnor2_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _12110_/A _11834_/A _11834_/B _11834_/C _09621_/A vssd1 vssd1 vccd1 vccd1
+ _11761_/B sky130_fd_sc_hd__a41o_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _07304_/A _12238_/C1 _10707_/X vssd1 vssd1 vccd1 vccd1 _10711_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__08916__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10642_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10644_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10573_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10577_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07461__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ _09293_/A _09130_/Y _09330_/A _12302_/B _12311_/Y vssd1 vssd1 vccd1 vccd1
+ _12312_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11793__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__B2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ _06585_/B _06905_/Y _12242_/X _12080_/A vssd1 vssd1 vccd1 vccd1 dest_val[29]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12174_ _12115_/A _06803_/Y _06817_/X _12173_/X vssd1 vssd1 vccd1 vccd1 _12175_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07267__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _11026_/A _11024_/X _11043_/A vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__o21a_1
X_11056_ _12095_/A fanout41/X _08135_/B fanout60/X vssd1 vssd1 vccd1 vccd1 _11057_/B
+ sky130_fd_sc_hd__o22a_1
X_10007_ _06977_/A fanout17/X fanout9/X _06985_/A vssd1 vssd1 vccd1 vccd1 _10008_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11958_ fanout15/X fanout9/A fanout4/A _07513_/B vssd1 vssd1 vccd1 vccd1 _11959_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11889_ _11889_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__and2_1
XANTENNA__11481__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ _11232_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _10909_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07080_ _07079_/B _07079_/C _07079_/A vssd1 vssd1 vccd1 vccd1 _07081_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__A2 _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout129 _06947_/X vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__buf_6
Xfanout118 _12704_/A vssd1 vssd1 vccd1 vccd1 _11295_/B2 sky130_fd_sc_hd__buf_6
X_07982_ _07982_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _07984_/B sky130_fd_sc_hd__xor2_1
Xfanout107 _07119_/X vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06933_ _06960_/A _07278_/A _07304_/A _07303_/B _07303_/A vssd1 vssd1 vccd1 vccd1
+ _06963_/B sky130_fd_sc_hd__o41a_4
X_09721_ fanout71/X fanout42/X _07239_/A fanout77/X vssd1 vssd1 vccd1 vccd1 _09722_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06864_ instruction[11] _06868_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
X_09652_ instruction[7] _09650_/Y _09651_/X vssd1 vssd1 vccd1 vccd1 _09652_/X sky130_fd_sc_hd__o21a_1
X_06795_ _06794_/A _06794_/B _11767_/A vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__a21o_1
X_08603_ _08603_/A _08603_/B vssd1 vssd1 vccd1 vccd1 _08616_/C sky130_fd_sc_hd__xor2_1
X_09583_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09583_/X sky130_fd_sc_hd__and2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ _08755_/A fanout83/X _08565_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08535_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08736__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08465_ _08465_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07416_ fanout42/X _12688_/A _07304_/Y _08333_/B vssd1 vssd1 vccd1 vccd1 _07417_/B
+ sky130_fd_sc_hd__o22a_1
X_08396_ _08607_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07347_ _10117_/A _11564_/A fanout38/X _12684_/A vssd1 vssd1 vccd1 vccd1 _07348_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07278_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07278_/Y sky130_fd_sc_hd__xnor2_1
X_09017_ _09017_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06703__B _07289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__buf_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _11983_/A _10321_/C _10053_/B vssd1 vssd1 vccd1 vccd1 _09919_/X sky130_fd_sc_hd__and3_1
X_12930_ _10156_/A _12962_/B2 hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__o21a_1
XANTENNA__10241__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ hold207/X _12885_/A2 _12885_/B1 hold205/X vssd1 vssd1 vccd1 vccd1 hold217/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07903__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11812_ fanout65/X _12029_/B _11812_/C vssd1 vssd1 vccd1 vccd1 _11895_/A sky130_fd_sc_hd__and3b_1
X_12792_ hold37/X hold35/X vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__nand2b_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11743_ _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__xnor2_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07682__A2 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11674_ _11674_/A _11674_/B _11674_/C vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__nor3_1
XANTENNA__11072__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ fanout76/X fanout50/X _07988_/B _11663_/A vssd1 vssd1 vccd1 vccd1 _10626_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09959__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _10557_/A _10557_/B _10557_/C vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08631__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _10488_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10663_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06613__B _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ reg1_val[28] reg1_val[29] _12226_/C vssd1 vssd1 vccd1 vccd1 _12269_/B sky130_fd_sc_hd__and3_1
X_12157_ _12157_/A _12157_/B _12155_/X vssd1 vssd1 vccd1 vccd1 _12158_/B sky130_fd_sc_hd__or3b_1
XANTENNA__08395__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10741__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__xnor2_1
X_12088_ _12141_/A fanout9/A fanout3/X fanout44/X vssd1 vssd1 vccd1 vccd1 _12089_/B
+ sky130_fd_sc_hd__o22a_1
X_11039_ hold273/A _12000_/A2 _11137_/B _11038_/Y _12313_/A1 vssd1 vssd1 vccd1 vccd1
+ _11039_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07370__B2 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07370__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ instruction[39] _06637_/B vssd1 vssd1 vccd1 vccd1 _12571_/B sky130_fd_sc_hd__and2_4
XFILLER_0_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12246__A2 fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ _08369_/A _08369_/B _08206_/Y vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ _07335_/A _07335_/B _07335_/C vssd1 vssd1 vccd1 vccd1 _07336_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08182_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07132_ _07132_/A _07132_/B _07132_/C _07132_/D vssd1 vssd1 vccd1 vccd1 _07138_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__A2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07063_ _08274_/A reg1_val[1] vssd1 vssd1 vccd1 vccd1 _07063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09178__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08386__B1 _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07965_ _07965_/A _07965_/B _07965_/C vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__and3_1
XANTENNA__08138__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ reg1_val[10] _06993_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _06917_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08689__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11142__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _10201_/S _09162_/X _09634_/Y vssd1 vssd1 vccd1 vccd1 _09635_/Y sky130_fd_sc_hd__a21oi_1
X_07896_ _07896_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08689__B2 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ _06850_/B _06863_/A vssd1 vssd1 vccd1 vccd1 _06847_/X sky130_fd_sc_hd__and2_4
X_06778_ _06777_/A _06777_/B _10570_/A vssd1 vssd1 vccd1 vccd1 _10689_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__12237__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_93_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09497_ _09501_/A _09497_/B vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07113__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _08841_/B _08517_/B vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11996__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07113__B2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _08714_/A _08448_/B vssd1 vssd1 vccd1 vccd1 _08500_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12716__A _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ _08755_/A fanout79/X _08430_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08380_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _11739_/A fanout37/X _08233_/B fanout64/X vssd1 vssd1 vccd1 vccd1 _10411_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07416__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11390_ _11390_/A _11390_/B _11390_/C vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ _10337_/Y _10340_/Y _12302_/A vssd1 vssd1 vccd1 vccd1 _10341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13060_ hold283/A _13059_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09169__A2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10272_ _10273_/A _10273_/B vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__nor2_1
X_12011_ curr_PC[25] _12079_/C vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__or2_1
XANTENNA__08377__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ hold144/X _12662_/A _13112_/B hold119/X _13121_/A vssd1 vssd1 vccd1 vccd1
+ hold145/A sky130_fd_sc_hd__o221a_1
XANTENNA__09341__A2 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ _13071_/A hold240/X vssd1 vssd1 vccd1 vccd1 _13163_/D sky130_fd_sc_hd__and2_1
XFILLER_0_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775_ hold74/X hold289/X vssd1 vssd1 vccd1 vccd1 _12775_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07280__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06608__B _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__xnor2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11440__A2_N _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09919__B _10321_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11588_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11590_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ fanout82/X fanout9/X fanout3/X _08565_/B vssd1 vssd1 vccd1 vccd1 _10609_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10539_ _10539_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09935__A _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10962__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ _13260_/CLK hold135/X vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13254_/CLK hold176/X vssd1 vssd1 vccd1 vccd1 _13189_/Q sky130_fd_sc_hd__dfxtp_1
X_12209_ _12253_/B _12209_/B vssd1 vssd1 vccd1 vccd1 _12211_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08907__A2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07750_/X sky130_fd_sc_hd__xor2_1
XANTENNA__07591__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ _06763_/B _06646_/A _12546_/B _06700_/X vssd1 vssd1 vccd1 vccd1 _06931_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09868__B1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08540__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06632_ _06980_/A vssd1 vssd1 vccd1 vccd1 _07002_/A sky130_fd_sc_hd__inv_2
XANTENNA__08286__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09420_ _09420_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09420_/Y sky130_fd_sc_hd__nor2_1
X_06563_ reg2_val[25] _06754_/B _06540_/Y _06562_/Y vssd1 vssd1 vccd1 vccd1 _07059_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09351_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08302_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__or2_1
X_09282_ _09282_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08233_ _08755_/A _08233_/B _08309_/B vssd1 vssd1 vccd1 vccd1 _08233_/X sky130_fd_sc_hd__or3_1
XFILLER_0_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06854__B1 _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout130_A _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08164_ _08164_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ _10920_/A _07091_/B _07091_/C _12600_/B _07128_/A vssd1 vssd1 vccd1 vccd1
+ _07284_/B sky130_fd_sc_hd__o41a_4
X_08095_ _11068_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07046_ _09423_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07082_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08071__A2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08997_ _09043_/A _09043_/B _08367_/A vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__a21oi_1
X_07948_ _09568_/A fanout37/X _08233_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _07949_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09580__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _07879_/A _07879_/B vssd1 vssd1 vccd1 vccd1 _07902_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _10320_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _09917_/B sky130_fd_sc_hd__or2_1
X_10890_ _10890_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ _09549_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09550_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _12560_/A _12568_/A vssd1 vssd1 vccd1 vccd1 _12562_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _12491_/A _12491_/B vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11511_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11442_ hold298/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__or2_1
XANTENNA__13041__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10929__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ fanout55/X fanout13/X fanout47/X fanout63/X vssd1 vssd1 vccd1 vccd1 _11374_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11197__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ hold100/X _13112_/B vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08062__A2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _10319_/X _10322_/Y _10323_/Y vssd1 vssd1 vccd1 vccd1 _10324_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06612__A3 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12697__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ _13085_/A hold254/X vssd1 vssd1 vccd1 vccd1 _13239_/D sky130_fd_sc_hd__and2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10256_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10255_/X sky130_fd_sc_hd__and2b_1
X_10186_ _10447_/B _10184_/X _10185_/Y vssd1 vssd1 vccd1 vccd1 _10186_/Y sky130_fd_sc_hd__a21oi_1
Xfanout290 _13085_/A vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ hold275/X hold49/X vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ hold267/X hold66/X vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__nand2b_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08825__A1 _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12689_ hold11/X _12692_/B _12688_/Y _13013_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XFILLER_0_72_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _11683_/Y _11684_/X _11685_/X _11686_/Y _11708_/X vssd1 vssd1 vccd1 vccd1
+ _11709_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10935__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10396__B1 _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12137__A1 _06890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07800__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08924_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07185__A _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _08267_/A _08267_/B _08850_/X vssd1 vssd1 vccd1 vccd1 _08851_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__09553__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _07855_/B _11955_/A _07855_/A vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__mux2_1
X_08782_ _08755_/A _08782_/A2 _08798_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08783_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ _07825_/A _07825_/B vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__nor2_1
X_07664_ _07664_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06615_ _06613_/Y _06540_/Y _06754_/B reg2_val[21] vssd1 vssd1 vccd1 vccd1 _06987_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_09403_ _10607_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _09405_/B sky130_fd_sc_hd__xnor2_2
X_07595_ _07595_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09334_ hold189/A _12190_/B _13160_/Q vssd1 vssd1 vccd1 vccd1 _09334_/Y sky130_fd_sc_hd__a21oi_1
X_06546_ _12297_/A vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09265_ _09266_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10623__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08216_ _08306_/A _08306_/B _08212_/Y vssd1 vssd1 vccd1 vccd1 _08229_/A sky130_fd_sc_hd__o21ba_1
X_09196_ _08914_/A _08913_/B _08913_/A vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__and2_1
XFILLER_0_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07252__B1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _08078_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07029_ _07059_/A _07029_/B vssd1 vssd1 vccd1 vccd1 _07065_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12679__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__B _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _09903_/A _09903_/B _09901_/Y vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__09544__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _11991_/Y sky130_fd_sc_hd__nor2_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12300__A1 _12299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ curr_PC[13] _11051_/C _11153_/A vssd1 vssd1 vccd1 vccd1 _10942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _10873_/A _10873_/B vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__and2_1
XFILLER_0_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08807__A1 _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__B2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ _12604_/Y _12608_/B _12606_/B vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12543_ _12548_/B _12550_/A vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__nand2_2
XANTENNA__07491__B1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11080__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _12466_/B _12471_/B _12464_/X vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 curr_PC[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _11424_/A _11424_/B _09061_/X vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__a21oi_1
X_11356_ hold298/A _11623_/B _11442_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10307_ _10308_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__nand2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ hold259/X _13025_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06621__B _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11287_ _11399_/A _11287_/B vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__nor2_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _11458_/A _10238_/B vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__xnor2_1
X_10169_ _10028_/A _10028_/B _10026_/Y vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07380_ _07380_/A _07380_/B vssd1 vssd1 vccd1 vccd1 _07381_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _11914_/B _11914_/C vssd1 vssd1 vccd1 vccd1 _11983_/C sky130_fd_sc_hd__or2_1
XANTENNA__12086__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ _08022_/A _08160_/A _08022_/C vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07908__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ _11135_/S _09951_/Y _09168_/A vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08730__C _08730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _08903_/A _08903_/B _08903_/C vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout295_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _11883_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__xnor2_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08724_/X _08835_/B _08706_/X vssd1 vssd1 vccd1 vccd1 _08834_/Y sky130_fd_sc_hd__a21oi_1
X_08765_ _08765_/A _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__or3_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _07916_/A _07716_/B vssd1 vssd1 vccd1 vccd1 _07718_/C sky130_fd_sc_hd__xnor2_1
X_08696_ _08696_/A _08696_/B vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07647_ _07203_/A _07203_/B _07206_/A vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ _09237_/A fanout8/X fanout6/X _08936_/A vssd1 vssd1 vccd1 vccd1 _07579_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06529_ instruction[0] instruction[1] _06850_/B pred_val vssd1 vssd1 vccd1 vccd1
+ _06529_/X sky130_fd_sc_hd__o31a_1
XANTENNA__12708__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _09161_/Y _09316_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09462__A1 _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _09444_/B _09248_/B vssd1 vssd1 vccd1 vccd1 _09266_/A sky130_fd_sc_hd__and2_1
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09179_ _11883_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09183_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09214__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ hold233/A _12190_/B _12275_/C vssd1 vssd1 vccd1 vccd1 _12190_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12140__A1_N _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _11086_/A _11086_/B _11085_/A vssd1 vssd1 vccd1 vccd1 _11212_/C sky130_fd_sc_hd__o21a_1
X_11141_ _11620_/B _11249_/B hold218/A vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07528__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _11072_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07528__B2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _10024_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11875__A3 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11974_ _11974_/A _11974_/B vssd1 vssd1 vccd1 vccd1 _11976_/C sky130_fd_sc_hd__nor2_1
X_10925_ _09473_/Y _10924_/X _11135_/S vssd1 vssd1 vccd1 vccd1 _10925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10835__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10835__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08384__A _08384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ _10856_/A _10948_/B _10856_/C vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__and3_1
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ _10787_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12526_ reg1_val[6] _12527_/B vssd1 vssd1 vccd1 vccd1 _12526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ _12458_/B vssd1 vssd1 vccd1 vccd1 _12457_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09205__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09205__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11408_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__or2_1
XFILLER_0_1_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12388_ _12389_/A _12389_/B _12389_/C vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06632__A _06980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _11339_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11339_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07231__A3 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A2 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ instruction[18] _06850_/Y _06879_/X _06637_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__o211a_4
X_13009_ _12769_/X _13009_/B vssd1 vssd1 vccd1 vccd1 _13010_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11079__A1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__B2 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ _08560_/A _08560_/B _08537_/X vssd1 vssd1 vccd1 vccd1 _08558_/B sky130_fd_sc_hd__a21oi_1
X_07501_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _07536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08481_ _08741_/A _08481_/B vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__xnor2_1
X_07432_ _07521_/A _07521_/B vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11713__A _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12028__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ _11955_/A _07363_/B vssd1 vssd1 vccd1 vccd1 _07364_/C sky130_fd_sc_hd__xor2_2
X_09102_ _09100_/X _09101_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11787__C1 _11786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ _07294_/A _07294_/B vssd1 vssd1 vccd1 vccd1 _07380_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09995__A2 _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout210_A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _11122_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07207__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__B1 _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09935_ _10924_/S _09935_/B vssd1 vssd1 vccd1 vccd1 _09935_/Y sky130_fd_sc_hd__nor2_1
X_09866_ _10481_/A fanout63/X fanout60/X _07000_/A vssd1 vssd1 vccd1 vccd1 _09867_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07373__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _08821_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__or2_1
XANTENNA__09380__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _09638_/X _09639_/Y _09641_/Y vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__o21a_1
X_08748_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _09005_/A sky130_fd_sc_hd__xnor2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08680_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__and2b_1
X_10710_ hold261/A _12304_/B1 _10820_/B _10709_/Y _09810_/A vssd1 vssd1 vccd1 vccd1
+ _10710_/X sky130_fd_sc_hd__a311o_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11689_/A _11689_/B _11689_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11708_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11778__C1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__A _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10641_ _11068_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _12297_/A _09141_/Y _12310_/X vssd1 vssd1 vccd1 vccd1 _12311_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11793__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _10450_/A _12217_/X _12218_/Y _12241_/X vssd1 vssd1 vccd1 vccd1 _12242_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _12263_/S _12173_/B vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__and2_1
XANTENNA__07267__B _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11124_ _11124_/A _11124_/B _11124_/C vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or3_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11055_ _11799_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__xnor2_1
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10014_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _12023_/A _11957_/B vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11481__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _10449_/C _11230_/A _11231_/B _11230_/B vssd1 vssd1 vccd1 vccd1 _10909_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11888_ _11889_/A _11889_/B vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11481__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ _10840_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ _12509_/A _12509_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xor2_4
XANTENNA__12364__A _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11536__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07981_ _07981_/A _07981_/B vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__xor2_2
Xfanout108 _11955_/A vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__buf_12
Xfanout119 _12704_/A vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06932_ _07137_/A _07109_/A _06932_/C _06942_/C vssd1 vssd1 vccd1 vccd1 _07303_/B
+ sky130_fd_sc_hd__or4_2
X_09720_ _09720_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__xor2_1
X_06863_ _06863_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _06868_/B sky130_fd_sc_hd__or2_2
X_09651_ _12263_/S _09651_/B _09651_/C vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__or3_1
X_06794_ _06794_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06794_/X sky130_fd_sc_hd__and2_1
X_08602_ _08638_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__nor2_1
X_09582_ _11796_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07921__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08533_ _08533_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _08563_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout160_A _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _06848_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07676__B1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08464_ _08464_/A _08464_/B _08464_/C vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__or3_1
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12973__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07415_ _07415_/A _07415_/B vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08395_ _08606_/A2 _08733_/B1 _08735_/A2 _08642_/B vssd1 vssd1 vccd1 vccd1 _08396_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _09979_/A _07346_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07277_/X sky130_fd_sc_hd__xor2_4
X_09016_ _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10506__B _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _11983_/A _10053_/B _10321_/C vssd1 vssd1 vccd1 vccd1 _09918_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09353__B1 _09350_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout73_A _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09704_/A _09704_/B _09702_/Y vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__a21oi_4
X_12860_ _13062_/A hold208/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__and2_1
XANTENNA__09105__A0 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11883_/A _11811_/B vssd1 vssd1 vccd1 vccd1 _11812_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08927__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ _12791_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__nor2_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ _11666_/A _11666_/B _11664_/Y vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11463__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11674_/A _11674_/B _11674_/C vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10624_ _12086_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09959__A2 _09955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _10555_/A _10555_/B vssd1 vssd1 vccd1 vccd1 _10557_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08631__A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12176__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07278__A _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10419_/A _10419_/B _10416_/A vssd1 vssd1 vccd1 vccd1 _10488_/B sky130_fd_sc_hd__a21oi_1
X_12225_ _12225_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12191__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12157_/A _12157_/B _12155_/X vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__08395__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__nand2b_1
X_12087_ _12146_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__and2_1
X_11038_ _12000_/A2 _11137_/B hold273/A vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07370__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ _12777_/X _12989_/B vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07200_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07335_/C sky130_fd_sc_hd__xnor2_1
X_08180_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__and2_1
XANTENNA__12954__A1 _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07131_ _07132_/C _07132_/D vssd1 vssd1 vccd1 vccd1 _07131_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10607__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07062_ _12499_/A _12501_/A vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07916__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A1 _08387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12541__B _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08138__A1 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12968__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07895_ _07896_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__or2_1
X_06915_ _10920_/A _06915_/B vssd1 vssd1 vccd1 vccd1 _06915_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08138__B2 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09704_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11157__B _11157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
X_06846_ instruction[5] _06846_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xor2_4
XFILLER_0_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06777_ _06777_/A _06777_/B vssd1 vssd1 vccd1 vccd1 _06777_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11173__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09565_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09496_ _12263_/S _09494_/Y _09495_/X vssd1 vssd1 vccd1 vccd1 _09497_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07113__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _08516_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08447_ _08670_/A2 _08735_/A2 _08735_/B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08448_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08378_ _08535_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07329_ _07330_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07649_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _11135_/S _10217_/X _10339_/X vssd1 vssd1 vccd1 vccd1 _10340_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__07098__A _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10273_/B sky130_fd_sc_hd__xnor2_1
X_12010_ _11980_/X _11981_/Y _11984_/Y _09145_/Y _12009_/Y vssd1 vssd1 vccd1 vccd1
+ _12010_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08377__A1 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__A1 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12912_ _07010_/B _12686_/B hold149/X vssd1 vssd1 vccd1 vccd1 _13197_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12843_ hold194/X _12885_/A2 _12885_/B1 hold239/X vssd1 vssd1 vccd1 vccd1 hold240/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12179__A _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ hold300/A hold27/X vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__nand2b_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ fanout17/X fanout13/X _07156_/X fanout9/A vssd1 vssd1 vccd1 vccd1 _11726_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11811__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12936__A1 _07301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout90 _12688_/A vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__buf_4
X_11656_ _11656_/A _11656_/B vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11674_/B sky130_fd_sc_hd__and2b_1
X_10607_ _10607_/A _10607_/B vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10538_ _10538_/A _10538_/B vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13257_ _13260_/CLK hold178/X vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10469_ hold279/A hold300/A _10469_/C vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__or3_2
XFILLER_0_110_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06672__A_N _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _12208_/A _12208_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12209_/B sky130_fd_sc_hd__nand3_1
X_13188_ _13188_/CLK _13188_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ _12080_/A _12082_/X _12113_/X _12138_/X vssd1 vssd1 vccd1 vccd1 dest_val[27]
+ sky130_fd_sc_hd__o22a_4
XANTENNA__07591__A2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ reg2_val[9] _06700_/B vssd1 vssd1 vccd1 vccd1 _06700_/X sky130_fd_sc_hd__and2_1
XANTENNA__09868__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07680_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07695_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08540__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ reg2_val[19] _06748_/B _06657_/B1 _06630_/X vssd1 vssd1 vccd1 vccd1 _06980_/A
+ sky130_fd_sc_hd__a22o_2
XANTENNA__12089__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08540__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ _06613_/A _12546_/B vssd1 vssd1 vccd1 vccd1 _06562_/Y sky130_fd_sc_hd__nor2_1
X_09350_ _09288_/X _09293_/Y _09349_/X _12080_/A vssd1 vssd1 vccd1 vccd1 _09350_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__xor2_4
X_08301_ _08535_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08354_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _11072_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09398__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__B _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08163_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _08202_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout123_A _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07114_ _12085_/A _07114_/B vssd1 vssd1 vccd1 vccd1 _07142_/A sky130_fd_sc_hd__xnor2_1
X_08094_ _08755_/A fanout37/X _08233_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08095_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ _12720_/A _09422_/A _09222_/B2 _12094_/A vssd1 vssd1 vccd1 vccd1 _07046_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11363__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08996_ _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__xor2_2
X_07947_ _07959_/B _07947_/B vssd1 vssd1 vccd1 vccd1 _07953_/B sky130_fd_sc_hd__nor2_2
XANTENNA__09861__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09072__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _07930_/A _07930_/B _07963_/B _07877_/B _07877_/A vssd1 vssd1 vccd1 vccd1
+ _07902_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_97_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06829_ _08823_/B _06829_/B vssd1 vssd1 vccd1 vccd1 _06833_/D sky130_fd_sc_hd__nand2_1
X_09617_ _09464_/A _09617_/B _09617_/C vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ _09547_/B _09547_/C _09547_/A vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08295__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout36_A fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _09086_/X _09090_/X _09479_/S vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _11509_/A _11509_/B _11547_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__o21ai_1
X_12490_ _12496_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12918__A1 _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _09120_/S _10925_/X _10938_/Y _09330_/A _11440_/X vssd1 vssd1 vccd1 vccd1
+ _11450_/A sky130_fd_sc_hd__o221a_1
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _11372_/A _11372_/B vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__xnor2_1
X_13111_ _13111_/A hold127/X vssd1 vssd1 vccd1 vccd1 _13254_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10323_ _10319_/X _10322_/Y _10450_/A vssd1 vssd1 vccd1 vccd1 _10323_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13042_ hold253/X _13084_/A2 _13041_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold254/A
+ sky130_fd_sc_hd__a22o_1
X_10254_ _10254_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10185_ _10447_/B _10184_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _10185_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11078__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout291 fanout298/X vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__clkbuf_4
Xfanout280 _06530_/X vssd1 vssd1 vccd1 vccd1 _06665_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__08387__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ _13090_/B _13091_/A _12738_/X vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12757_ hold66/X hold267/X vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__and2b_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12688_ _12688_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _12688_/Y sky130_fd_sc_hd__nand2_1
X_11708_ _11708_/A _11708_/B _11708_/C _11700_/X vssd1 vssd1 vccd1 vccd1 _11708_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_72_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11639_ fanout65/X fanout8/X fanout6/X fanout68/X vssd1 vssd1 vccd1 vccd1 _11640_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09250__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12372__A _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08210__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _08267_/A _08267_/B _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08850_/X
+ sky130_fd_sc_hd__a211o_1
X_07801_ _07916_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07855_/B sky130_fd_sc_hd__xnor2_1
X_08781_ _08771_/C _08771_/B _08770_/Y vssd1 vssd1 vccd1 vccd1 _08784_/B sky130_fd_sc_hd__a21bo_1
X_07732_ _07732_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07825_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11716__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06614_ reg2_val[21] _06754_/B _06540_/Y _06613_/Y vssd1 vssd1 vccd1 vccd1 _07012_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_09402_ _10481_/A fanout64/X fanout58/X _07000_/A vssd1 vssd1 vccd1 vccd1 _09403_/B
+ sky130_fd_sc_hd__o22a_1
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09333_/Y sky130_fd_sc_hd__xnor2_1
X_07594_ _07594_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12073__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06545_ _06545_/A _06545_/B vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__or2_4
XANTENNA__08277__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10084__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09264_ _09264_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09266_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10623__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _08535_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__xnor2_1
X_09195_ _08956_/A _08956_/B _08953_/A vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ _08146_/A _08146_/B vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07252__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__B2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _08077_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08078_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12128__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ _07028_/A _07028_/B _07028_/C _07028_/D vssd1 vssd1 vccd1 vccd1 _07065_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11336__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _07658_/A _07658_/B _07656_/X vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__a21oi_4
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _11924_/A _11921_/Y _11923_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__o21a_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11639__B2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _12179_/A _10912_/X _10913_/Y _10940_/X _10911_/Y vssd1 vssd1 vccd1 vccd1
+ _10941_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12611_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _12620_/C sky130_fd_sc_hd__nand2_2
X_10872_ _10873_/A _10873_/B vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12064__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__A2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ reg1_val[9] _12542_/B vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _12496_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12478_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__07491__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 curr_PC[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11623_/B _11442_/B hold298/A vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07286__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ _11286_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11287_/B sky130_fd_sc_hd__nor2_1
X_10306_ _10443_/B _10306_/B vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__and2_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13025_ _13025_/A _13025_/B vssd1 vssd1 vccd1 vccd1 _13025_/Y sky130_fd_sc_hd__xnor2_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ fanout8/A _07763_/B fanout6/X _10370_/A vssd1 vssd1 vccd1 vccd1 _10238_/B
+ sky130_fd_sc_hd__o22a_1
X_10168_ _10168_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__nand2_1
X_10099_ _10099_/A1 fanout51/X _07988_/B _10359_/B2 vssd1 vssd1 vccd1 vccd1 _10100_/B
+ sky130_fd_sc_hd__o22a_1
X_12809_ _13044_/B _13045_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _13050_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11271__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ _08159_/A _08159_/B _07999_/Y vssd1 vssd1 vccd1 vccd1 _08022_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09676__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09951_ _11033_/A _09486_/X _09166_/B vssd1 vssd1 vccd1 vccd1 _09951_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08902_ _08903_/A _08903_/B _08903_/C vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _12684_/A _07183_/A _07183_/B fanout45/X _10370_/A vssd1 vssd1 vccd1 vccd1
+ _09883_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_57_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _09005_/A _09005_/B _08747_/X vssd1 vssd1 vccd1 vccd1 _09004_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout288_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06760__A3 _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07715_ _09568_/A fanout49/X _09428_/A fanout51/X vssd1 vssd1 vccd1 vccd1 _07716_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07135__S _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08695_ _08693_/A _08693_/B _08694_/Y vssd1 vssd1 vccd1 vccd1 _08696_/B sky130_fd_sc_hd__o21a_1
X_07646_ _07404_/A _07404_/B _07402_/Y vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08755__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ _07268_/A _12245_/A _12029_/B vssd1 vssd1 vccd1 vccd1 fanout6/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11254__C1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06528_ reg2_val[31] _06700_/B vssd1 vssd1 vccd1 vccd1 _06528_/X sky130_fd_sc_hd__and2_1
X_09316_ _09114_/X _09116_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10057__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _09444_/A _09246_/C _09246_/A vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _09698_/A _12141_/A fanout45/X _09885_/A vssd1 vssd1 vccd1 vccd1 _09179_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11557__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09586__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08129_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ hold171/A _11140_/B vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07528__A2 _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ fanout43/X fanout9/X fanout3/X _08333_/B vssd1 vssd1 vccd1 vccd1 _11072_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07834__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12285__A1 _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _11973_/A _11973_/B _11973_/C vssd1 vssd1 vccd1 vccd1 _11974_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10924_ _09934_/Y _09938_/Y _10924_/S vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10835__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _10855_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _10856_/C sky130_fd_sc_hd__or2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__A _11091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12524_/A _12521_/Y _12523_/B vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__o21a_2
X_10786_ _10787_/B _10787_/A vssd1 vssd1 vccd1 vccd1 _10904_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ _12478_/A _12480_/A vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09205__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ _12396_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12389_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _11407_/A _11407_/B vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _06785_/Y _11337_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13253_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__09508__A3 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _11654_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__xor2_1
X_13008_ _13013_/A hold256/X vssd1 vssd1 vccd1 vccd1 _13232_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07500_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07501_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11079__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _08755_/B _08715_/A2 _08735_/B1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 _08481_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07431_ _08916_/A _07431_/B vssd1 vssd1 vccd1 vccd1 _07521_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12028__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12028__B2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ _07099_/X _07154_/X _07799_/B _07110_/Y vssd1 vssd1 vccd1 vccd1 _07363_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ reg1_val[11] reg1_val[20] _09120_/S vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07455__A1 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07455__B2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07293_ _07875_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07294_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__A3 _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07919__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ _08587_/X _09032_/B vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__and2b_1
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07207__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__A1 _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10762__B2 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ _10201_/S _09303_/X _09933_/Y vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__o21ai_1
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__xor2_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _09423_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09380__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _11696_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__nand2_1
X_08747_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08747_/X sky130_fd_sc_hd__and2b_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10278__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _11068_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__xnor2_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08891__B1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ _11876_/A fanout37/X _08233_/B _11950_/A vssd1 vssd1 vccd1 vccd1 _10641_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _10570_/A _10570_/B _10570_/Y _09498_/A vssd1 vssd1 vccd1 vccd1 _10571_/X
+ sky130_fd_sc_hd__a211o_1
X_12310_ reg1_val[31] _07184_/B _09147_/X _12309_/X _12280_/A vssd1 vssd1 vccd1 vccd1
+ _12310_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _09145_/Y _12225_/Y _12240_/X _12222_/X vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _06559_/Y _12114_/X _06560_/A vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11123_ _11232_/A _11122_/B _11122_/C vssd1 vssd1 vccd1 vccd1 _11123_/Y sky130_fd_sc_hd__o21ai_1
X_11054_ _11739_/A fanout13/X fanout47/X fanout64/X vssd1 vssd1 vccd1 vccd1 _11055_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10005_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07382__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11956_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__and2_1
XFILLER_0_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10907_ _11014_/B _10907_/B vssd1 vssd1 vccd1 vccd1 _11230_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11887_ _11887_/A _11887_/B vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11481__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838_ _11799_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10840_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ _10770_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10894_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _12506_/Y _12508_/B vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_124_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12439_ _12439_/A _12439_/B vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06948__B1 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _07980_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__nor2_1
Xfanout109 _11955_/A vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__clkbuf_8
X_06931_ _07296_/A _06931_/B vssd1 vssd1 vccd1 vccd1 _06942_/C sky130_fd_sc_hd__or2_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ reg1_val[2] _09634_/A _09649_/X vssd1 vssd1 vccd1 vccd1 _09650_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06862_ instruction[13] _06862_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
X_08601_ _08601_/A _08601_/B vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__xnor2_1
X_06793_ _06792_/A _06792_/B _11689_/A vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__a21o_1
X_09581_ _10377_/A1 fanout49/X fanout92/X fanout50/X vssd1 vssd1 vccd1 vccd1 _09582_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08532_ _08533_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _08532_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07676__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08463_ _08514_/A _08462_/B _08459_/X vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__a21o_1
X_07414_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07415_/B sky130_fd_sc_hd__and2_1
XANTENNA__07676__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08394_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07345_ _07238_/Y fanout92/X _12690_/A fanout42/X vssd1 vssd1 vccd1 vccd1 _07346_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ _07276_/A _07276_/B vssd1 vssd1 vccd1 vccd1 _07332_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09015_ _09015_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _09621_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B2 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__A _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07600__B2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07600__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _10321_/A _09917_/B _10320_/B vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__or3_1
XANTENNA__09353__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__xnor2_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07903__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _10320_/B _09778_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _09779_/Y sky130_fd_sc_hd__o21ai_1
X_12790_ hold249/A hold53/X vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__and2b_1
X_11810_ fanout63/X fanout11/X fanout44/X _12094_/A vssd1 vssd1 vccd1 vccd1 _11811_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A _11741_/B vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__xnor2_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11463__A2 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11674_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10623_ _11169_/A fanout14/X fanout52/X _11297_/A vssd1 vssd1 vccd1 vccd1 _10624_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13060__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10554_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10555_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10485_ _10663_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10488_/A sky130_fd_sc_hd__or2_1
X_12224_ _12223_/A _12223_/B _12223_/C vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12155_ _12155_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _12155_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11809__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11108_/B sky130_fd_sc_hd__xnor2_1
X_12086_ _12086_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__nand2_1
X_11037_ hold297/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11137_/B sky130_fd_sc_hd__or2_1
XANTENNA__07355__B1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ _13103_/A hold286/X vssd1 vssd1 vccd1 vccd1 _13228_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07107__B1 _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11939_ _11918_/Y _11919_/X _11926_/X _11938_/X vssd1 vssd1 vccd1 vccd1 _11939_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07130_ reg1_val[22] _07284_/B _07130_/C vssd1 vssd1 vccd1 vccd1 _07132_/D sky130_fd_sc_hd__nor3_1
XANTENNA__08083__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12094__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__B2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07061_ _09862_/B _07061_/B vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _07963_/A _07963_/B vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08138__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07894_ _07892_/A _07892_/B _07893_/X vssd1 vssd1 vccd1 vccd1 _07896_/B sky130_fd_sc_hd__a21oi_1
X_06914_ _10920_/A _06915_/B vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__xor2_4
X_09702_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09702_/Y sky130_fd_sc_hd__nor2_1
X_09633_ _09316_/X _09318_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09623__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ instruction[3] _06825_/X _06839_/X _06843_/Y _06841_/X vssd1 vssd1 vccd1
+ vccd1 _06846_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__xnor2_2
X_06776_ _06775_/A _06775_/B _06830_/C vssd1 vssd1 vccd1 vccd1 _06777_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08515_ _08516_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__nand2_1
X_09495_ _09495_/A _09495_/B _09495_/C vssd1 vssd1 vccd1 vccd1 _09495_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ _08741_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09859__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08377_ _08565_/B _08737_/A2 _08813_/B1 fanout83/X vssd1 vssd1 vccd1 vccd1 _08378_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07328_ _07649_/A _07328_/B vssd1 vssd1 vccd1 vccd1 _07330_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_46_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07259_ _07259_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08377__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08003__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ hold146/X _12662_/A _13112_/B hold144/X _13013_/A vssd1 vssd1 vccd1 vccd1
+ hold149/A sky130_fd_sc_hd__o221a_1
XANTENNA__07842__A _07842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _13071_/A hold195/X vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__and2_1
XFILLER_0_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12773_ hold27/X hold300/A vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__and2b_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11724_ _11724_/A _11724_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08673__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ fanout51/X fanout9/A fanout3/X _07138_/Y vssd1 vssd1 vccd1 vccd1 _11656_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07289__A _07289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout80 fanout81/X vssd1 vssd1 vccd1 vccd1 fanout80/X sky130_fd_sc_hd__buf_6
Xfanout91 _07296_/Y vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ _11674_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11588_/B sky130_fd_sc_hd__nor2_1
X_10606_ _10607_/A _10607_/B vssd1 vssd1 vccd1 vccd1 _10606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10537_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10538_/B sky130_fd_sc_hd__nor3_1
X_13256_ _13260_/CLK hold165/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__dfxtp_1
X_10468_ _06706_/B _09141_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _10468_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12208_/A _12208_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06921__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _13188_/CLK _13187_/D vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__dfxtp_1
X_10399_ _10399_/A _10399_/B vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__nor2_1
X_12138_ _12265_/C1 _12117_/Y _12119_/X _12137_/Y vssd1 vssd1 vccd1 vccd1 _12138_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13113__A2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ hold235/A _12190_/B _12129_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12069_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09868__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__C1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _06646_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _06630_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06561_ instruction[35] _06637_/B vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__and2_4
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09280_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09280_/X sky130_fd_sc_hd__and2_1
X_08300_ fanout83/X _08733_/B1 _08735_/A2 _08565_/B vssd1 vssd1 vccd1 vccd1 _08301_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09679__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08231_ _09237_/A fanout43/X _08333_/B _09428_/A vssd1 vssd1 vccd1 vccd1 _08232_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07113_ _09568_/A fanout15/X _09698_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _07114_/B
+ sky130_fd_sc_hd__o22a_1
X_08093_ _08093_/A _08093_/B vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11060__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _07044_/A _07044_/B vssd1 vssd1 vccd1 vccd1 _07044_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12552__B _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11363__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__C1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__xnor2_1
X_07946_ _07946_/A _07946_/B vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__and2_1
XANTENNA__07319__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__B1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _07877_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11184__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ _06828_/A _12668_/A vssd1 vssd1 vccd1 vccd1 _06829_/B sky130_fd_sc_hd__nand2_1
X_09616_ _09616_/A _09616_/B vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__xnor2_4
X_06759_ _06753_/B _06537_/Y _12507_/B _06754_/X reg1_val[1] vssd1 vssd1 vccd1 vccd1
+ _06759_/Y sky130_fd_sc_hd__a311oi_2
X_09547_ _09547_/A _09547_/B _09547_/C vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__and3_1
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08295__A1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _09083_/X _09109_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09478_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08295__B2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout29_A _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13222_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08429_ _08535_/A _08429_/B vssd1 vssd1 vccd1 vccd1 _08497_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12918__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ reg1_val[18] _06980_/B _09138_/X _11439_/X vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11372_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13110_ hold301/X _13110_/A2 _13109_/X _06858_/B hold126/X vssd1 vssd1 vccd1 vccd1
+ hold127/A sky130_fd_sc_hd__a32o_1
XANTENNA__07837__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _10447_/A _10447_/B _10447_/C _12223_/A vssd1 vssd1 vccd1 vccd1 _10322_/Y
+ sky130_fd_sc_hd__o31ai_1
X_13041_ hold267/A _13040_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12000__C1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _10254_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10374_/A sky130_fd_sc_hd__nand2_1
X_10184_ _10447_/A _10053_/X _10449_/A vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__o21a_1
Xfanout281 _12498_/C vssd1 vssd1 vccd1 vccd1 _06637_/B sky130_fd_sc_hd__buf_4
Xfanout270 _13084_/B2 vssd1 vssd1 vccd1 vccd1 _13070_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout292 _13111_/A vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__buf_4
XANTENNA__08387__B _08387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08522__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ _12742_/B _13086_/B _12740_/X vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__a21o_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12756_ hold253/X hold5/X vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__nand2b_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ hold25/X _12686_/B _12686_/Y _13121_/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__o211a_1
X_11707_ _11702_/Y _11703_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11708_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__06635__B _06980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ _12089_/A _11638_/B vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09786__A1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _11739_/A fanout7/X fanout5/X _11663_/A vssd1 vssd1 vccd1 vccd1 _11649_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ _13241_/CLK _13239_/D vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11269__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07800_ fanout51/X _09237_/A _09428_/A fanout49/X vssd1 vssd1 vccd1 vccd1 _07801_/B
+ sky130_fd_sc_hd__o22a_1
X_08780_ _08784_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08795_/A sky130_fd_sc_hd__xor2_2
X_07731_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07825_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07482__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _07662_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__nand2_1
X_06613_ _06613_/A _12527_/B vssd1 vssd1 vccd1 vccd1 _06613_/Y sky130_fd_sc_hd__nor2_1
X_07593_ _07594_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07593_/Y sky130_fd_sc_hd__nor2_1
X_09401_ _10126_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06544_ reg1_val[31] _07604_/A vssd1 vssd1 vccd1 vccd1 _06545_/B sky130_fd_sc_hd__nor2_1
X_09332_ _08814_/A _12112_/A _09331_/X vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08277__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10608__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08277__B2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _09263_/A _09263_/B vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09202__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13022__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08214_ fanout83/X _08735_/A2 _08735_/B1 _08565_/B vssd1 vssd1 vccd1 vccd1 _08215_/B
+ sky130_fd_sc_hd__o22a_1
X_09194_ _09194_/A _09194_/B vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09226__B1 _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _08154_/B _08154_/A vssd1 vssd1 vccd1 vccd1 _08145_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07252__A2 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ _09423_/A vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__clkinv_8
XFILLER_0_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09083__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ _08978_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__xnor2_4
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _07929_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11639__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10940_ _12303_/A _10926_/X _10939_/X _10918_/X vssd1 vssd1 vccd1 vccd1 _10940_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07712__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ reg1_val[22] _12615_/B vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11642__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _11296_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10873_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12541_ reg1_val[9] _12542_/B vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__or2_1
XANTENNA__11272__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ reg1_val[23] curr_PC[23] _12495_/S vssd1 vssd1 vccd1 vccd1 _12473_/B sky130_fd_sc_hd__mux2_2
XANTENNA__07491__A2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ _11233_/A _12110_/A _11331_/X _11235_/A vssd1 vssd1 vccd1 vccd1 _11424_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 curr_PC[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11354_ hold253/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07286__B _07286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _11286_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__and2_1
X_10305_ _10305_/A _10305_/B _10305_/C vssd1 vssd1 vccd1 vccd1 _10306_/B sky130_fd_sc_hd__or3_1
X_13024_ _12763_/X _13024_/B vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__nand2b_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _10236_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10273_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08398__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _09974_/A _09974_/B _09975_/Y vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10098_ _09994_/A _09993_/B _09991_/X vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07703__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12808_ _13039_/B _13040_/A _12757_/X vssd1 vssd1 vccd1 vccd1 _13045_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12739_ hold265/X hold95/X vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__nand2b_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09950_ _09152_/Y _09944_/Y _09949_/X vssd1 vssd1 vccd1 vccd1 _09950_/Y sky130_fd_sc_hd__a21oi_1
Xmax_cap256 _08276_/A vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__buf_4
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08901_ _08901_/A _08901_/B vssd1 vssd1 vccd1 vccd1 _08903_/C sky130_fd_sc_hd__xor2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _11885_/A _09881_/B vssd1 vssd1 vccd1 vccd1 _09888_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _09006_/A _09006_/B _08761_/X vssd1 vssd1 vccd1 vccd1 _09005_/B sky130_fd_sc_hd__a21o_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08101__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ _08763_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _08772_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07714_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07714_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08694_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08694_/Y sky130_fd_sc_hd__nand2b_1
X_07645_ _07334_/A _07334_/B _07333_/A vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11462__A _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__B _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _11124_/A _07574_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _07576_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06527_ instruction[0] _06850_/B instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06527_/X sky130_fd_sc_hd__or4bb_2
X_09315_ _09314_/X _09311_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__A1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ _09246_/A _09444_/A _09246_/C vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09867__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08670__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09177_ _09194_/B _08925_/B _08934_/B _08935_/B _08935_/A vssd1 vssd1 vccd1 vccd1
+ _09193_/A sky130_fd_sc_hd__a32o_2
XANTENNA__11557__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11557__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _08128_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08059_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08077_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout96_A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _11184_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11073_/A sky130_fd_sc_hd__xnor2_1
X_10021_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__and2_1
XANTENNA__12285__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11974_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10923_ _10923_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10923_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ _10855_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _10948_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11091__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12524_/A _12524_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
X_10785_ _10785_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10787_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ _12455_/A _12455_/B _12455_/C vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__and3_1
XFILLER_0_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06913__B _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11548__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _12546_/B _12386_/B vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _11407_/A _11407_/B vssd1 vssd1 vccd1 vccd1 _11504_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _06662_/B _11237_/Y _06660_/Y vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _12148_/A _11564_/A fanout38/X _12201_/A vssd1 vssd1 vccd1 vccd1 _11269_/B
+ sky130_fd_sc_hd__o22a_1
X_13007_ hold255/X _12663_/B _13006_/X hold177/X vssd1 vssd1 vccd1 vccd1 hold256/A
+ sky130_fd_sc_hd__a22o_1
X_10219_ _12073_/B2 _10204_/Y _10218_/Y _09124_/S _10216_/X vssd1 vssd1 vccd1 vccd1
+ _10219_/X sky130_fd_sc_hd__o221a_1
X_11199_ _11200_/B _11199_/B vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12378__A _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ fanout80/X _06940_/A _10490_/B2 fanout82/X vssd1 vssd1 vccd1 vccd1 _07431_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12028__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09429__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07361_ _07361_/A _07361_/B _07361_/C vssd1 vssd1 vccd1 vccd1 _07364_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09100_ reg1_val[10] reg1_val[21] _09120_/S vssd1 vssd1 vccd1 vccd1 _09100_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07455__A2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07292_ _12684_/A _11564_/A _12686_/A fanout38/X vssd1 vssd1 vccd1 vccd1 _07293_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07207__A2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__A2 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07000__A _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09626__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10762__A2 _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ _09314_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09933_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__nand2_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _09313_/S _08815_/B vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__or2_1
XANTENNA__07915__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _11135_/S _09793_/X _09794_/X vssd1 vssd1 vccd1 vccd1 _09796_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__10278__A1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ _08732_/A _08732_/B _08745_/X vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__o21bai_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11475__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _08655_/A _08655_/B _08676_/Y vssd1 vssd1 vccd1 vccd1 _08680_/A sky130_fd_sc_hd__o21a_1
XANTENNA__10278__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07628_ fanout92/X fanout37/X fanout34/X _12694_/A vssd1 vssd1 vccd1 vccd1 _07629_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08891__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07559_ _07559_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07560_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10570_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10570_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout11_A _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09229_ _09228_/B _09228_/C _09563_/A vssd1 vssd1 vccd1 vccd1 _09231_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ _12240_/A _12240_/B _12240_/C _12236_/X vssd1 vssd1 vccd1 vccd1 _12240_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12112_/A _12258_/C _12169_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _12171_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ _11232_/A _11122_/B _11122_/C vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__or3_1
X_11053_ _11153_/A _11152_/B _11052_/Y _11050_/X vssd1 vssd1 vccd1 vccd1 dest_val[14]
+ sky130_fd_sc_hd__o31ai_4
X_10004_ _09848_/A _09848_/B _09844_/X vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__07382__B2 _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _11955_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11466__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06908__B _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10906_ _11014_/A _10796_/B _10791_/A vssd1 vssd1 vccd1 vccd1 _10907_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ _12201_/A fanout15/X _07513_/B fanout9/A vssd1 vssd1 vccd1 vccd1 _11887_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10837_ fanout76/X fanout13/X fanout47/X _11663_/A vssd1 vssd1 vccd1 vccd1 _10838_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ _10894_/A _10768_/B vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_124_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ reg1_val[2] _12507_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12438_ _12455_/A _12438_/B vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__nand2_1
X_10699_ _10699_/A vssd1 vssd1 vccd1 vccd1 _10699_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06643__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12369_ _12375_/B _12369_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
XANTENNA__06948__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06930_ _07137_/A _07109_/A _06932_/C vssd1 vssd1 vccd1 vccd1 _06930_/X sky130_fd_sc_hd__or3_1
XANTENNA__08570__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ instruction[12] _06862_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
X_08600_ _08741_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__xnor2_1
X_06792_ _06792_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06792_/X sky130_fd_sc_hd__and2_1
X_09580_ _11183_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11457__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _08607_/A _08531_/B vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08462_ _08459_/X _08462_/B vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__nand2b_1
X_07413_ _07540_/A _07412_/Y _07408_/X vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07676__A2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12836__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08393_ _08458_/A _08392_/B _08388_/X vssd1 vssd1 vccd1 vccd1 _08404_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout146_A _07122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12957__B1 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ _07344_/A _07344_/B vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07275_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07276_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12185__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08389__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08928__A2 _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold186 hold203/X vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _10321_/C sky130_fd_sc_hd__xnor2_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _11183_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__xnor2_4
X_09778_ _10321_/A _09917_/B _11983_/A vssd1 vssd1 vccd1 vccd1 _09778_/X sky130_fd_sc_hd__o21a_1
X_08729_ _08729_/A _08752_/A vssd1 vssd1 vccd1 vccd1 _08732_/A sky130_fd_sc_hd__xnor2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11741_/A _11741_/B vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__and2_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10120__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11671_ _11671_/A _11671_/B vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ _10622_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__xnor2_2
X_10553_ _10554_/A _10554_/B vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__and2_1
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10974__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10484_ _10484_/A _10484_/B _10621_/A vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__and3_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ _12223_/A _12223_/B _12223_/C vssd1 vssd1 vccd1 vccd1 _12225_/A sky130_fd_sc_hd__and3_1
X_12154_ _12155_/B _12155_/A vssd1 vssd1 vccd1 vccd1 _12211_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11105_ _11106_/B _11106_/A vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09344__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _12085_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__or2_1
XANTENNA__07355__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _11032_/Y _11035_/Y _11696_/A vssd1 vssd1 vccd1 vccd1 _11036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11439__A0 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ hold285/X _06858_/B _12986_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold286/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06638__B _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__S _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11938_ _11932_/Y _11933_/X _11937_/X _11930_/X vssd1 vssd1 vccd1 vccd1 _11938_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ _11869_/A _11871_/B _11869_/C vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11611__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07060_ _12716_/A _09727_/A _08798_/B _12718_/A vssd1 vssd1 vccd1 vccd1 _07061_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08083__A2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07962_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/A sky130_fd_sc_hd__or2_1
X_09701_ _11885_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07893_ _07972_/B _07972_/A vssd1 vssd1 vccd1 vccd1 _07893_/X sky130_fd_sc_hd__and2b_1
X_06913_ _07128_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _06915_/B sky130_fd_sc_hd__and2_2
XFILLER_0_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ _09631_/X _09630_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09632_/X sky130_fd_sc_hd__mux2_1
X_06844_ _06892_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__or2_2
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09563_ _09563_/A _09563_/B vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06548__B _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ _06775_/A _06775_/B vssd1 vssd1 vccd1 vccd1 _06775_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout263_A _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__xnor2_1
X_09494_ _06761_/A _08823_/B _06759_/Y vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ _08740_/A2 _08715_/A2 _08689_/B1 _08755_/B vssd1 vssd1 vccd1 vccd1 _08446_/B
+ sky130_fd_sc_hd__o22a_1
X_08376_ _08350_/A _08349_/C _08349_/B vssd1 vssd1 vccd1 vccd1 _08376_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11470__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ _07327_/A _07327_/B _07327_/C vssd1 vssd1 vccd1 vccd1 _07328_/B sky130_fd_sc_hd__or3_1
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07258_ _07259_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07189_ _12142_/A _07189_/B vssd1 vssd1 vccd1 vccd1 _07200_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _08688_/A _12686_/B hold147/X vssd1 vssd1 vccd1 vccd1 _13196_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__08534__B1 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ hold247/A _12885_/A2 _12885_/B1 hold194/X vssd1 vssd1 vccd1 vccd1 hold195/A
+ sky130_fd_sc_hd__a22o_1
X_12772_ hold279/A hold25/X vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__nand2b_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11723_ _11723_/A _11723_/B _11723_/C vssd1 vssd1 vccd1 vccd1 _11724_/B sky130_fd_sc_hd__nand3_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11654_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout92 fanout93/X vssd1 vssd1 vccd1 vccd1 fanout92/X sky130_fd_sc_hd__buf_6
Xfanout81 _06937_/X vssd1 vssd1 vccd1 vccd1 fanout81/X sky130_fd_sc_hd__clkbuf_8
Xfanout70 _12706_/A vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__buf_6
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10605_ _11184_/A _10605_/B vssd1 vssd1 vccd1 vccd1 _10607_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ _11585_/A _11585_/B _11585_/C vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__and3_1
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12149__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10536_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13255_ _13260_/CLK hold102/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__dfxtp_1
X_10467_ hold197/A _10208_/B _10583_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _10467_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12253_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12208_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13188_/CLK hold227/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07576__A1 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10398_ _10398_/A _10398_/B _10398_/C vssd1 vssd1 vccd1 vccd1 _10399_/B sky130_fd_sc_hd__and3_1
X_12137_ _06890_/X _12125_/X _12136_/X vssd1 vssd1 vccd1 vccd1 _12137_/Y sky130_fd_sc_hd__o21ai_1
X_12068_ _12190_/B _12129_/B hold235/A vssd1 vssd1 vccd1 vccd1 _12068_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08525__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _11230_/D _11017_/X _11018_/Y vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06560_ _06560_/A _06560_/B vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12386__A _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08755_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08309_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _08160_/A _08160_/B _08160_/C vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07112_ _11955_/A _07112_/B vssd1 vssd1 vccd1 vccd1 _07112_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08092_ _08093_/A _08093_/B vssd1 vssd1 vccd1 vccd1 _08092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11060__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11060__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07043_ _07064_/B _07044_/B vssd1 vssd1 vccd1 vccd1 _07043_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11363__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08994_ _08996_/A _08996_/B _08251_/Y vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07319__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _07941_/Y _07985_/B _07940_/Y vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12312__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07319__B2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__nand2_1
X_09615_ _09771_/B _09463_/B _09457_/Y vssd1 vssd1 vccd1 vccd1 _09616_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__07154__S _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__B _11184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10323__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06542__A2 _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06827_ _06700_/B _06762_/X _06763_/X _12499_/A vssd1 vssd1 vccd1 vccd1 _08823_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06758_ _06753_/B _06752_/Y _06753_/Y _12501_/A vssd1 vssd1 vccd1 vccd1 _06761_/A
+ sky130_fd_sc_hd__a211o_1
X_09546_ _10126_/A _09546_/B _09546_/C vssd1 vssd1 vccd1 vccd1 _09547_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09475_/X _09476_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08295__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06689_ _06763_/B _06613_/A _12559_/B _06688_/X vssd1 vssd1 vccd1 vccd1 _07304_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08428_ fanout83/X _08782_/B2 _08813_/B1 _08565_/B vssd1 vssd1 vccd1 vccd1 _08429_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11370_ _11370_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11371_/B sky130_fd_sc_hd__or2_1
X_10321_ _10321_/A _10321_/B _10321_/C _10321_/D vssd1 vssd1 vccd1 vccd1 _10447_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13040_ _13040_/A _13040_/B vssd1 vssd1 vccd1 vccd1 _13040_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07007__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10183_ _10309_/B _10183_/B vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__xor2_4
Xfanout282 _06529_/X vssd1 vssd1 vccd1 vccd1 _12498_/C sky130_fd_sc_hd__buf_4
Xfanout271 hold177/X vssd1 vssd1 vccd1 vccd1 _13084_/B2 sky130_fd_sc_hd__buf_4
Xfanout260 _12080_/A vssd1 vssd1 vccd1 vccd1 _12495_/S sky130_fd_sc_hd__buf_4
Xfanout293 fanout298/X vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09180__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _13081_/B _13082_/A _12743_/X vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__a21o_1
X_12755_ hold5/X hold253/X vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__and2b_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ _09124_/S _10581_/X _11696_/B _09330_/A _11705_/X vssd1 vssd1 vccd1 vccd1
+ _11706_/X sky130_fd_sc_hd__o221a_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10719__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ _12686_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ _11876_/A _12141_/A fanout44/X fanout55/X vssd1 vssd1 vccd1 vccd1 _11638_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06932__A _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _11666_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__or2_1
XFILLER_0_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ _10519_/A _10519_/B vssd1 vssd1 vccd1 vccd1 _10520_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13238_ _13241_/CLK _13238_/D vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _13169_/CLK _13169_/D vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08210__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07763__A _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _07730_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07732_/B sky130_fd_sc_hd__xnor2_1
X_07661_ _07661_/A _07661_/B _07661_/C vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__nand3_1
X_06612_ instruction[0] instruction[1] _06850_/B instruction[31] pred_val vssd1 vssd1
+ vccd1 vccd1 _12527_/B sky130_fd_sc_hd__o311a_4
X_07592_ _07832_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__xnor2_1
X_09400_ _10009_/A fanout60/X _07070_/Y _09725_/B2 vssd1 vssd1 vccd1 vccd1 _09401_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06543_ reg1_val[31] _07604_/A vssd1 vssd1 vccd1 vccd1 _06545_/A sky130_fd_sc_hd__and2_1
X_09331_ _12115_/A _12297_/A _08276_/A _08823_/B vssd1 vssd1 vccd1 vccd1 _09331_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10608__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10608__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08277__A2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10084__A2 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _09263_/A _09263_/B vssd1 vssd1 vccd1 vccd1 _09262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11281__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13022__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12844__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__xnor2_1
X_09193_ _09193_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09268_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout226_A _08936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ reg1_val[3] _07026_/B vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__buf_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08977_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11195__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _08026_/A _08026_/B _08026_/C vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07859_ _07859_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _07961_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07712__B2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ fanout81/X fanout7/X fanout5/X _10957_/A vssd1 vssd1 vccd1 vccd1 _10871_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ _09396_/A _09396_/B _09395_/A vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12540_ _12539_/A _12536_/Y _12538_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11272__B2 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__A1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ _12478_/B _12471_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07228__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ _11509_/B _11422_/B vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__or2_1
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _06653_/B _11351_/X _11352_/Y _11350_/X vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _11656_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__xnor2_1
X_10304_ _10305_/A _10305_/B _10305_/C vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__o21ai_2
X_13023_ _13111_/A hold260/X vssd1 vssd1 vccd1 vccd1 _13235_/D sky130_fd_sc_hd__and2_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10235_ _10236_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__and2b_1
X_10166_ _10032_/A _10031_/B _10029_/Y vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__a21o_1
X_10097_ _10014_/A _10014_/B _10005_/Y vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07703__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__A1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _13034_/B _13035_/A _12759_/X vssd1 vssd1 vccd1 vccd1 _13040_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06927__A _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06646__B _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ _10999_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _11000_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12738_ hold95/X hold265/X vssd1 vssd1 vccd1 vccd1 _12738_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ hold35/X _12692_/B _12668_/Y _12970_/A vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__o211a_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12664__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__A1 _10796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08900_ _07588_/Y _07595_/B _07593_/Y vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__a21o_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _10117_/A fanout8/X fanout6/X _09880_/B2 vssd1 vssd1 vccd1 vccd1 _09881_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08777_/Y _09007_/B _08779_/A vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__o21ai_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11727__B fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08762_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10829__B2 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _09563_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07830_/B sky130_fd_sc_hd__xnor2_2
X_08693_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08712_/B sky130_fd_sc_hd__xor2_1
X_07644_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__and2_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout176_A _07011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12558__B _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _11124_/A _07574_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12248_/B sky130_fd_sc_hd__o21a_2
XANTENNA__11462__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ instruction[0] _06850_/B instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06526_/X sky130_fd_sc_hd__and4bb_1
X_09314_ _09312_/X _09313_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _09356_/B _09244_/B _09244_/C vssd1 vssd1 vccd1 vccd1 _09246_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08670__A2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _08973_/A _08973_/B _08974_/Y vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__11557__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08127_ _08741_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _08128_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07630__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _08741_/A _08058_/B vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09883__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _08688_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07015_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09094__S _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout89_A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _11794_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__xnor2_1
X_11971_ _11973_/A _11973_/B _11973_/C vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10922_ reg1_val[12] curr_PC[12] _10813_/X vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10847__C_N _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _10853_/A _10853_/B vssd1 vssd1 vccd1 vccd1 _10855_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10784_ _10785_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__and2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12523_ _12521_/Y _12523_/B vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__or3_1
XANTENNA__08949__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11548__A2 _11164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _12546_/B _12386_/B vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _11504_/A _11405_/B vssd1 vssd1 vccd1 vccd1 _11407_/B sky130_fd_sc_hd__and2_1
XFILLER_0_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _11838_/A _09039_/B _09039_/C _12179_/A vssd1 vssd1 vccd1 vccd1 _11336_/X
+ sky130_fd_sc_hd__a31o_1
X_13006_ hold279/A _13005_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__mux2_1
X_11267_ _11454_/B _11266_/Y _11636_/S vssd1 vssd1 vccd1 vccd1 _11267_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10508__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ _10203_/S _10217_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10218_/Y sky130_fd_sc_hd__o21ai_2
X_11198_ _12086_/A _11198_/B vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__xnor2_1
X_10149_ fanout82/X fanout63/X fanout60/X _06940_/A vssd1 vssd1 vccd1 vccd1 _10150_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08856__B _08858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07688__B1 _06984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09429__A1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09429__B2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07360_ _07361_/B _07361_/C _07361_/A vssd1 vssd1 vccd1 vccd1 _07364_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07291_ _07291_/A _07291_/B vssd1 vssd1 vccd1 vccd1 _07291_/Y sky130_fd_sc_hd__nand2_2
X_09030_ _09030_/A _09030_/B vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12197__C1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ _09299_/X _09306_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout293_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__A1 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _09862_/B _09863_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__nand2b_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08112__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ _10203_/S _09794_/B vssd1 vssd1 vccd1 vccd1 _09794_/X sky130_fd_sc_hd__or2_1
X_08814_ _08814_/A _08814_/B vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07915__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07951__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ _08749_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__and2b_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11475__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _08681_/B _08681_/A vssd1 vssd1 vccd1 vccd1 _08676_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10278__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07627_/A _07627_/B vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07558_ _07559_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07560_/A sky130_fd_sc_hd__and2_1
XANTENNA__08891__A2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06509_ _12664_/A vssd1 vssd1 vccd1 vccd1 _06509_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _07489_/A _07489_/B _07668_/A vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__or3_1
XANTENNA__09840__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09228_ _09563_/A _09228_/B _09228_/C vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__and3_1
XFILLER_0_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12727__A1 _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _10809_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09159_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ _12112_/A _12169_/X _12258_/C vssd1 vssd1 vccd1 vccd1 _12170_/Y sky130_fd_sc_hd__o21ai_1
X_11121_ _11231_/C _11119_/X _11120_/Y vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ curr_PC[13] _11051_/C curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11052_/Y sky130_fd_sc_hd__a21oi_1
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07382__A2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _12089_/A _11954_/B vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11466__B2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ _11885_/A _11885_/B vssd1 vssd1 vccd1 vccd1 _11889_/A sky130_fd_sc_hd__xnor2_1
X_10905_ _10905_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08882__A2 _08985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10836_ _12089_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08692__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _10767_/A _10767_/B _10767_/C vssd1 vssd1 vccd1 vccd1 _10768_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10698_ _09628_/X _09632_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ reg1_val[2] _12507_/B vssd1 vssd1 vccd1 vccd1 _12506_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ _12496_/A _12437_/B vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__or2_1
XANTENNA__11926__C1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ _12368_/A _12368_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12369_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06948__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06940__A _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__and2_1
XANTENNA__11558__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11319_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11320_/B sky130_fd_sc_hd__nor3_1
X_06860_ instruction[11] _06862_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
XFILLER_0_38_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08570__B2 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ _06790_/A _06790_/B _06837_/D vssd1 vssd1 vccd1 vccd1 _06792_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11457__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _08642_/B _08737_/A2 _08813_/B1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 _08531_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08461_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__or2_1
X_07412_ _07540_/B vssd1 vssd1 vccd1 vccd1 _07412_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09698__A _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08388_/X _08392_/B vssd1 vssd1 vccd1 vccd1 _08458_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07343_ _07343_/A _07343_/B vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10637__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07833__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ _07635_/S _07274_/B vssd1 vssd1 vccd1 vccd1 _07275_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12709__A1 _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09013_ _09013_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__or2_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12852__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08389__B2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12571__B _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08928__A3 _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11468__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09777_/A _09777_/B _10049_/A vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__a21oi_2
X_09846_ _11387_/A fanout36/X fanout34/X fanout71/X vssd1 vssd1 vccd1 vccd1 _09847_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _10252_/A _06989_/B vssd1 vssd1 vccd1 vccd1 _07023_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12299__A _12299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__xor2_4
X_08728_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08801_/A _08659_/B vssd1 vssd1 vccd1 vccd1 _08662_/A sky130_fd_sc_hd__xnor2_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10120__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10120__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__A1 _07152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ _11671_/A _11671_/B vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09401__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _10552_/A _10552_/B vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ instruction[4] vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
XFILLER_0_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08017__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ _12221_/A _12221_/B _12221_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12222_/X
+ sky130_fd_sc_hd__o211a_1
X_10483_ _10484_/A _10484_/B _10621_/A vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13069__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _12211_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09329__B1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ _12095_/B _12084_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__xnor2_1
X_11104_ _11104_/A _11104_/B vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__xnor2_1
X_11035_ _11135_/S _09291_/X _11034_/X vssd1 vssd1 vccd1 vccd1 _11035_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__07355__A2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ hold294/A _12985_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11439__A1 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11937_ _09293_/A _10204_/Y _10218_/Y _12073_/B2 _11936_/X vssd1 vssd1 vccd1 vccd1
+ _11937_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11868_ _06847_/X _11864_/X _11867_/X vssd1 vssd1 vccd1 vccd1 dest_val[23] sky130_fd_sc_hd__o21ai_4
X_10819_ hold207/A _11781_/B _10927_/B _10818_/Y _11448_/A vssd1 vssd1 vccd1 vccd1
+ _10826_/A sky130_fd_sc_hd__a311o_1
X_11799_ _11799_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11801_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11375__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13116__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _07961_/A _07961_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08791__A1 _08784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09981__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06912_ reg1_val[10] reg1_val[11] reg1_val[12] _06993_/B vssd1 vssd1 vccd1 vccd1
+ _07091_/B sky130_fd_sc_hd__or4_4
XANTENNA__11127__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _09880_/B2 fanout8/X fanout6/X _09885_/A vssd1 vssd1 vccd1 vccd1 _09701_/B
+ sky130_fd_sc_hd__o22a_2
X_07892_ _07892_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07972_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10920__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _09310_/X _09312_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__mux2_1
X_06843_ _09151_/A vssd1 vssd1 vccd1 vccd1 _06843_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06774_ _10328_/B _10328_/C _10331_/A vssd1 vssd1 vccd1 vccd1 _06775_/B sky130_fd_sc_hd__o21ai_1
X_09562_ _09563_/A _09563_/B vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08513_ _08513_/A _08513_/B vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__xor2_1
X_09493_ _09493_/A _09493_/B vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08444_ _08607_/A _08444_/B vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _08417_/A _08417_/B vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07326_ _07327_/B _07327_/C _07327_/A vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ _09420_/A _07257_/B vssd1 vssd1 vccd1 vccd1 _07259_/B sky130_fd_sc_hd__xnor2_4
X_07188_ _12668_/A _12141_/A _09237_/A _07391_/B vssd1 vssd1 vccd1 vccd1 _07189_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08231__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11198__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__and2_1
XANTENNA__08534__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ _13071_/A hold248/X vssd1 vssd1 vccd1 vccd1 _13161_/D sky130_fd_sc_hd__and2_1
XANTENNA__06739__B _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12771_ hold25/X hold279/A vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11722_ _11723_/A _11723_/B _11723_/C vssd1 vssd1 vccd1 vccd1 _11724_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10277__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout60 _12094_/A vssd1 vssd1 vccd1 vccd1 fanout60/X sky130_fd_sc_hd__buf_6
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout71 _12706_/A vssd1 vssd1 vccd1 vccd1 fanout71/X sky130_fd_sc_hd__buf_4
X_10604_ fanout78/X _12148_/A _12201_/A _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10605_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout82 fanout83/X vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_6
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 _07278_/Y vssd1 vssd1 vccd1 vccd1 fanout93/X sky130_fd_sc_hd__buf_8
XFILLER_0_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11584_ _11585_/A _11585_/B _11585_/C vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _10535_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10537_/C sky130_fd_sc_hd__xor2_1
X_13254_ _13254_/CLK _13254_/D vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
X_10466_ _10208_/B _10583_/B hold197/A vssd1 vssd1 vccd1 vccd1 _10466_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12149__A2 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _13185_/CLK _13185_/D vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__dfxtp_1
X_12205_ _12205_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12206_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _12130_/Y _12131_/X _12135_/X _12128_/X vssd1 vssd1 vccd1 vccd1 _12136_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09970__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10397_ _10398_/B _10398_/C _10398_/A vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ hold228/A _12067_/B vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__or2_1
XANTENNA__10740__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _11230_/D _11017_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _11018_/Y sky130_fd_sc_hd__o21ai_1
X_12969_ hold243/X _12663_/B _12968_/X _12664_/A vssd1 vssd1 vccd1 vccd1 hold244/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08289__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _08160_/A _08160_/B _08160_/C vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__and3_1
XFILLER_0_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _11072_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08093_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11060__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07042_ _07064_/A _07065_/A _07065_/B _07065_/C _07058_/B1 vssd1 vssd1 vccd1 vccd1
+ _07044_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07016__A1 _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08993_ _09043_/A _08998_/A _09043_/B _08849_/X vssd1 vssd1 vccd1 vccd1 _08996_/B
+ sky130_fd_sc_hd__a31o_1
X_07944_ _10853_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07319__A2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _07875_/A _07875_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__or2_4
X_09614_ _09614_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09616_/A sky130_fd_sc_hd__nor2_2
XANTENNA__10323__A1 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__C fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ reg1_val[1] _09479_/S vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12076__A1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09545_ _09546_/B _09546_/C _10126_/A vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__a21o_1
X_09476_ _09075_/X _09093_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06688_ reg2_val[11] _06748_/B vssd1 vssd1 vccd1 vccd1 _06688_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08427_ _08427_/A _08427_/B _08427_/C _08427_/D vssd1 vssd1 vccd1 vccd1 _08427_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08358_ _08358_/A _08427_/A vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ _07294_/A _07294_/B _07381_/A vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__a21oi_1
X_08289_ _08740_/A2 _12688_/A _12690_/A _09725_/B2 vssd1 vssd1 vccd1 vccd1 _08290_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10320_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10321_/D sky130_fd_sc_hd__or2_1
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _10251_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06766__B1 _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _10051_/A _10309_/A _10051_/B _10047_/Y vssd1 vssd1 vccd1 vccd1 _10183_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout250 _09146_/X vssd1 vssd1 vccd1 vccd1 _12179_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11656__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _13110_/A2 vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__buf_4
Xfanout261 _06848_/Y vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__clkbuf_16
Xfanout283 _06700_/B vssd1 vssd1 vccd1 vccd1 _06748_/B sky130_fd_sc_hd__clkbuf_4
Xfanout294 fanout298/X vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__buf_4
XANTENNA__09180__A1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__B2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__C_N _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _13077_/A _12822_/B _12745_/X vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ hold298/A hold3/X vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ _09138_/X _11704_/X _06619_/B vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__a21o_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ hold27/X _12686_/B _12684_/Y _13013_/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__o211a_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11027__C1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08691__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09796__A _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ _11632_/X _11635_/Y _11636_/S vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__mux2_8
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11566_/B _11567_/B vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08443__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13111__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _10519_/A _10519_/B vssd1 vssd1 vccd1 vccd1 _10518_/Y sky130_fd_sc_hd__nand2_1
X_13237_ _13241_/CLK _13237_/D vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11498_ _11499_/B _11499_/A vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10449_ _10449_/A _10681_/A _10449_/C vssd1 vssd1 vccd1 vccd1 _10450_/C sky130_fd_sc_hd__nand3_1
X_13168_ _13169_/CLK hold199/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13099_ _12735_/X _13099_/B vssd1 vssd1 vccd1 vccd1 _13100_/B sky130_fd_sc_hd__nand2b_1
X_12119_ _12112_/A _09053_/Y _09055_/Y _09145_/Y _12118_/Y vssd1 vssd1 vccd1 vccd1
+ _12119_/X sky130_fd_sc_hd__o311a_1
XANTENNA__07763__B _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _07660_/A _07662_/A _07660_/C vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__and3_1
X_06611_ _11782_/S _06611_/B vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__nor2_1
X_07591_ fanout77/X _10481_/A _07000_/A fanout74/X vssd1 vssd1 vccd1 vccd1 _07592_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06542_ _06753_/B _06665_/A2 _06540_/B _06528_/X vssd1 vssd1 vccd1 vccd1 _07184_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09330_ _09330_/A _09330_/B vssd1 vssd1 vccd1 vccd1 _09330_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10608__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _08942_/A _08942_/B _08940_/Y vssd1 vssd1 vccd1 vccd1 _09263_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__B2 _07137_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11281__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _09193_/B _09193_/A vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11569__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout121_A _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _08143_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ _08074_/A _08074_/B vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ reg1_val[0] reg1_val[1] reg1_val[2] _07128_/A vssd1 vssd1 vccd1 vccd1 _07026_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08115__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11476__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _08977_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08976_/X sky130_fd_sc_hd__and2_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__A1 _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _07927_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _08026_/C sky130_fd_sc_hd__xnor2_1
X_07858_ _07858_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07961_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06809_ _12117_/A _06808_/X _06803_/Y vssd1 vssd1 vccd1 vccd1 _06809_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07712__A2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _09568_/A _11564_/A fanout38/X _09698_/A vssd1 vssd1 vccd1 vccd1 _07790_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09528_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__or2_2
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout34_A _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09459_ _08981_/A _08981_/B _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09459_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11272__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _12457_/Y _12478_/C _12480_/B vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07228__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__A1 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _11547_/A _11421_/B _11421_/C vssd1 vssd1 vccd1 vccd1 _11422_/B sky130_fd_sc_hd__and3_1
X_11352_ _06978_/A _12280_/A _09147_/X _06653_/A _06847_/X vssd1 vssd1 vccd1 vccd1
+ _11352_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10305_/C sky130_fd_sc_hd__xor2_1
X_11283_ _12095_/A fanout50/X _07988_/B fanout60/X vssd1 vssd1 vccd1 vccd1 _11284_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ hold259/X _06858_/B _13021_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold260/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07864__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _10108_/A _10108_/B _10105_/A vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10096_ _10041_/A _10041_/B _10042_/X vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__09832__A1_N _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12806_ _13029_/B _13030_/A _12761_/X vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06927__B _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10998_ _10997_/A _10997_/B _10999_/A vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10449__B _10681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12737_ hold49/X hold275/X vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ _12668_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _12668_/Y sky130_fd_sc_hd__nand2_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ hold168/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11701_/B sky130_fd_sc_hd__or2_1
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _12599_/A _12599_/B _12599_/C vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__or3_2
XANTENNA__10223__B1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07774__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08830_ _09008_/A _09008_/B _08794_/X vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__o21ba_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09144__A1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__A1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08762_/B _08762_/A vssd1 vssd1 vccd1 vccd1 _08761_/X sky130_fd_sc_hd__and2b_1
X_07712_ _06828_/A _12716_/A _08765_/A _12714_/A vssd1 vssd1 vccd1 vccd1 _07713_/B
+ sky130_fd_sc_hd__o22a_1
X_08692_ _08734_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _08712_/A sky130_fd_sc_hd__xnor2_1
X_07643_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__or2_1
XFILLER_0_88_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09313_ _09105_/X _09107_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07574_ reg1_val[30] _07574_/B vssd1 vssd1 vccd1 vccd1 _07574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06525_ instruction[0] pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06863_/A
+ sky130_fd_sc_hd__and3b_1
XANTENNA__07014__A _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07949__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ _09356_/B _09244_/B _09244_/C vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__or3_2
X_09175_ _08978_/A _08978_/B _08976_/X vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08126_ _10876_/A1 _08740_/A2 _08755_/B _10957_/A vssd1 vssd1 vccd1 vccd1 _08127_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07630__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07630__B2 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _08755_/B fanout93/X _10647_/A _08740_/A2 vssd1 vssd1 vccd1 vccd1 _08058_/B
+ sky130_fd_sc_hd__o22a_1
X_07008_ reg1_val[6] _07008_/B vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06736__A3 _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__xnor2_1
X_11970_ _11970_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11973_/C sky130_fd_sc_hd__xnor2_1
X_10921_ _10921_/A _10921_/B vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10852_ fanout78/X fanout9/X fanout3/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10853_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ reg1_val[5] _12522_/B vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ _12453_/A _12453_/B vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08949__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12384_ reg1_val[10] curr_PC[10] _12495_/S vssd1 vssd1 vccd1 vccd1 _12386_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08949__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _11404_/A _11404_/B _11404_/C vssd1 vssd1 vccd1 vccd1 _11405_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11953__B1 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11335_ _11838_/A _09039_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _11335_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ curr_PC[16] _11265_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11266_/Y sky130_fd_sc_hd__a21oi_1
X_13005_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13005_/Y sky130_fd_sc_hd__xnor2_1
X_10217_ _11033_/A _09127_/X _09166_/B vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10508__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10508__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11197_ _11663_/A fanout14/X fanout52/X _11739_/A vssd1 vssd1 vccd1 vccd1 _11198_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09374__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _09972_/A _09972_/B _09969_/A vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__a21o_1
X_10079_ hold213/A _10208_/B _10207_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _10079_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07688__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__A _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__A1 _07157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__B2 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B1 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09429__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ _06931_/B _07295_/A _07295_/B _06930_/X vssd1 vssd1 vccd1 vccd1 _07290_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09062__B1 _09464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _09931_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11172__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ _09863_/B _09862_/B vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__nand2b_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07009__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09793_ _09792_/X _09655_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__mux2_1
X_08813_ _08813_/A1 _09237_/A _08813_/B1 _06828_/A vssd1 vssd1 vccd1 vccd1 _08814_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07915__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08744_ _08744_/A _08753_/A vssd1 vssd1 vccd1 vccd1 _08749_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06848__A _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06567__B _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _08682_/A _08708_/A _08708_/B _08668_/Y vssd1 vssd1 vccd1 vccd1 _08681_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07627_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07557_ _07916_/A _07557_/B vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__xnor2_1
X_06508_ _13219_/Q vssd1 vssd1 vccd1 vccd1 _06508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07679__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07488_ _07489_/B _07668_/A _07489_/A vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09840__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ _09862_/B _09227_/B _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/C sky130_fd_sc_hd__nand3_1
XANTENNA__12727__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ _11135_/S _09158_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ reg1_val[10] reg1_val[21] _09092_/S vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08109_ _08109_/A _08110_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__nor2_2
X_11120_ _11231_/C _11119_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__o21ai_1
X_11051_ curr_PC[13] curr_PC[14] _11051_/C vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__and3_1
X_10002_ _10850_/A _10002_/B vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _12148_/A fanout11/X _07391_/B _12201_/A vssd1 vssd1 vccd1 vccd1 _11954_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11466__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06878__C1 _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11884_ _12095_/A fanout8/X fanout6/X _11950_/A vssd1 vssd1 vccd1 vccd1 _11885_/B
+ sky130_fd_sc_hd__o22a_1
X_10904_ _10904_/A _10904_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10905_/B sky130_fd_sc_hd__nor3_1
X_10835_ _11169_/A fanout11/X fanout44/X _11297_/A vssd1 vssd1 vccd1 vccd1 _10836_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10767_/A _10767_/B _10767_/C vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12504_/A _12503_/B _12501_/Y vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__a21oi_4
X_10697_ _10574_/Y _10578_/B _10694_/Y _10695_/X vssd1 vssd1 vccd1 vccd1 _10697_/Y
+ sky130_fd_sc_hd__a211oi_2
X_12436_ _12496_/A _12437_/B vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12367_ _12368_/A _12368_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12375_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12298_ _12267_/A _12223_/B _12223_/C _12223_/A vssd1 vssd1 vccd1 vccd1 _12299_/B
+ sky130_fd_sc_hd__o31a_1
X_11318_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__o21a_1
X_11249_ hold218/A _11249_/B vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__or2_1
XANTENNA__11154__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__A2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06790_ _06790_/A _06790_/B vssd1 vssd1 vccd1 vccd1 _06790_/X sky130_fd_sc_hd__and2_1
XFILLER_0_54_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11457__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09979__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07540_/B sky130_fd_sc_hd__and2_1
X_08391_ _08388_/B _08388_/C _08388_/A vssd1 vssd1 vccd1 vccd1 _08392_/B sky130_fd_sc_hd__a21o_1
X_07342_ _07343_/A _07343_/B vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09698__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__A2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07833__B2 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _12142_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12709__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__and2_1
XFILLER_0_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08389__A2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06850__B _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold148/X vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__B1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__buf_2
XFILLER_0_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__buf_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__A1_N _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11145__A1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09914_ _10310_/A _10311_/A vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10091__C _10091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__xor2_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _06977_/A fanout77/X _06985_/A _12710_/A vssd1 vssd1 vccd1 vccd1 _06989_/B
+ sky130_fd_sc_hd__o22a_1
X_09776_ _08982_/A _09775_/Y _09773_/Y vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__a21bo_2
X_08727_ _08727_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _09004_/A sky130_fd_sc_hd__nor2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__A1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ _08782_/A2 _08733_/B1 _08735_/A2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08659_/B
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13208_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10120__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08589_ _08589_/A _08589_/B vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10620_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10620_/X sky130_fd_sc_hd__and2_1
XFILLER_0_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10552_/A _10552_/B vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11081__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10482_ _10607_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10621_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12221_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10592__C1 _10591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _12205_/A _12152_/B vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__nand2_1
X_12083_ _12201_/A fanout8/X fanout6/X _12148_/A vssd1 vssd1 vccd1 vccd1 _12084_/B
+ sky130_fd_sc_hd__o22a_1
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__nor2_1
X_11034_ _11134_/S _10073_/X _11033_/Y _10809_/A vssd1 vssd1 vccd1 vccd1 _11034_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07760__B1 _06999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _12985_/A _12985_/B vssd1 vssd1 vccd1 vccd1 _12985_/Y sky130_fd_sc_hd__xnor2_1
X_11936_ _07029_/B _06905_/Y _11625_/B _06579_/A _11935_/Y vssd1 vssd1 vccd1 vccd1
+ _11936_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ _12080_/A _11867_/B _11941_/B vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__or3_1
X_10818_ _11781_/B _10927_/B hold207/A vssd1 vssd1 vccd1 vccd1 _10818_/Y sky130_fd_sc_hd__a21oi_1
X_11798_ fanout13/X fanout9/A fanout4/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11799_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07112__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _10749_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12672__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12419_ reg1_val[15] curr_PC[15] _12444_/S vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__B2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13116__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _07960_/A _07960_/B vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06911_ reg1_val[7] reg1_val[8] reg1_val[9] _06970_/B vssd1 vssd1 vccd1 vccd1 _06993_/B
+ sky130_fd_sc_hd__or4_2
X_07891_ _07889_/A _07889_/B _07890_/Y vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__o21ai_2
X_09630_ _09309_/X _09319_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__mux2_1
X_06842_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__nand2_4
X_06773_ _06772_/A _06772_/B _06830_/D vssd1 vssd1 vccd1 vccd1 _10328_/C sky130_fd_sc_hd__a21boi_1
X_09561_ _09862_/B _09561_/B vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__xnor2_1
X_08512_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08841_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _09490_/Y _09492_/B vssd1 vssd1 vccd1 vccd1 _09493_/B sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout151_A _06984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _08606_/A2 _08737_/A2 _08733_/B1 _08642_/B vssd1 vssd1 vccd1 vccd1 _08444_/B
+ sky130_fd_sc_hd__o22a_1
X_08374_ _08374_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _08417_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09256__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07325_ _07337_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07327_/C sky130_fd_sc_hd__and2_1
XFILLER_0_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07256_ _08765_/A _12201_/A fanout9/A _06828_/A vssd1 vssd1 vccd1 vccd1 _07257_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07187_ _12085_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07187_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08231__B2 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__A1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08782__A2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _11794_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09830_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08534__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09760_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10629__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ hold255/X hold11/X vssd1 vssd1 vccd1 vccd1 _13009_/B sky130_fd_sc_hd__nand2b_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11805_/A _11721_/B vssd1 vssd1 vccd1 vccd1 _11723_/C sky130_fd_sc_hd__nand2_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11652_ _11956_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout61 _07043_/Y vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__clkbuf_8
Xfanout72 _07002_/Y vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__clkbuf_8
Xfanout50 fanout51/X vssd1 vssd1 vccd1 vccd1 fanout50/X sky130_fd_sc_hd__buf_6
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _10504_/A _10504_/B _10506_/X vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__o21ai_2
Xfanout83 _06923_/Y vssd1 vssd1 vccd1 vccd1 fanout83/X sky130_fd_sc_hd__buf_6
XANTENNA__11054__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _11668_/B _11583_/B vssd1 vssd1 vccd1 vccd1 _11585_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout94 _08333_/B vssd1 vssd1 vccd1 vccd1 _07239_/A sky130_fd_sc_hd__buf_6
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ _11184_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10535_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12003__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13253_ _13253_/CLK _13253_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
X_10465_ hold200/A hold241/A _10465_/C vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__or3_1
X_13184_ _13185_/CLK hold230/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12204_ _12205_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10396_ _10395_/B _10395_/C _10529_/A vssd1 vssd1 vccd1 vccd1 _10398_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ _09293_/A _09796_/B _09815_/X _09330_/A _12134_/Y vssd1 vssd1 vccd1 vccd1
+ _12135_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09970__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09970__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08525__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11230_/C _10909_/B _11232_/A vssd1 vssd1 vccd1 vccd1 _11017_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ hold249/A _12967_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08289__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ hold90/X _12663_/B _12686_/B _12499_/A vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__a22o_1
X_11919_ _11918_/A _11918_/B _09498_/A vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07110_ _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _07110_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _08737_/A2 _08333_/B _08813_/B1 fanout43/X vssd1 vssd1 vccd1 vccd1 _08091_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07041_ _07041_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07041_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__11299__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08992_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _11983_/B sky130_fd_sc_hd__and2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ fanout79/X _08715_/A2 _08689_/B1 _08430_/B vssd1 vssd1 vccd1 vccd1 _07944_/B
+ sky130_fd_sc_hd__o22a_1
X_07874_ _09428_/A fanout41/X _08135_/B _09568_/A vssd1 vssd1 vccd1 vccd1 _07875_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11520__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06825_ instruction[6] _06824_/X _06813_/X vssd1 vssd1 vccd1 vccd1 _06825_/X sky130_fd_sc_hd__a21bo_1
X_09613_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__and3_1
XANTENNA__12858__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06856__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06756_ _06753_/B _06752_/Y _06753_/Y vssd1 vssd1 vccd1 vccd1 _06756_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _07075_/A _07075_/B _09725_/B2 vssd1 vssd1 vccd1 vccd1 _09546_/C sky130_fd_sc_hd__a21o_1
X_09475_ _09071_/X _09078_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09475_/X sky130_fd_sc_hd__mux2_1
X_06687_ _10823_/A _06687_/B vssd1 vssd1 vccd1 vccd1 _06831_/D sky130_fd_sc_hd__nand2_1
XANTENNA__10378__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _08358_/A _08357_/C _08357_/B vssd1 vssd1 vccd1 vccd1 _08427_/D sky130_fd_sc_hd__a21o_1
XANTENNA__09229__B1 _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _08358_/A _08357_/B _08357_/C vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07308_ _07380_/A _07380_/B vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__and2_1
X_08288_ _08714_/A _08288_/B vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07687__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ _07239_/A vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__inv_2
X_10250_ _10607_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06766__B2 _06511_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10181_/A _10181_/B vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__xor2_4
Xfanout240 _06736_/X vssd1 vssd1 vccd1 vccd1 _07108_/C sky130_fd_sc_hd__buf_4
Xfanout273 hold177/X vssd1 vssd1 vccd1 vccd1 _13110_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout251 _09139_/Y vssd1 vssd1 vccd1 vccd1 _12265_/C1 sky130_fd_sc_hd__buf_4
Xfanout262 _06847_/X vssd1 vssd1 vccd1 vccd1 _11636_/S sky130_fd_sc_hd__clkbuf_16
Xfanout295 fanout298/X vssd1 vssd1 vccd1 vccd1 _12955_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout284 _06754_/B vssd1 vssd1 vccd1 vccd1 _06700_/B sky130_fd_sc_hd__buf_6
XANTENNA__07715__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A2 _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__B2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__A1 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ _12745_/X _12822_/B vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__nand2b_1
X_12753_ hold287/A hold1/X vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__nand2b_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11704_ _09501_/B _11625_/B _11704_/S vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__mux2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12684_ _12684_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12684_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08691__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08691__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _11712_/B _11635_/B vssd1 vssd1 vccd1 vccd1 _11635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _11567_/B _11566_/B vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08443__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08443__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10519_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _13251_/CLK _13236_/D vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ _10449_/A _10449_/C _10681_/A vssd1 vssd1 vccd1 vccd1 _10450_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _13169_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07954__B1 _07953_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ fanout7/X _10647_/A fanout5/X _10506_/A vssd1 vssd1 vccd1 vccd1 _10380_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13098_ _13103_/A _13098_/B vssd1 vssd1 vccd1 vccd1 _13251_/D sky130_fd_sc_hd__and2_1
X_12118_ _12112_/A _09053_/Y _09055_/Y vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__o21ai_1
X_12049_ _09465_/A _09056_/C _09056_/B vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07706__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07182__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ reg1_val[22] _07028_/B vssd1 vssd1 vccd1 vccd1 _06611_/B sky130_fd_sc_hd__nor2_1
X_07590_ _10126_/A _07590_/B vssd1 vssd1 vccd1 vccd1 _07594_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06541_ _06665_/A2 _06657_/B1 _06528_/X vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09260_ _09394_/B _09260_/B vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__nand2_2
XANTENNA__13007__B2 hold177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _10853_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11018__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _09191_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11569__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11569__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ _08143_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ _08074_/A _08074_/B vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__or2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ _07415_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _08975_/A _08975_/B vssd1 vssd1 vccd1 vccd1 _08977_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09227__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__buf_1
X_07926_ _08012_/A _08012_/B vssd1 vssd1 vccd1 vccd1 _08026_/B sky130_fd_sc_hd__and2b_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _07857_/A _07857_/B vssd1 vssd1 vccd1 vccd1 _07858_/B sky130_fd_sc_hd__and2_1
X_06808_ _12056_/A _06807_/X _12115_/B vssd1 vssd1 vccd1 vccd1 _06808_/X sky130_fd_sc_hd__o21a_1
X_07788_ _09979_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__xnor2_1
X_06739_ reg1_val[4] _07108_/C vssd1 vssd1 vccd1 vccd1 _06739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09527_ _09526_/B _09527_/B vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08122__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _09458_/A _09458_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08409_ _08411_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08412_/A sky130_fd_sc_hd__and2_1
X_09389_ _09389_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__or2_1
XANTENNA__10836__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__A2 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _11421_/B _11421_/C _11547_/A vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__a21oi_1
X_11351_ _06653_/A _09501_/B _09138_/X vssd1 vssd1 vccd1 vccd1 _11351_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07210__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__or2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _12086_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__xnor2_1
X_13021_ hold261/A _13020_/Y hold246/X vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__mux2_1
X_10233_ _10429_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__or2_1
XANTENNA__07936__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _10164_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__nor2_2
X_10095_ _10046_/A _10046_/B _10044_/X vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_107_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _13024_/B _13025_/A _12763_/X vssd1 vssd1 vccd1 vccd1 _13030_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10997_ _10997_/A _10997_/B vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__nor2_1
X_12736_ hold293/X hold81/X vssd1 vssd1 vccd1 vccd1 _13099_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07104__B _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12667_ _12248_/B _12926_/A2 hold34/X _13013_/A vssd1 vssd1 vccd1 vccd1 _13126_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10746__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ _10713_/Y _11617_/Y _12125_/S vssd1 vssd1 vccd1 vccd1 _11618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12598_ reg1_val[20] _12615_/B vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap215 _06889_/Y vssd1 vssd1 vccd1 vccd1 _09156_/B sky130_fd_sc_hd__buf_4
X_11549_ _11415_/Y _11506_/X _11547_/X _11421_/B _11508_/B vssd1 vssd1 vccd1 vccd1
+ _11600_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ _13222_/CLK hold140/X vssd1 vssd1 vccd1 vccd1 _13219_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10481__A _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13217_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _08759_/A _08776_/A vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__and2b_1
X_07711_ _09564_/A _07711_/B vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__xnor2_2
X_08691_ _08219_/B _08735_/A2 _08735_/B1 _08815_/B vssd1 vssd1 vccd1 vccd1 _08692_/B
+ sky130_fd_sc_hd__o22a_1
X_07642_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12201__A _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ _09101_/X _09104_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09312_/X sky130_fd_sc_hd__mux2_1
X_07573_ _08897_/B _07573_/B vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08104__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06524_ _06892_/A _06524_/B vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__nor2_8
XFILLER_0_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout231_A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09244_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _06520_/Y _09173_/X _11713_/A vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__mux2_8
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _08607_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07630__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08714_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__xnor2_1
X_07007_ reg1_val[4] reg1_val[5] _07050_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _07008_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11714__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _08959_/B _08959_/A vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12675__C1 _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _07909_/A _07909_/B _07909_/C vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__nand3_2
X_08889_ _11726_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10920_ _10920_/A curr_PC[13] vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11950__A _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _10948_/A _10851_/B vssd1 vssd1 vccd1 vccd1 _10855_/A sky130_fd_sc_hd__and2_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ reg1_val[5] _12522_/B vssd1 vssd1 vccd1 vccd1 _12521_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09420__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12452_ _12496_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12453_/B sky130_fd_sc_hd__or2_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _11404_/A _11404_/B _11404_/C vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__a21o_1
X_12383_ _12389_/B _12383_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XANTENNA__11953__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07875__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__B2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ _11331_/X _11332_/X _11333_/Y vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ curr_PC[16] curr_PC[17] _11265_/C vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__and3_1
X_13004_ _12771_/X _13004_/B vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__nand2b_1
X_10216_ _11448_/A _10208_/X _10209_/Y _10215_/X vssd1 vssd1 vccd1 vccd1 _10216_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11705__A1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10508__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11196_ _11196_/A _11196_/B vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__xor2_1
X_10147_ _10146_/B _10146_/C _10146_/A vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10078_ _10208_/B _10207_/B hold213/A vssd1 vssd1 vccd1 vccd1 _10078_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11469__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__B _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__A2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06954__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ hold19/X _12720_/B _12718_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__o211a_1
XANTENNA__09330__A _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11641__B1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06673__B _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12197__A1 _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09930_ _09928_/Y _09930_/B vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09861_ _10252_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__xnor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _09103_/X _09126_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__mux2_1
X_08812_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__xnor2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08744_/A _08743_/B _08743_/C vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__nand3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout279_A _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09224__B _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__nor2_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07625_/X sky130_fd_sc_hd__or2_1
X_07556_ fanout51/X _07137_/Y fanout49/X _12686_/A vssd1 vssd1 vccd1 vccd1 _07557_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09825__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__inv_2
XANTENNA__09240__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _09227_/B _09227_/C _09862_/B vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06654__A3 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ _09165_/B vssd1 vssd1 vccd1 vccd1 _09158_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ reg1_val[11] reg1_val[20] _09092_/S vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _08535_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08110_/B sky130_fd_sc_hd__xnor2_4
X_08039_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08042_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11148__C1 _11146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout94_A _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11050_ _11019_/X _11022_/X _11027_/X _11049_/X _11636_/S vssd1 vssd1 vccd1 vccd1
+ _11050_/X sky130_fd_sc_hd__a41o_1
X_10001_ _06940_/A fanout63/X fanout55/X fanout83/X vssd1 vssd1 vccd1 vccd1 _10002_/B
+ sky130_fd_sc_hd__o22a_2
X_11952_ _11948_/A _11877_/B _11880_/A vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10123__B1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11883_ _11883_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10903_ _10904_/A _10904_/B _10904_/C vssd1 vssd1 vccd1 vccd1 _10905_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10834_ _11636_/S _10831_/X _11051_/C _10833_/Y vssd1 vssd1 vccd1 vccd1 dest_val[12]
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _12504_/A _12504_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xnor2_4
X_10765_ _10873_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _10767_/C sky130_fd_sc_hd__or2_1
XANTENNA__06645__A3 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _10694_/Y _10695_/X _10574_/Y _10578_/B vssd1 vssd1 vccd1 vccd1 _10696_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ reg1_val[18] curr_PC[18] _12444_/S vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11926__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _12375_/A _12366_/B vssd1 vssd1 vccd1 vccd1 _12368_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09296__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11319_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _12297_/A _12297_/B vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12016__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09347__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _11696_/A _11246_/Y _11247_/X _06889_/Y vssd1 vssd1 vccd1 vccd1 _11248_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ _11180_/A _11180_/B _11180_/C vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06949__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12686__A _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07410_ _12668_/A _07391_/B _07391_/C _07391_/D vssd1 vssd1 vccd1 vccd1 _07411_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ _09564_/A _08390_/B vssd1 vssd1 vccd1 vccd1 _08458_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07343_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10417__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07272_ _12141_/A _09237_/A _07391_/B _09428_/A vssd1 vssd1 vccd1 vccd1 _07273_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07833__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09017_/A sky130_fd_sc_hd__and2_1
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07597__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__C1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _10311_/A vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__inv_2
XANTENNA__11145__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__D _10091_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__and2_1
XANTENNA__10353__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _06987_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _06987_/Y sky130_fd_sc_hd__xnor2_1
X_09775_ _11163_/A vssd1 vssd1 vccd1 vccd1 _09775_/Y sky130_fd_sc_hd__inv_2
X_08726_ _08726_/A _08726_/B _08726_/C vssd1 vssd1 vccd1 vccd1 _08727_/B sky130_fd_sc_hd__and3_1
XANTENNA__11853__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08657_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08669_/A sky130_fd_sc_hd__or2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _07608_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08588_ _08588_/A _08588_/B _08588_/C vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__or3_1
X_07539_ _07546_/A _07546_/B _07546_/C vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11605__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10550_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11081__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11081__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ _09209_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09210_/B sky130_fd_sc_hd__nand2_1
X_10481_ _10481_/A fanout3/X vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _06819_/X _12219_/X _12263_/S vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08785__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _12205_/A _12152_/B vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12082_ curr_PC[27] _12082_/B vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__xor2_1
X_11102_ _11102_/A _11102_/B _11102_/C vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__and3_1
X_11033_ _11033_/A _11033_/B vssd1 vssd1 vccd1 vccd1 _11033_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07760__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ _13111_/A hold295/X vssd1 vssd1 vccd1 vccd1 _13227_/D sky130_fd_sc_hd__and2_1
XANTENNA__07760__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11935_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11866_ curr_PC[22] curr_PC[23] _11866_/C vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__and3_1
X_10817_ _13170_/Q _10817_/B vssd1 vssd1 vccd1 vccd1 _10927_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11797_ _11879_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10748_ _10749_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10748_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12418_ _12424_/B _12418_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XFILLER_0_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10679_ _10794_/A _10562_/B _10793_/B vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11375__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ reg1_val[5] curr_PC[5] _12495_/S vssd1 vssd1 vccd1 vccd1 _12351_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ reg1_val[4] reg1_val[5] reg1_val[6] _07050_/B vssd1 vssd1 vccd1 vccd1 _06970_/B
+ sky130_fd_sc_hd__or4_2
X_07890_ _07900_/B _07900_/A vssd1 vssd1 vccd1 vccd1 _07890_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__06679__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ instruction[6] _06839_/X _06840_/Y vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06772_ _06772_/A _06772_/B vssd1 vssd1 vccd1 vccd1 _06772_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12088__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _09727_/A fanout9/X fanout4/X _07056_/Y vssd1 vssd1 vccd1 vccd1 _09561_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09491_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09492_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11835__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08511_ _08553_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__and2_1
XFILLER_0_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _08452_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08464_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11048__D1 _11039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout144_A _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _08310_/B _08373_/B vssd1 vssd1 vccd1 vccd1 _08374_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09256__B2 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09256__A1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _11955_/A _07324_/B vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12260__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07255_ _07255_/A _07255_/B vssd1 vssd1 vccd1 vccd1 _12728_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06861__B _06862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ _07186_/A _07186_/B vssd1 vssd1 vccd1 vccd1 _07186_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__12012__B1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B1 _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12315__A1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__B _08788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10326__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ fanout15/X _07763_/B _12690_/A fanout52/X vssd1 vssd1 vccd1 vccd1 _09828_/B
+ sky130_fd_sc_hd__o22a_1
X_09758_ _09757_/A _09757_/B _09759_/A vssd1 vssd1 vccd1 vccd1 _09758_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout57_A _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _08709_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08711_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10629__B2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11719_/B _11720_/B vssd1 vssd1 vccd1 vccd1 _11721_/B sky130_fd_sc_hd__nand2b_1
X_09689_ _09689_/A _09689_/B vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__xnor2_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 fanout41/X vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__buf_6
X_11651_ _07069_/X _07154_/X _07799_/B _07075_/Y vssd1 vssd1 vccd1 vccd1 _11652_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout62 _12720_/A vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__clkbuf_8
Xfanout73 _12710_/A vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__buf_6
Xfanout51 _07135_/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__buf_8
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__or2_1
X_10602_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10674_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11054__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout84 _11235_/A vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__buf_4
XFILLER_0_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout95 _07238_/Y vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__buf_8
X_10533_ fanout78/X fanout60/X _12148_/A _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10534_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13252_ _13254_/CLK _13252_/D vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dfxtp_1
X_10464_ _10461_/Y _10463_/X _11696_/A vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _13185_/CLK _13183_/D vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__dfxtp_1
X_12203_ _12203_/A _12203_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10395_ _10529_/A _10395_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__or3_1
X_12134_ _06559_/Y _12132_/Y _12133_/X vssd1 vssd1 vccd1 vccd1 _12134_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07430__B1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13096__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12065_ hold265/A _12304_/B1 _12126_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _12066_/B
+ sky130_fd_sc_hd__a31o_1
X_11016_ _11155_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11230_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08930__B1 _07842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ _12967_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08289__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12898_ _13085_/A hold129/X vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__and2_1
X_11918_ _11918_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11918_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08219__A _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ _11849_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07123__A _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A1 _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06962__A _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07040_ _07041_/A _07041_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07421__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08889__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08991_ _08870_/A _08991_/B _09049_/A vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__nand3b_1
X_07942_ _07942_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__xnor2_1
X_07873_ _11183_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__xnor2_2
X_06824_ _08983_/B _06823_/A _06823_/B _06545_/A vssd1 vssd1 vccd1 vccd1 _06824_/X
+ sky130_fd_sc_hd__a31o_1
X_09612_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09771_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08921__B1 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ _10009_/A _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__nand3b_1
XANTENNA_fanout261_A _06848_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06755_ _06753_/B _06752_/Y _06753_/Y vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__11808__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _10809_/A _09473_/A _09159_/Y vssd1 vssd1 vccd1 vccd1 _09474_/X sky130_fd_sc_hd__o21a_1
X_06686_ reg1_val[12] _07278_/A vssd1 vssd1 vccd1 vccd1 _06687_/B sky130_fd_sc_hd__or2_1
XANTENNA__12874__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ _08416_/A _08414_/X _08475_/A _08412_/A vssd1 vssd1 vccd1 vccd1 _08427_/C
+ sky130_fd_sc_hd__a211o_1
X_08356_ _08353_/A _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08357_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _11183_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07380_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06591__B _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _08670_/A2 _08689_/B1 _12686_/A _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08288_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07238_ _10156_/A _11184_/B vssd1 vssd1 vccd1 vccd1 _07238_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07169_ _08698_/A _07169_/B vssd1 vssd1 vccd1 vccd1 _07174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10181_/B sky130_fd_sc_hd__xnor2_4
Xfanout241 _12302_/A vssd1 vssd1 vccd1 vccd1 _11696_/A sky130_fd_sc_hd__buf_4
Xfanout263 _12271_/S vssd1 vssd1 vccd1 vccd1 _12125_/S sky130_fd_sc_hd__buf_4
XANTENNA__07208__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 _07050_/A vssd1 vssd1 vccd1 vccd1 _07128_/A sky130_fd_sc_hd__buf_4
Xfanout252 _08765_/A vssd1 vssd1 vccd1 vccd1 _08813_/A1 sky130_fd_sc_hd__buf_6
Xfanout296 fanout298/X vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__buf_4
Xfanout285 _06527_/X vssd1 vssd1 vccd1 vccd1 _06754_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__07715__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ hold292/A hold29/X vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07191__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ hold1/X hold287/A vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07479__B1 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11703_ _13180_/Q _11781_/B _11779_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _11703_/X
+ sky130_fd_sc_hd__a31o_1
X_12683_ _07123_/Y _12926_/A2 hold75/X _12970_/A vssd1 vssd1 vccd1 vccd1 _13134_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ curr_PC[19] _11633_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08691__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11565_ _11654_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08443__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11496_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__or2_1
X_10516_ _11470_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10517_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13235_ _13251_/CLK _13235_/D vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10447_ _10447_/A _10447_/B _10447_/C _10319_/X vssd1 vssd1 vccd1 vccd1 _10449_/C
+ sky130_fd_sc_hd__or4b_2
X_13166_ _13169_/CLK _13166_/D vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__dfxtp_1
X_10378_ _12089_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13097_ hold293/X _06858_/B _13096_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 _13098_/B
+ sky130_fd_sc_hd__a22o_1
X_12117_ _12117_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _12047_/A _12047_/B _12113_/A vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07706__B2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07182__A2 _07187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _06753_/B _06540_/B vssd1 vssd1 vccd1 vccd1 _06540_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13007__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12694__A _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09479__S _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ fanout79/X _08737_/A2 _08733_/B1 _08430_/B vssd1 vssd1 vccd1 vccd1 _08211_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _08901_/A _08901_/B _08904_/A vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11569__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08141_ _08137_/A _08137_/B _08148_/A vssd1 vssd1 vccd1 vccd1 _08143_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07300__B _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ _08814_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08074_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _07023_/A _07023_/B vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _08975_/B _08975_/A vssd1 vssd1 vccd1 vccd1 _08974_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _07925_/A _07925_/B vssd1 vssd1 vccd1 vccd1 _08012_/B sky130_fd_sc_hd__xor2_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ _07859_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _07856_/Y sky130_fd_sc_hd__nor2_1
X_06807_ _11988_/A _06806_/Y _06805_/Y vssd1 vssd1 vccd1 vccd1 _06807_/X sky130_fd_sc_hd__o21a_1
X_07787_ _10117_/A fanout42/X _08333_/B _12684_/A vssd1 vssd1 vccd1 vccd1 _07788_/B
+ sky130_fd_sc_hd__o22a_1
X_06738_ _07051_/A _07108_/C vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09527_/B _09526_/B vssd1 vssd1 vccd1 vccd1 _09528_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_93_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ _09458_/B _09458_/A vssd1 vssd1 vccd1 vccd1 _09457_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08122__A1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06669_ _11143_/S _06669_/B vssd1 vssd1 vccd1 vccd1 _06831_/A sky130_fd_sc_hd__nand2_2
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _09389_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__A1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _08606_/A2 _08735_/A2 _08735_/B1 _08642_/B vssd1 vssd1 vccd1 vccd1 _08340_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ hold179/A _11781_/B _11445_/B _11349_/Y _11448_/A vssd1 vssd1 vccd1 vccd1
+ _11350_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ _13020_/A _13020_/B vssd1 vssd1 vccd1 vccd1 _13020_/Y sky130_fd_sc_hd__xnor2_1
X_11281_ _11739_/A fanout14/X fanout52/X fanout64/X vssd1 vssd1 vccd1 vccd1 _11282_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07936__A1 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _10232_/A _10232_/B _10232_/C vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__and3_1
XANTENNA__07936__B2 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ _10162_/A _10162_/B _10162_/C vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__a21oi_1
X_10094_ _10354_/C _10093_/Y _11153_/A _10091_/X vssd1 vssd1 vccd1 vccd1 dest_val[6]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09153__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ _13019_/B _13020_/A _12765_/X vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06927__D _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10996_ _10868_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12735_ hold81/X hold293/X vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__and2b_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ hold33/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07872__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11617_/Y sky130_fd_sc_hd__xnor2_1
X_12597_ _12597_/A _12599_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06678__A_N _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ _11164_/A _11164_/B _11418_/Y _11547_/X vssd1 vssd1 vccd1 vccd1 _11600_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10759__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ _11480_/A _11480_/B vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13218_ _13222_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08232__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10481__B fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13149_ _13246_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12133__C1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ _12710_/A _09422_/A _09222_/B2 _12712_/A vssd1 vssd1 vccd1 vccd1 _07711_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08690_ _08814_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__xnor2_1
X_07641_ _07641_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11239__A1 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _07572_/A _07572_/B _07572_/C vssd1 vssd1 vccd1 vccd1 _07573_/B sky130_fd_sc_hd__or3_1
XANTENNA__12201__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _09309_/X _09310_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__mux2_1
X_06523_ instruction[3] _06524_/B vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__nor2_8
XANTENNA__10002__A _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12987__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07863__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ _09309_/S _12280_/A _06907_/A _09172_/X vssd1 vssd1 vccd1 vccd1 _09173_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10214__A2 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout224_A _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _08606_/A2 _09180_/B2 _10506_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08125_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _08670_/A2 _09180_/B2 _10506_/A _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08056_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ reg1_val[5] _07006_/B vssd1 vssd1 vccd1 vccd1 _07006_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07918__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08957_ _07585_/A _07585_/B _07583_/X vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07908_ _08741_/A _07908_/B _07908_/C vssd1 vssd1 vccd1 vccd1 _07909_/C sky130_fd_sc_hd__nand3_1
X_08888_ _10117_/A fanout13/X fanout47/X _12684_/A vssd1 vssd1 vccd1 vccd1 _08889_/B
+ sky130_fd_sc_hd__o22a_1
X_07839_ _07839_/A _07839_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_79_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ _10850_/A _10850_/B _10850_/C vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09701__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _09152_/Y _09500_/Y _09501_/Y _09508_/X vssd1 vssd1 vccd1 vccd1 _09509_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11950__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10781_ _10781_/A _10781_/B vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12519_/A _12516_/Y _12518_/B vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__o21a_2
X_12451_ _12496_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12453_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07221__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11404_/C sky130_fd_sc_hd__xnor2_1
X_12382_ _12382_/A _12382_/B _12382_/C vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11953__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _11331_/X _11332_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _11333_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _11713_/A _11261_/X _11262_/Y _11263_/X vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__08052__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__B1 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _13013_/A hold280/X vssd1 vssd1 vccd1 vccd1 _13231_/D sky130_fd_sc_hd__and2_1
XANTENNA__12902__A1 _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _06830_/D _09501_/B _09148_/X _06719_/B _10214_/Y vssd1 vssd1 vccd1 vccd1
+ _10215_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11166__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11195_ _11799_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11196_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _10146_/A _10146_/B _10146_/C vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__or3_1
X_10077_ hold222/A hold239/A _10077_/C vssd1 vssd1 vccd1 vccd1 _10207_/B sky130_fd_sc_hd__or3_1
XANTENNA__12302__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__A1 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__B2 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12969__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06954__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ fanout17/X fanout42/X _07239_/A fanout9/A vssd1 vssd1 vccd1 vccd1 _10980_/B
+ sky130_fd_sc_hd__o22a_1
X_12718_ _12718_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09330__B _09330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12197__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ reg1_val[30] _12656_/A vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__or2_1
XFILLER_0_5_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06970__A _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _06977_/A _07070_/Y fanout17/X _06985_/A vssd1 vssd1 vccd1 vccd1 _09861_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09789_/X _09790_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09794_/B sky130_fd_sc_hd__mux2_1
X_08811_ _08811_/A _08811_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__xor2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08763_/A _08763_/B _08738_/X vssd1 vssd1 vccd1 vccd1 _08743_/C sky130_fd_sc_hd__o21bai_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _08741_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__xnor2_1
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout174_A _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09224__C _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07555_ _12085_/A _07555_/B vssd1 vssd1 vccd1 vccd1 _07559_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09825__A1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__inv_2
X_07486_ _11068_/A _07486_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07836__B1 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _07075_/A _07075_/B _08798_/B vssd1 vssd1 vccd1 vccd1 _09227_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ reg1_val[31] _09156_/B vssd1 vssd1 vccd1 vccd1 _09165_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09087_ _09083_/X _09086_/X _09479_/S vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__mux2_1
X_08107_ fanout83/X _08715_/A2 _08689_/B1 _08565_/B vssd1 vssd1 vccd1 vccd1 _08108_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08038_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08042_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout87_A _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__xor2_4
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08600__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__S _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10123__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11882_ _12094_/A _12141_/A fanout45/X _12148_/A vssd1 vssd1 vccd1 vccd1 _11883_/B
+ sky130_fd_sc_hd__o22a_1
X_10902_ _10902_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10904_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__09816__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ curr_PC[12] _10719_/C _11636_/S vssd1 vssd1 vccd1 vccd1 _10833_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09150__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ _10764_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__and2_1
XFILLER_0_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _12501_/Y _12503_/B vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08047__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__and2_1
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12434_ _12439_/B _12434_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12365_ _12532_/B _12365_/B vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__or2_1
X_11316_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11139__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12296_ _12115_/A _06823_/Y _12295_/Y vssd1 vssd1 vccd1 vccd1 _12297_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _12125_/S _11247_/B vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__or2_1
XANTENNA__08004__B1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11280_/A _11178_/B vssd1 vssd1 vccd1 vccd1 _11180_/C sky130_fd_sc_hd__nand2_1
X_10129_ _10128_/B _10128_/C _10128_/A vssd1 vssd1 vccd1 vccd1 _10130_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11862__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06965__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07340_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07340_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09060__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10417__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__C_N _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07271_ _09634_/A _07271_/B vssd1 vssd1 vccd1 vccd1 _07271_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09010_ _09010_/A _09010_/B _09013_/A vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__or3_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13119__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A2 _07070_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09991__B1 _07157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__nor2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _11654_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09845_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout291_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11550__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06982_/A _07065_/A _07028_/C _07058_/B1 vssd1 vssd1 vccd1 vccd1 _06987_/B
+ sky130_fd_sc_hd__o31a_1
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _11163_/A sky130_fd_sc_hd__nand2_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _08706_/B _08706_/C _08706_/A vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_96_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08656_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__and2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _07608_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _07607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09251__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ _08588_/B _08588_/C _08588_/A vssd1 vssd1 vccd1 vccd1 _08587_/X sky130_fd_sc_hd__o21a_1
X_07538_ _07538_/A _07538_/B vssd1 vssd1 vccd1 vccd1 _07546_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ _07542_/B _07542_/A vssd1 vssd1 vccd1 vccd1 _07469_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11081__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ _09209_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10480_ _10434_/A _10434_/B _10435_/Y vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09139_ _09146_/A _09140_/B vssd1 vssd1 vccd1 vccd1 _09139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08785__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _12208_/B _12150_/B vssd1 vssd1 vccd1 vccd1 _12152_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ _11102_/A _11102_/B _11102_/C vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__a21oi_1
X_12081_ _12078_/Y _12080_/X _12080_/A _12077_/X vssd1 vssd1 vccd1 vccd1 dest_val[26]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11956__A _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11032_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08330__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ hold294/X _06858_/B _12982_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold295/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11934_ _06579_/A _09141_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ curr_PC[22] _11866_/C curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__a21oi_1
X_10816_ _12125_/S _10810_/Y _10813_/X _10815_/Y vssd1 vssd1 vccd1 vccd1 _10816_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11796_ _11796_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ _10747_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _10680_/A vssd1 vssd1 vccd1 vccd1 _10794_/C sky130_fd_sc_hd__inv_2
XFILLER_0_125_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12417_ _12417_/A _12417_/B _12417_/C vssd1 vssd1 vccd1 vccd1 _12418_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12348_ _12354_/B _12348_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ _09138_/X _12278_/X _06572_/B vssd1 vssd1 vccd1 vccd1 _12280_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09336__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B1 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ instruction[6] _12297_/A _09146_/A vssd1 vssd1 vccd1 vccd1 _06840_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06679__B _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _06730_/Y _06770_/Y _06832_/A vssd1 vssd1 vccd1 vccd1 _06772_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12088__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A1 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11835__A1 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ _08510_/A _08510_/B vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10099__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08498_/A _08498_/B _08437_/Y vssd1 vssd1 vccd1 vccd1 _08452_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08417_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09256__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10010__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07323_ _07110_/Y _07154_/X _07799_/B _07147_/Y vssd1 vssd1 vccd1 vccd1 _07324_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _06585_/B _06592_/B _07068_/A _07303_/A vssd1 vssd1 vccd1 vccd1 _07255_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA_fanout137_A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07185_ _09479_/S _07186_/B vssd1 vssd1 vccd1 vccd1 _07185_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__08767__A1 _08768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _11796_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__xnor2_1
X_06969_ _10252_/A vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__inv_6
X_09757_ _09757_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__nor2_2
XANTENNA__12400__A _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08709_/B sky130_fd_sc_hd__and2_1
XANTENNA__10629__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09688_ _09689_/B _09689_/A vssd1 vssd1 vccd1 vccd1 _09688_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08639_ _08640_/A _08657_/A _08640_/C vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11039__C1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 _12095_/B vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__clkbuf_8
X_11650_ _11650_/A _11650_/B vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout41 _07287_/X vssd1 vssd1 vccd1 vccd1 fanout41/X sky130_fd_sc_hd__buf_8
Xfanout74 _12710_/A vssd1 vssd1 vccd1 vccd1 fanout74/X sky130_fd_sc_hd__clkbuf_4
Xfanout63 _12720_/A vssd1 vssd1 vccd1 vccd1 fanout63/X sky130_fd_sc_hd__buf_4
Xfanout52 _07513_/B vssd1 vssd1 vccd1 vccd1 fanout52/X sky130_fd_sc_hd__buf_6
X_11581_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__and2_1
XFILLER_0_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _10555_/A _10555_/B _10553_/X vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11054__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout85 _09621_/A vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout96 _12142_/A vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__buf_8
X_10532_ _10532_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08325__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13251_ _13251_/CLK _13251_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
X_10463_ _10087_/X _10462_/X _11135_/S vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08758__A1 _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ _13185_/CLK _13182_/D vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10565__A1 _10681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _07075_/A _07075_/B _08565_/B vssd1 vssd1 vccd1 vccd1 _10395_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12133_ _07064_/B _12238_/C1 _09147_/X _06560_/A _06847_/X vssd1 vssd1 vccd1 vccd1
+ _12133_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07430__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07430__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _12304_/B1 _12126_/B hold265/A vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09707__B1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _10796_/B _11156_/A _11158_/A vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10317__A1 _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ _12970_/A hold250/X vssd1 vssd1 vccd1 vccd1 _13223_/D sky130_fd_sc_hd__and2_1
X_12897_ _13189_/Q _13084_/B2 _13084_/A2 hold128/X vssd1 vssd1 vccd1 vccd1 hold129/A
+ sky130_fd_sc_hd__a22o_1
X_11917_ _06798_/X _11916_/X _12263_/S vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08219__B _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11769_/Y _11773_/B _11771_/B vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__A1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _13180_/Q _11779_/B vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07421__A1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__B2 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ _08991_/B _09049_/A _08870_/A vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07941_ _07942_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07941_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09174__A1 _09173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _09698_/A fanout37/X _08233_/B _09885_/A vssd1 vssd1 vccd1 vccd1 _07873_/B
+ sky130_fd_sc_hd__o22a_1
X_06823_ _06823_/A _06823_/B vssd1 vssd1 vccd1 vccd1 _06823_/Y sky130_fd_sc_hd__nand2_1
X_09611_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08921__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A1 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06754_ reg2_val[1] _06754_/B vssd1 vssd1 vccd1 vccd1 _06754_/X sky130_fd_sc_hd__and2_1
XANTENNA__11808__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ _10607_/A _09542_/B vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11808__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ _09473_/A vssd1 vssd1 vccd1 vccd1 _09473_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout254_A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ reg1_val[12] _07278_/A vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__and2_1
XANTENNA__10492__B1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07306_ _12688_/A fanout36/X _12690_/A _07305_/X vssd1 vssd1 vccd1 vccd1 _07307_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08286_ _08688_/A _08286_/B vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__xnor2_1
X_07237_ _07237_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _10845_/C sky130_fd_sc_hd__nand2_1
X_07168_ _12710_/A _10009_/A _12712_/A _09725_/B2 vssd1 vssd1 vccd1 vccd1 _07169_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07099_ _07099_/A _07099_/B vssd1 vssd1 vccd1 vccd1 _07099_/X sky130_fd_sc_hd__xor2_2
Xfanout220 _06856_/Y vssd1 vssd1 vccd1 vccd1 _13084_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout231 _09634_/A vssd1 vssd1 vccd1 vccd1 _10201_/S sky130_fd_sc_hd__buf_4
Xfanout242 _06727_/X vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__buf_4
Xfanout264 _06726_/X vssd1 vssd1 vccd1 vccd1 _12271_/S sky130_fd_sc_hd__clkbuf_4
Xfanout253 _07063_/Y vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__clkbuf_8
Xfanout297 fanout298/X vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__clkbuf_2
X_09809_ _09808_/B _10080_/C hold294/A vssd1 vssd1 vccd1 vccd1 _09810_/C sky130_fd_sc_hd__a21oi_1
Xfanout286 _06753_/B vssd1 vssd1 vccd1 vccd1 _06763_/B sky130_fd_sc_hd__buf_6
Xfanout275 _06908_/X vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__buf_4
XANTENNA__07715__A2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _13072_/B _13073_/A _12746_/X vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ hold166/X hold283/A vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07479__A1 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07479__B2 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ hold74/X _12686_/B vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__or2_1
X_11702_ _11781_/B _11779_/B _13180_/Q vssd1 vssd1 vccd1 vccd1 _11702_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ curr_PC[19] curr_PC[20] _11633_/C vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__and3_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08428__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11432__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ _11564_/A fanout3/X vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ _11402_/A _11402_/B _11400_/Y vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__a21boi_1
X_10515_ _11663_/A fanout41/X _08135_/B _11739_/A vssd1 vssd1 vccd1 vccd1 _10516_/B
+ sky130_fd_sc_hd__o22a_1
X_13234_ _13234_/CLK _13234_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
X_10446_ _10560_/B _10446_/B vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11735__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13165_ _13169_/CLK hold215/X vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
X_10377_ _10377_/A1 fanout44/X fanout92/X fanout11/X vssd1 vssd1 vccd1 vccd1 _10378_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13096_ hold275/X _13095_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__mux2_1
X_12116_ _12053_/A _12114_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__a21oi_1
X_12047_ _12047_/A _12047_/B vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07706__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ hold92/X _12665_/A _12955_/B1 hold106/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold109/A sky130_fd_sc_hd__o221a_1
XFILLER_0_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12694__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06692__B _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10226__B1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07300__C _07301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ _08274_/A _11462_/A _08813_/A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 _08072_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _07023_/A _07023_/B vssd1 vssd1 vccd1 vccd1 _07216_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_24_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08973_ _08973_/A _08973_/B vssd1 vssd1 vccd1 vccd1 _08975_/B sky130_fd_sc_hd__xnor2_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__B _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07924_ _08734_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _08012_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _07855_/A _07855_/B vssd1 vssd1 vccd1 vccd1 _07859_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06806_ reg1_val[24] _07029_/B vssd1 vssd1 vccd1 vccd1 _06806_/Y sky130_fd_sc_hd__nand2_1
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__nor2_1
X_06737_ _06763_/B _06646_/A _12522_/B _06735_/X vssd1 vssd1 vccd1 vccd1 _06737_/Y
+ sky130_fd_sc_hd__a31oi_4
X_09525_ _11794_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08658__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06668_ reg1_val[15] _06941_/A vssd1 vssd1 vccd1 vccd1 _06669_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08122__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08407_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__xnor2_1
X_06599_ reg2_val[23] _06754_/B _06657_/B1 _06598_/X vssd1 vssd1 vccd1 vccd1 _06601_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09387_ _09387_/A _09387_/B vssd1 vssd1 vccd1 vccd1 _09389_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08338_ _08328_/Y _08332_/X _08336_/X _08337_/Y vssd1 vssd1 vccd1 vccd1 _08350_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08269_ _08223_/B _08223_/C _08223_/A vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11280_ _11280_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__xnor2_1
X_10300_ _10300_/A _10300_/B vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11717__B1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _10232_/A _10232_/B _10232_/C vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07219__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _10162_/A _10162_/B _10162_/C vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__and3_1
XANTENNA__10940__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ curr_PC[6] _10092_/B _11636_/S vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12693__A1 _07277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12498__C _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _13014_/B _13015_/A _12767_/X vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ _12832_/B _12734_/B vssd1 vssd1 vccd1 vccd1 _13104_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10995_ _10885_/A _10885_/B _10884_/A vssd1 vssd1 vccd1 vccd1 _11000_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07872__A1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11616_ _11523_/Y _11527_/B _11525_/B vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__o21a_1
X_12596_ reg1_val[19] _12615_/B vssd1 vssd1 vccd1 vccd1 _12599_/C sky130_fd_sc_hd__xnor2_4
XANTENNA__10759__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10759__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _11799_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11480_/B sky130_fd_sc_hd__xnor2_1
X_13217_ _13217_/CLK _13217_/D vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__or2_1
X_13148_ _13243_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ hold271/X _13084_/A2 _13078_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold272/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12133__B1 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08888__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _07640_/A _07640_/B vssd1 vssd1 vccd1 vccd1 _07641_/B sky130_fd_sc_hd__nor2_1
X_07571_ _07572_/A _07572_/B _07572_/C vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12987__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06522_ instruction[0] instruction[1] _06850_/B pred_val vssd1 vssd1 vccd1 vccd1
+ _06524_/B sky130_fd_sc_hd__or4bb_4
X_09310_ _09098_/X _09100_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09310_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07799__A _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07863__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__B2 _06939_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09241_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ _06824_/X _06905_/B _09171_/X vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08123_ _08714_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08050_/A _08050_/B _08239_/A vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07005_ reg1_val[4] _07050_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _07006_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09519__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _08956_/A _08956_/B vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__xor2_1
X_07907_ _07908_/B _07908_/C _08741_/A vssd1 vssd1 vccd1 vccd1 _07909_/B sky130_fd_sc_hd__a21o_1
X_08887_ _08890_/A vssd1 vssd1 vccd1 vccd1 _08887_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _07839_/A _07839_/B vssd1 vssd1 vccd1 vccd1 _07838_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ reg1_val[2] _09634_/A _09147_/X _09504_/X _09505_/X vssd1 vssd1 vccd1 vccd1
+ _09508_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07769_ _06940_/A fanout92/X _10647_/A fanout82/X vssd1 vssd1 vccd1 vccd1 _07770_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10781_/A _10781_/B vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09440_/B sky130_fd_sc_hd__nand2_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ reg1_val[20] curr_PC[20] _12495_/S vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__mux2_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11959__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _12382_/A _12382_/B _12382_/C vssd1 vssd1 vccd1 vccd1 _12389_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08333__A _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ _11233_/A _12110_/A _11232_/A vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11263_ curr_PC[16] _11265_/C _11636_/S vssd1 vssd1 vccd1 vccd1 _11263_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09359__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__A1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13002_ hold279/X _12663_/B _13001_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold280/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12902__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ _06719_/A _12309_/B1 _10213_/X vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11166__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11194_ fanout64/X fanout13/X fanout47/X _11876_/A vssd1 vssd1 vccd1 vccd1 _11195_/B
+ sky130_fd_sc_hd__o22a_1
X_10145_ _10275_/B _10144_/B _10144_/C vssd1 vssd1 vccd1 vccd1 _10146_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ _10067_/Y _10075_/Y _11696_/A vssd1 vssd1 vccd1 vccd1 _10076_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11469__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12969__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11626__C1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10978_ _11065_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ hold29/X _12720_/B _12716_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11641__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06954__C _06961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12648_ _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ _12579_/A _12579_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
XANTENNA__08270__A1 _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08270__B2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08810_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09087_/X _09110_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09790_/X sky130_fd_sc_hd__mux2_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08741_/A _08741_/B vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__xor2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08672_ _08755_/B _08737_/A2 _08813_/B1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 _08673_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11163__D_N _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07623_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout167_A _07056_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ fanout15/X _09698_/A _07513_/B _09885_/A vssd1 vssd1 vccd1 vccd1 _07555_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ hold251/X vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__inv_2
X_07485_ _10117_/A fanout36/X fanout34/X _07137_/Y vssd1 vssd1 vccd1 vccd1 _07486_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07836__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _09224_/A _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ _09155_/A _09155_/B vssd1 vssd1 vccd1 vccd1 _09155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _09084_/X _09085_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08106_ _08110_/A vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__inv_2
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08037_ _08037_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08860_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07992__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__nand2_1
X_08939_ _12029_/B _08939_/B vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ _11950_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__nor2_1
X_10901_ _10902_/B _10902_/A vssd1 vssd1 vccd1 vccd1 _10901_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10123__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _11803_/A _11879_/B _11802_/B _11806_/A vssd1 vssd1 vccd1 vccd1 _11897_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10832_ curr_PC[11] curr_PC[12] _10832_/C vssd1 vssd1 vccd1 vccd1 _11051_/C sky130_fd_sc_hd__and3_2
XFILLER_0_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _10764_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ reg1_val[1] _12502_/B vssd1 vssd1 vccd1 vccd1 _12503_/B sky130_fd_sc_hd__or2_2
XFILLER_0_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10831__B1 _10830_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12433_ _12496_/A _12427_/B _12439_/A vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12364_ _12532_/B _12365_/B vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08063__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _11214_/A _11214_/B _11213_/A vssd1 vssd1 vccd1 vccd1 _11317_/B sky130_fd_sc_hd__a21o_1
X_12295_ _12264_/A _12262_/X _12115_/A _12278_/S vssd1 vssd1 vccd1 vccd1 _12295_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__08004__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11246_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11246_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08004__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _11177_/A _11177_/B vssd1 vssd1 vccd1 vccd1 _11178_/B sky130_fd_sc_hd__or2_1
X_10128_ _10128_/A _10128_/B _10128_/C vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nand3_1
X_10059_ instruction[7] _10059_/B vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09504__A1 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ _09634_/A _07271_/B vssd1 vssd1 vccd1 vccd1 _07270_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13119__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09911_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _10310_/A sky130_fd_sc_hd__and2_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12223__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _10099_/A1 _11564_/A fanout38/X _10359_/B2 vssd1 vssd1 vccd1 vccd1 _09843_/B
+ sky130_fd_sc_hd__o22a_1
X_09773_ _09460_/Y _09774_/B _09772_/Y vssd1 vssd1 vccd1 vccd1 _09773_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11550__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11550__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08724_ _08726_/A _08726_/B _08726_/C vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__a21o_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _06985_/A vssd1 vssd1 vccd1 vccd1 _08700_/C sky130_fd_sc_hd__inv_2
XANTENNA__06875__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08655_ _08655_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__xor2_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _09420_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07608_/B sky130_fd_sc_hd__xnor2_2
X_08586_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08588_/C sky130_fd_sc_hd__and2b_1
XANTENNA__07052__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07468_ _07468_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07399_ _07396_/A _07395_/B _07395_/A vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ _09209_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__or2_1
X_09138_ _09153_/B _09142_/B vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__or2_4
XANTENNA__08234__A1 _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08785__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ reg1_val[3] reg1_val[28] _09092_/S vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _11065_/A _10978_/B _10986_/B _10989_/A vssd1 vssd1 vccd1 vccd1 _11102_/C
+ sky130_fd_sc_hd__o31a_1
X_12080_ _12080_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__or2_1
XANTENNA__08611__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11031_ _10923_/A _10923_/B _10921_/B vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10344__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ hold257/X _12981_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__mux2_1
X_11933_ hold271/A _11623_/B _11998_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11933_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _06601_/B _06905_/Y _06907_/Y _11863_/X vssd1 vssd1 vccd1 vccd1 _11864_/X
+ sky130_fd_sc_hd__o22a_1
X_10815_ _12125_/S _10815_/B vssd1 vssd1 vccd1 vccd1 _10815_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08058__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _11796_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _11879_/A sky130_fd_sc_hd__or2_1
XANTENNA__10804__B1 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ _11799_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10747_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10677_ _10677_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__or2_2
X_12416_ _12417_/A _12417_/B _12417_/C vssd1 vssd1 vccd1 vccd1 _12424_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12309__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _12347_/A _12347_/B _12347_/C vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _09501_/B _09148_/X _12278_/S vssd1 vssd1 vccd1 vccd1 _12278_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08521__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _11229_/A _11418_/A vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09725__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07137__A _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _09924_/B _09924_/C _09926_/A vssd1 vssd1 vccd1 vccd1 _06770_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__12088__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10498__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__B2 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _08440_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08996_/A _08995_/A _09043_/A _08998_/A vssd1 vssd1 vccd1 vccd1 _08371_/Y
+ sky130_fd_sc_hd__nand4_1
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07337_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ _09862_/B _07253_/B vssd1 vssd1 vccd1 vccd1 _07259_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07184_ _09495_/A _07184_/B _09309_/S vssd1 vssd1 vccd1 vccd1 _07186_/B sky130_fd_sc_hd__and3_2
XFILLER_0_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08767__A2 _08768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09413__B1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09825_ _10490_/B2 fanout51/X fanout49/X fanout80/X vssd1 vssd1 vccd1 vccd1 _09826_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06968_ reg1_val[9] _06968_/B vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__06950__A1 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _09577_/A _09577_/B _09575_/Y vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__a21o_2
X_08707_ _08707_/A _08731_/A vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__xor2_1
X_09687_ _09687_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09689_/B sky130_fd_sc_hd__xnor2_1
X_06899_ _12080_/A _06899_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08638_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _08640_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout20 _09465_/A vssd1 vssd1 vccd1 vccd1 _11838_/A sky130_fd_sc_hd__buf_4
Xfanout31 _12095_/B vssd1 vssd1 vccd1 vccd1 _11885_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__xor2_1
Xfanout53 _07112_/Y vssd1 vssd1 vccd1 vccd1 _07513_/B sky130_fd_sc_hd__buf_6
Xfanout64 _12714_/A vssd1 vssd1 vccd1 vccd1 fanout64/X sky130_fd_sc_hd__buf_6
X_11580_ _11668_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout42 fanout43/X vssd1 vssd1 vccd1 vccd1 fanout42/X sky130_fd_sc_hd__clkbuf_8
X_10600_ _11636_/S _10596_/X _10599_/X vssd1 vssd1 vccd1 vccd1 dest_val[10] sky130_fd_sc_hd__o21ai_4
Xfanout86 _11235_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__clkbuf_4
Xfanout75 _06987_/Y vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__clkbuf_8
Xfanout97 _12142_/A vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__buf_8
XANTENNA_fanout9_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ _10531_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__and2_1
X_13250_ _13250_/CLK _13250_/D vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ _09307_/X _09315_/X _10924_/S vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__mux2_1
X_12201_ _12201_/A _12245_/B _12142_/A vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13181_ _13185_/CLK hold193/X vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09955__A1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10871__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10393_ _10393_/A _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__and3_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ _06560_/A _09501_/B _09138_/X vssd1 vssd1 vccd1 vccd1 _12132_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07430__A2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ hold299/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__or2_1
XANTENNA__09156__B _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11156_/A sky130_fd_sc_hd__and2_1
XANTENNA__08930__A2 _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12965_ _12664_/A _12963_/Y _12964_/X _12663_/B hold249/X vssd1 vssd1 vccd1 vccd1
+ hold250/A sky130_fd_sc_hd__a32o_1
X_11916_ _06837_/A _11841_/X _11858_/S vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12896_ _13085_/A hold175/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11847_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ hold291/A _11623_/B _11931_/C _11777_/Y _12313_/A1 vssd1 vssd1 vccd1 vccd1
+ _11778_/X sky130_fd_sc_hd__a311o_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09643__B1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _11271_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12071__A2_N _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13250_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__07421__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _07942_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07871_ _07932_/A _07932_/B _07867_/X vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__08382__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ _06821_/A _06821_/B _12264_/A vssd1 vssd1 vccd1 vccd1 _06823_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08921__A2 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _09610_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09613_/C sky130_fd_sc_hd__xnor2_1
X_06753_ reg2_val[1] _06753_/B vssd1 vssd1 vccd1 vccd1 _06753_/Y sky130_fd_sc_hd__nor2_1
X_09541_ _10481_/A fanout58/X fanout55/X _07000_/A vssd1 vssd1 vccd1 vccd1 _09542_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11808__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ _11134_/S _09471_/Y _09166_/B vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__o21a_1
X_06684_ _07278_/A reg1_val[12] vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09882__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__C _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__or2_1
XANTENNA__10492__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07305_ _07305_/A _11385_/A vssd1 vssd1 vccd1 vccd1 _07305_/X sky130_fd_sc_hd__or2_4
XFILLER_0_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ _12694_/A _08798_/B fanout93/X _09727_/A vssd1 vssd1 vccd1 vccd1 _08286_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _07237_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07236_/X sky130_fd_sc_hd__and2_1
X_07167_ _07832_/A _07167_/B vssd1 vssd1 vccd1 vccd1 _07174_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07948__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09257__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ _07099_/A _07099_/B vssd1 vssd1 vccd1 vccd1 _07098_/Y sky130_fd_sc_hd__xnor2_2
Xfanout221 _06858_/B vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__buf_4
Xfanout210 _08688_/A vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__buf_12
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout232 _09634_/A vssd1 vssd1 vccd1 vccd1 _10073_/S sky130_fd_sc_hd__clkbuf_8
Xfanout243 _06539_/X vssd1 vssd1 vccd1 vccd1 _06657_/B1 sky130_fd_sc_hd__buf_8
Xfanout265 _06613_/A vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__buf_6
Xfanout254 _09420_/A vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__buf_12
Xfanout298 _06521_/Y vssd1 vssd1 vccd1 vccd1 fanout298/X sky130_fd_sc_hd__clkbuf_4
Xfanout276 _12484_/A vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__buf_8
X_09808_ hold294/A _09808_/B _10080_/C vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__and3_1
Xfanout287 _06526_/X vssd1 vssd1 vccd1 vccd1 _06753_/B sky130_fd_sc_hd__buf_4
XANTENNA_fanout62_A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _10377_/A1 fanout50/X _07988_/B _10490_/B2 vssd1 vssd1 vccd1 vccd1 _09740_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06923__A1 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ hold263/X hold13/X vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07479__A2 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ hold210/A _11701_/B vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__or2_1
X_12681_ _07157_/X _12926_/A2 hold69/X _12970_/A vssd1 vssd1 vccd1 vccd1 _13133_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10866__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ _09145_/Y _11607_/X _11608_/Y _11631_/Y _11606_/Y vssd1 vssd1 vccd1 vccd1
+ _11632_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08428__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08428__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07100__A1 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _11656_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11567_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ _11494_/A _11494_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__xor2_1
X_10514_ _10514_/A _10514_/B vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__nor2_1
X_13233_ _13260_/CLK _13233_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__and2_1
XFILLER_0_110_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _13169_/CLK hold224/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11735__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11735__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _12115_/A _12115_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__and3_1
X_10376_ _10376_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__xor2_1
X_13095_ _13095_/A _13095_/B vssd1 vssd1 vccd1 vccd1 _13095_/Y sky130_fd_sc_hd__xnor2_1
X_12046_ _11909_/Y _11910_/X _11980_/A _12112_/A vssd1 vssd1 vccd1 vccd1 _12047_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11636__S _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__B1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ _07152_/B _12962_/B2 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o21a_1
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _13180_/Q _12885_/A2 _12885_/B1 hold191/X vssd1 vssd1 vccd1 vccd1 hold192/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07150__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11423__B1 _11235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ _08801_/A _08070_/B vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07021_ _07021_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07023_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10934__C1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08972_ _07652_/A _07652_/B _07650_/Y vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10016__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _11462_/A _09422_/A _08815_/B fanout76/X vssd1 vssd1 vccd1 vccd1 _07924_/B
+ sky130_fd_sc_hd__o22a_1
X_07854_ _07854_/A _07854_/B vssd1 vssd1 vccd1 vccd1 _07859_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06805_ reg1_val[25] _07059_/A vssd1 vssd1 vccd1 vccd1 _06805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07785_ _07785_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__and2_1
XANTENNA__08107__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06736_ _06763_/B _06646_/A _12522_/B _06735_/X vssd1 vssd1 vccd1 vccd1 _06736_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09524_ fanout15/X _12684_/A _10370_/A fanout52/X vssd1 vssd1 vccd1 vccd1 _09525_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08658__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ reg1_val[15] _06941_/A vssd1 vssd1 vccd1 vccd1 _11143_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09455_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09540__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _08394_/X _08405_/X _08350_/B _08376_/X vssd1 vssd1 vccd1 vccd1 _08416_/A
+ sky130_fd_sc_hd__o211ai_2
X_06598_ _06613_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _06598_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ _09387_/A _09387_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08337_ _11072_/A _08408_/A vssd1 vssd1 vccd1 vccd1 _08337_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ _08268_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07995__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07219_ _10252_/A _07219_/B vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13001__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__A _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__B2 _07070_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__A1 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ _08200_/B _08200_/A vssd1 vssd1 vccd1 vccd1 _08199_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10230_ _10371_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10232_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08594__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__xnor2_1
X_10092_ curr_PC[6] _10092_/B vssd1 vssd1 vccd1 vccd1 _10354_/C sky130_fd_sc_hd__and2_1
XANTENNA__12693__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12141__A _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _13009_/B _13010_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__a21o_1
X_10994_ _10880_/B _10886_/B _10880_/A vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__09846__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ _13105_/A hold7/X vssd1 vssd1 vccd1 vccd1 _12734_/B sky130_fd_sc_hd__nand2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12664_ _12664_/A _12664_/B vssd1 vssd1 vccd1 vccd1 _12664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07872__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11615_/A _11615_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__nand2_1
X_12595_ _12591_/A _12594_/B _12591_/B vssd1 vssd1 vccd1 vccd1 _12597_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ _11713_/A _11543_/X _11544_/X _11545_/Y vssd1 vssd1 vccd1 vccd1 dest_val[19]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10759__A2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13216_ _13217_/CLK _13216_/D vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ _12095_/A fanout13/X fanout47/X fanout60/X vssd1 vssd1 vccd1 vccd1 _11478_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _10289_/A _10289_/B _10287_/Y vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ _13254_/CLK _13147_/D vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__dfxtp_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _06946_/X _07154_/X fanout47/X _10359_/B2 vssd1 vssd1 vccd1 vccd1 _10360_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13078_ hold292/A _13077_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__mux2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12029_ _12095_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08888__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__B2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _08897_/A _07570_/B vssd1 vssd1 vccd1 vccd1 _07572_/C sky130_fd_sc_hd__and2_1
X_06521_ rst vssd1 vssd1 vccd1 vccd1 _06521_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07799__B _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07312__B2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ _11885_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07863__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _09062_/Y _09063_/X _09170_/X vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09464__C_N _09617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07076__B1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ _08699_/A2 fanout93/X _10647_/A _08670_/A2 vssd1 vssd1 vccd1 vccd1 _08123_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__nor2_1
X_07004_ _07832_/A _07004_/B vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout112_A _11887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ _11654_/A _08955_/B vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__xnor2_1
X_07906_ _11169_/A _08755_/B vssd1 vssd1 vccd1 vccd1 _07908_/C sky130_fd_sc_hd__or2_1
XANTENNA__12675__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _11883_/A _08886_/B vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12896__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _10252_/A _07837_/B vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07055__A _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _07768_/A _07768_/B _07768_/C vssd1 vssd1 vccd1 vccd1 _07771_/B sky130_fd_sc_hd__nand3_1
X_06719_ _06719_/A _06719_/B vssd1 vssd1 vccd1 vccd1 _06830_/D sky130_fd_sc_hd__nand2_1
X_09507_ _09488_/X _09493_/X _12125_/S vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07699_ _07699_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09438_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ _09370_/A _09370_/B _09370_/C vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _12389_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12382_/C sky130_fd_sc_hd__nand2_1
X_11400_ _11399_/A _11399_/B _11401_/A vssd1 vssd1 vccd1 vccd1 _11400_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__and2_1
XANTENNA__08333__B _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ curr_PC[16] _11265_/C vssd1 vssd1 vccd1 vccd1 _11262_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09359__A2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ hold300/A _13000_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__mux2_1
X_10213_ _10211_/Y _10212_/X _07123_/A _12238_/C1 vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11166__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _11196_/A vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__inv_2
X_10144_ _10275_/B _10144_/B _10144_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__and3_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ _10203_/S _10074_/X _10072_/X vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11874__B1 _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ _12716_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ _12647_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__or2_2
XFILLER_0_26_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12578_ _12578_/A _12578_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__and3_2
XFILLER_0_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11529_ hold182/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__or2_1
XANTENNA__08270__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11885__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06698__B _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08740_ _08755_/A _08740_/A2 _08755_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08741_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _08714_/A _08671_/B vssd1 vssd1 vccd1 vccd1 _08708_/A sky130_fd_sc_hd__xnor2_1
X_07622_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _07622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ _07249_/A _07249_/B _07261_/B _07262_/B _07262_/A vssd1 vssd1 vccd1 vccd1
+ _07567_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__09286__A1 _09464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ hold245/X vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__inv_2
X_07484_ _07484_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07836__A2 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _09564_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09223_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ hold249/A _09150_/Y _09152_/Y hold189/A _09149_/Y vssd1 vssd1 vccd1 vccd1
+ _09155_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08434__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ _10853_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__xnor2_2
X_09085_ reg1_val[12] reg1_val[19] _09092_/S vssd1 vssd1 vccd1 vccd1 _09085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ _08036_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11795__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _10168_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__and2_1
X_08938_ fanout8/X _09428_/A fanout6/X _09237_/A vssd1 vssd1 vccd1 vccd1 _08939_/B
+ sky130_fd_sc_hd__o22a_1
X_08869_ _08870_/B vssd1 vssd1 vccd1 vccd1 _09048_/D sky130_fd_sc_hd__inv_2
XFILLER_0_99_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07513__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _11880_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__or2_1
XANTENNA__08609__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _12179_/A _10800_/Y _10801_/X _10830_/X _10799_/X vssd1 vssd1 vccd1 vccd1
+ _10831_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ _06921_/X _11385_/B _10761_/Y _10850_/A vssd1 vssd1 vccd1 vccd1 _10764_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _12501_/A _12501_/B vssd1 vssd1 vccd1 vccd1 _12501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__A1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12432_ _12496_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12439_/B sky130_fd_sc_hd__xnor2_4
X_10693_ _10692_/A _10692_/B _10692_/Y _09498_/A vssd1 vssd1 vccd1 vccd1 _10715_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ reg1_val[7] curr_PC[7] _12495_/S vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__mux2_1
X_12294_ _12286_/Y _12289_/X _12291_/Y _12293_/X _10450_/A vssd1 vssd1 vccd1 vccd1
+ _12294_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11314_ _11314_/A _11314_/B vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ _11243_/Y _11245_/B vssd1 vssd1 vccd1 vccd1 _11246_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08004__A2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11176_ _11177_/A _11177_/B vssd1 vssd1 vccd1 vccd1 _11280_/A sky130_fd_sc_hd__nand2_1
X_10127_ _10126_/B _10126_/C _10126_/A vssd1 vssd1 vccd1 vccd1 _10128_/C sky130_fd_sc_hd__a21o_1
X_10058_ _06732_/X _09923_/Y _06734_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09504__A2 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A0 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09841_ _09979_/A _09841_/B vssd1 vssd1 vccd1 vccd1 _09845_/A sky130_fd_sc_hd__xnor2_4
X_06984_ _06984_/A _06984_/B vssd1 vssd1 vccd1 vccd1 _06984_/Y sky130_fd_sc_hd__nand2_2
X_09772_ _09457_/Y _09771_/C _09614_/B vssd1 vssd1 vccd1 vccd1 _09772_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11550__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10353__A3 _10332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ _08726_/A _08726_/B _08726_/C vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__a21oi_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08655_/B sky130_fd_sc_hd__or2_1
XANTENNA__10510__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08429__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _08765_/A fanout9/A fanout4/X _06828_/A vssd1 vssd1 vccd1 vccd1 _07606_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08585_ _08588_/B _08585_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__nor2_1
X_07536_ _07536_/A _07536_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ _07675_/A _07502_/B _07460_/X vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _10126_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07398_ _07344_/A _07344_/B _07397_/B _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1
+ _07475_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07690__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__B1 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _09153_/B _09142_/B vssd1 vssd1 vccd1 vccd1 _09137_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07442__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _09066_/X _09067_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08019_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08156_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12414__A _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout92_A fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _11030_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__nand2_1
X_12981_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _12981_/Y sky130_fd_sc_hd__xnor2_1
X_11932_ _11623_/B _11998_/B hold271/A vssd1 vssd1 vccd1 vccd1 _11932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _11836_/Y _11837_/X _11840_/X _12179_/A _11862_/X vssd1 vssd1 vccd1 vccd1
+ _11863_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _10811_/X _10812_/Y _10695_/X _10697_/Y vssd1 vssd1 vccd1 vccd1 _10815_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ _11794_/A _11794_/B vssd1 vssd1 vccd1 vccd1 _11796_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10745_ _11462_/A fanout13/X fanout47/X fanout76/X vssd1 vssd1 vccd1 vccd1 _10746_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12006__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12424_/A _12415_/B vssd1 vssd1 vccd1 vccd1 _12417_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_63_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ _12347_/A _12347_/B _12347_/C vssd1 vssd1 vccd1 vccd1 _12354_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12277_ _13189_/Q _12190_/B _12275_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12277_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09617__B _09617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__C _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _11164_/A _11164_/B _11418_/A vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__09725__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11160_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10099__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07321_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07327_/B sky130_fd_sc_hd__and2_1
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _12095_/A _08798_/B _11950_/A _09727_/A vssd1 vssd1 vccd1 vccd1 _07253_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07183_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__or2_1
XANTENNA__09413__A1 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09413__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _09734_/A _09734_/B _09733_/A vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__a21o_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ reg1_val[7] reg1_val[8] _06970_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _06968_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__10689__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09530_/A _09530_/B _09531_/Y vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__o21ai_4
X_06898_ instruction[24] _09495_/A is_load _06727_/B _06897_/X vssd1 vssd1 vccd1 vccd1
+ _06899_/B sky130_fd_sc_hd__a32o_2
XANTENNA__06950__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _08706_/A _08706_/B _08706_/C vssd1 vssd1 vccd1 vccd1 _08706_/X sky130_fd_sc_hd__and3_1
X_09686_ _09538_/A _09538_/B _09536_/Y vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__a21oi_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08637_ _08656_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07063__A _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06526__B_N _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout21 _09465_/A vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__buf_2
Xfanout10 _12728_/A vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__buf_6
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ _08603_/B _08535_/A _08603_/A vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ _11955_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout54 _12718_/A vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__clkbuf_8
Xfanout32 _07576_/Y vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__clkbuf_8
Xfanout65 _12714_/A vssd1 vssd1 vccd1 vccd1 fanout65/X sky130_fd_sc_hd__buf_4
X_08499_ _08502_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _08503_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10798__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout43 _07236_/X vssd1 vssd1 vccd1 vccd1 fanout43/X sky130_fd_sc_hd__buf_8
XFILLER_0_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout87 _12690_/A vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__buf_8
Xfanout98 _07178_/Y vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__buf_8
Xfanout76 fanout77/X vssd1 vssd1 vccd1 vccd1 fanout76/X sky130_fd_sc_hd__buf_6
XFILLER_0_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _10531_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10461_/Y sky130_fd_sc_hd__xnor2_1
X_12200_ _07075_/Y _12029_/B _12142_/A vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ _13185_/CLK hold212/X vssd1 vssd1 vccd1 vccd1 _13180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _10607_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09718__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ hold237/A _12190_/B _12188_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12131_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12144__A _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12062_ _09952_/X _12061_/Y _12271_/S vssd1 vssd1 vccd1 vccd1 _12062_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07238__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A2 _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _10791_/A _10905_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10722__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10599__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ hold35/X fanout1/X hold37/X vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11915_ _11983_/A _11914_/B _11914_/C vssd1 vssd1 vccd1 vccd1 _11915_/Y sky130_fd_sc_hd__a21oi_1
X_12895_ hold174/X _13084_/B2 _13084_/A2 _13189_/Q vssd1 vssd1 vccd1 vccd1 hold175/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11847_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11777_ _11623_/B _11931_/C hold291/A vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__A _12499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10728_ _10845_/A _10845_/B _07239_/Y _10845_/C _07044_/Y vssd1 vssd1 vccd1 vccd1
+ _10729_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_125_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12950__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ _12507_/B _12330_/B vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06987__A _06987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _10156_/A _07870_/B vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08382__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _06821_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__and2_1
XANTENNA__08382__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06752_ _06512_/Y _06532_/X _06535_/Y _12507_/B vssd1 vssd1 vccd1 vccd1 _06752_/Y
+ sky130_fd_sc_hd__o211ai_4
X_09540_ _10252_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09550_/A sky130_fd_sc_hd__xnor2_2
X_09471_ _09471_/A vssd1 vssd1 vccd1 vccd1 _09471_/Y sky130_fd_sc_hd__inv_2
X_06683_ _06763_/B _06613_/A _12565_/B _06682_/X vssd1 vssd1 vccd1 vccd1 _07278_/A
+ sky130_fd_sc_hd__a31o_4
X_08422_ _08422_/A _08556_/A vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09882__B2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__A1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09302__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _08353_/A _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__or3_1
XANTENNA_fanout142_A _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07611__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ _07304_/A _07304_/B vssd1 vssd1 vccd1 vccd1 _07304_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08284_ _08283_/B _08283_/C _08272_/X vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11441__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07235_ _11184_/A _11184_/B _11271_/A vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_116_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07166_ _12704_/A _07000_/A _12702_/A _10481_/A vssd1 vssd1 vccd1 vccd1 _07167_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07097_ _09634_/A _07186_/A _09309_/S _07184_/B _09495_/A vssd1 vssd1 vccd1 vccd1
+ _07099_/B sky130_fd_sc_hd__o311a_2
XANTENNA__07948__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout200 _12692_/B vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__buf_4
Xfanout211 _07006_/Y vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__buf_8
Xfanout222 _06856_/Y vssd1 vssd1 vccd1 vccd1 _06858_/B sky130_fd_sc_hd__buf_6
Xfanout244 _09342_/X vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__buf_4
Xfanout255 _07842_/A vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__buf_12
Xfanout233 _06749_/X vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__buf_6
Xfanout288 fanout298/X vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__clkbuf_4
Xfanout277 _06665_/A2 vssd1 vssd1 vccd1 vccd1 _12484_/A sky130_fd_sc_hd__buf_4
X_09807_ hold257/A hold296/A hold243/A hold249/A vssd1 vssd1 vccd1 vccd1 _10080_/C
+ sky130_fd_sc_hd__or4_2
Xfanout266 _06537_/Y vssd1 vssd1 vccd1 vccd1 _06613_/A sky130_fd_sc_hd__buf_4
Xfanout299 _12263_/S vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__clkbuf_8
X_07999_ _11656_/A _08159_/A vssd1 vssd1 vccd1 vccd1 _07999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09570__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _09520_/Y _09523_/B _09528_/A vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout55_A _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ curr_PC[3] _09669_/B vssd1 vssd1 vccd1 vccd1 _09957_/C sky130_fd_sc_hd__and2_1
X_11700_ hold269/A _11623_/B _11776_/B _11699_/Y _12313_/A1 vssd1 vssd1 vccd1 vccd1
+ _11700_/X sky130_fd_sc_hd__a311o_1
X_12680_ hold68/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__or2_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _12303_/A _11618_/X _11630_/X _11612_/X vssd1 vssd1 vccd1 vccd1 _11631_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08428__A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11562_ fanout17/X fanout50/X _07988_/B _12728_/A vssd1 vssd1 vccd1 vccd1 _11563_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07100__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10514_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11493_ _11494_/B _11494_/A vssd1 vssd1 vccd1 vccd1 _11585_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13232_ _13260_/CLK _13232_/D vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ _10444_/A _10444_/B vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__nor2_2
X_13163_ _13169_/CLK _13163_/D vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12932__A1 _11184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10375_ _10376_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _06552_/B _12053_/B _06552_/A vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__a21bo_1
X_13094_ _13103_/A hold276/X vssd1 vssd1 vccd1 vccd1 _13250_/D sky130_fd_sc_hd__and2_1
X_12045_ _12107_/B _12045_/B vssd1 vssd1 vccd1 vccd1 _12047_/A sky130_fd_sc_hd__or2_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08116__B2 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ hold113/A _12665_/A _12955_/B1 hold92/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold93/A sky130_fd_sc_hd__o221a_1
XFILLER_0_62_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11120__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _13062_/A hold211/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__and2_1
XANTENNA__07431__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _11828_/A _11828_/B _11828_/C vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07150__B _07152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A2 _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07020_ _07021_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07216_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07577__S _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09358__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__xnor2_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _07925_/A _07925_/B vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__nor2_1
X_07853_ _07771_/A _07771_/B _07771_/C vssd1 vssd1 vccd1 vccd1 _07854_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07606__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _07103_/A _07064_/A vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07784_ _07884_/A _07884_/B _07783_/A vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08107__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06735_ reg2_val[4] _06748_/B vssd1 vssd1 vccd1 vccd1 _06735_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ _09523_/A _09523_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08658__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06666_ reg1_val[15] _06936_/A vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__nand2_1
X_09454_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08405_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__and2b_1
X_09385_ _09243_/A _09243_/B _09241_/Y vssd1 vssd1 vccd1 vccd1 _09387_/B sky130_fd_sc_hd__a21oi_1
X_06597_ instruction[33] _06637_/B vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__and2_4
XFILLER_0_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ _08335_/A _08335_/B _08408_/A vssd1 vssd1 vccd1 vccd1 _08336_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08267_ _08267_/A _08267_/B vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_117_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _06977_/A _12710_/A _12712_/A _06985_/A vssd1 vssd1 vccd1 vccd1 _07219_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08172__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12914__A1 _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _07149_/A _07149_/B _07152_/B vssd1 vssd1 vccd1 vccd1 _07156_/A sky130_fd_sc_hd__and3_2
XANTENNA__11717__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10160_ _10158_/X _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08594__B2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _10091_/A _10091_/B _10091_/C _10091_/D vssd1 vssd1 vccd1 vccd1 _10091_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__12141__B fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07235__B _11184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _13004_/B _13005_/A _12771_/X vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09846__A1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _10993_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__xor2_1
X_12732_ _13105_/A hold7/X vssd1 vssd1 vccd1 vccd1 _12832_/B sky130_fd_sc_hd__or2_1
XFILLER_0_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09846__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07251__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ rst _12663_/B _12663_/C vssd1 vssd1 vccd1 vccd1 _13125_/D sky130_fd_sc_hd__nor3_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11614_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11615_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12599_/A _12594_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11545_ curr_PC[19] _11633_/C _11713_/A vssd1 vssd1 vccd1 vccd1 _11545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ _12089_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13215_ _13217_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08082__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10427_ _10298_/A _10298_/B _10296_/Y vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10117__A _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13146_ _13188_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09782__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _10301_/A _10301_/B _10299_/Y vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13077_ _13077_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13077_/Y sky130_fd_sc_hd__xnor2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12133__A2 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _12148_/A fanout8/X fanout5/X _12094_/A vssd1 vssd1 vccd1 vccd1 _12030_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08888__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06520_ curr_PC[0] vssd1 vssd1 vccd1 vccd1 _06520_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07312__A2 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09170_ instruction[5] _06813_/X _09151_/A _09134_/X _09169_/X vssd1 vssd1 vccd1
+ vccd1 _09170_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07076__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08121_/X sky130_fd_sc_hd__and2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _08535_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08238_/B sky130_fd_sc_hd__xnor2_1
X_07003_ _12704_/A _10481_/A _07000_/A _12706_/A vssd1 vssd1 vccd1 vccd1 _07004_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08954_ fanout92/X fanout38/X _10647_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _08955_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07905_ _06938_/A _06938_/B _08740_/A2 vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08879__A2 _08985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ _09568_/A _12141_/A _07391_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _08886_/B
+ sky130_fd_sc_hd__o22a_1
X_07836_ _10957_/A _06977_/A _06985_/A fanout80/X vssd1 vssd1 vccd1 vccd1 _07837_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07767_ _07768_/B _07768_/C _07768_/A vssd1 vssd1 vccd1 vccd1 _07771_/A sky130_fd_sc_hd__a21o_1
X_06718_ reg1_val[7] _07123_/A vssd1 vssd1 vccd1 vccd1 _06719_/B sky130_fd_sc_hd__nand2_1
X_09506_ _09474_/X _09488_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07698_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06649_ reg1_val[17] _07165_/A vssd1 vssd1 vccd1 vccd1 _06787_/A sky130_fd_sc_hd__nand2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09439_/B sky130_fd_sc_hd__xnor2_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09578_/B _09368_/B vssd1 vssd1 vccd1 vccd1 _09370_/C sky130_fd_sc_hd__or2_1
X_09299_ _09297_/X _09298_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09299_/X sky130_fd_sc_hd__mux2_1
X_08319_ _08319_/A _08319_/B vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout18_A _07070_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_60 pred_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ _11329_/A _11329_/B _11418_/B vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _11233_/Y _11234_/X _11236_/Y _09145_/Y _11260_/X vssd1 vssd1 vccd1 vccd1
+ _11261_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08016__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13000_ _13000_/A _13000_/B vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__xnor2_1
X_10212_ hold300/A _09808_/B _10469_/C _09810_/A vssd1 vssd1 vccd1 vccd1 _10212_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08630__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _12089_/A _11192_/B vssd1 vssd1 vccd1 vccd1 _11196_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10144_/C sky130_fd_sc_hd__xnor2_1
X_10074_ _10073_/X _09290_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _10074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__and2_1
X_12715_ hold17/X _12720_/B _12714_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__o211a_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ _12578_/A _12578_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _10828_/A _11527_/Y _12125_/S vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08007__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ _11460_/B _11459_/B vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10365__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ _13208_/CLK _13129_/D vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07230__A1 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10365__B2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06995__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08670_ _08755_/A _08670_/A2 _08699_/A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08671_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07621_ _08903_/B _07621_/B vssd1 vssd1 vccd1 vccd1 _07623_/B sky130_fd_sc_hd__nor2_2
X_07552_ _07473_/A _07473_/B _07474_/Y vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07483_ _07484_/A _07484_/B vssd1 vssd1 vccd1 vccd1 _07489_/B sky130_fd_sc_hd__and2_1
XFILLER_0_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09222_ _09422_/A fanout9/X fanout4/X _09222_/B2 vssd1 vssd1 vccd1 vccd1 _09223_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ fanout79/X _08735_/A2 _08735_/B1 _08430_/B vssd1 vssd1 vccd1 vccd1 _08105_/B
+ sky130_fd_sc_hd__o22a_1
X_09084_ _10920_/A reg1_val[18] _09092_/S vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ _08853_/B _08853_/A vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10980__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10356__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _09986_/A _09986_/B _09986_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__nand3_1
X_08937_ _07599_/Y _07609_/B _07607_/Y vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__a21o_1
X_08868_ _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08870_/B sky130_fd_sc_hd__xnor2_1
X_07819_ _07819_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__xnor2_2
X_08799_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07513__B _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _12303_/A _10816_/X _10829_/X _10807_/Y vssd1 vssd1 vccd1 vccd1 _10830_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__A1 _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__B2 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08485__B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _10761_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _10692_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10692_/Y sky130_fd_sc_hd__nor2_1
X_12500_ _12504_/A _12500_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__nor2_8
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ reg1_val[17] curr_PC[17] _12444_/S vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12362_ _12368_/B _12362_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
XANTENNA__10595__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12293_ _12257_/Y _12258_/X _12290_/Y _12292_/X _12112_/A vssd1 vssd1 vccd1 vccd1
+ _12293_/X sky130_fd_sc_hd__a221o_1
X_11313_ _11314_/B _11314_/A vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__nand2b_1
X_11244_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11245_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11175_ _11654_/A _11175_/B vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__xnor2_1
X_10126_ _10126_/A _10126_/B _10126_/C vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__nand3_1
X_10057_ _09621_/A _09019_/A _09019_/B _09145_/Y _10056_/Y vssd1 vssd1 vccd1 vccd1
+ _10091_/B sky130_fd_sc_hd__o311a_1
XANTENNA__07704__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07279__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07279__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10959_ _11102_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10961_/B sky130_fd_sc_hd__and2_1
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10348__A2_N _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ _12629_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10586__A1 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ fanout77/X fanout42/X _07239_/A fanout74/X vssd1 vssd1 vccd1 vccd1 _09841_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06983_ _07012_/B _06983_/B vssd1 vssd1 vccd1 vccd1 _06983_/Y sky130_fd_sc_hd__xnor2_4
X_09771_ _09614_/B _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__and3b_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10353__A4 _10352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08726_/C sky130_fd_sc_hd__xnor2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07614__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__and2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10510__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 fanout4/A sky130_fd_sc_hd__or2_2
X_08584_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__and2_1
X_07535_ _07731_/A _07731_/B _07534_/A vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10975__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09205_ _10009_/A fanout63/X fanout60/X _09725_/B2 vssd1 vssd1 vccd1 vccd1 _09206_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ _07397_/A _07397_/B vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07690__A1 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__B2 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12015__B2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _12053_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07442__A1 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ reg1_val[1] reg1_val[30] _09092_/S vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08018_ _08166_/A _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout85_A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__nor2_2
X_12980_ _13111_/A hold258/X vssd1 vssd1 vccd1 vccd1 _13226_/D sky130_fd_sc_hd__and2_1
X_11931_ hold292/A hold291/A _11931_/C vssd1 vssd1 vccd1 vccd1 _11998_/B sky130_fd_sc_hd__or3_1
X_11862_ _12303_/A _11850_/X _11861_/X _11844_/X vssd1 vssd1 vccd1 vccd1 _11862_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _10695_/X _10697_/Y _10811_/X _10812_/Y vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11793_ _12148_/A fanout15/X _07112_/Y fanout17/X vssd1 vssd1 vccd1 vccd1 _11794_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ _10744_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__and2_1
X_12414_ _12571_/B _12414_/B vssd1 vssd1 vccd1 vccd1 _12415_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10017__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12345_ _12354_/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12347_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12309__A2 _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09186__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12276_ _12190_/B _12275_/X _13189_/Q vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09617__C _09617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11517__B1 _09146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ _11329_/A _11227_/B vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__and2_1
XANTENNA__10125__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _11158_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__nor2_1
X_11089_ _11087_/X _11089_/B vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08697__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07320_ _12085_/A _07320_/B vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09661__A2 _09637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _09423_/A _07251_/B vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__B1 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07182_ _11794_/A _07187_/B _11883_/A vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09413__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07188__B1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _09762_/A _09762_/B _09763_/Y vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__06935__B1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__nor2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09596_/A _09596_/B _09595_/A vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09543__B _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ instruction[40] _06532_/X _06895_/X _06896_/Y vssd1 vssd1 vccd1 vccd1 _06897_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _09685_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__or2_2
X_08705_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08706_/C sky130_fd_sc_hd__nand2_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08741_/A _08636_/B vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06702__A3 _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout22 _12223_/A vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__buf_2
XFILLER_0_49_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout11 _12141_/A vssd1 vssd1 vccd1 vccd1 fanout11/X sky130_fd_sc_hd__clkbuf_8
X_08567_ _08607_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _08603_/B sky130_fd_sc_hd__xnor2_1
X_07518_ _07154_/X _07185_/Y _07271_/X _07799_/B vssd1 vssd1 vccd1 vccd1 _07519_/B
+ sky130_fd_sc_hd__a22o_1
Xfanout33 _12248_/B vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__buf_8
Xfanout55 _12718_/A vssd1 vssd1 vccd1 vccd1 fanout55/X sky130_fd_sc_hd__buf_4
Xfanout44 _07391_/B vssd1 vssd1 vccd1 vccd1 fanout44/X sky130_fd_sc_hd__buf_6
XFILLER_0_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08498_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__xor2_1
X_07449_ _07449_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11995__B1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout66 _07017_/Y vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__clkbuf_8
Xfanout77 _06983_/Y vssd1 vssd1 vccd1 vccd1 fanout77/X sky130_fd_sc_hd__buf_8
Xfanout88 _07304_/Y vssd1 vssd1 vccd1 vccd1 _12690_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout99 _12702_/A vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__buf_6
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _10458_/Y _10460_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09115_/X _09118_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10391_ _10481_/A fanout9/X fanout3/X _07000_/A vssd1 vssd1 vccd1 vccd1 _10392_/B
+ sky130_fd_sc_hd__o22a_1
X_12130_ _12190_/B _12188_/B hold237/A vssd1 vssd1 vccd1 vccd1 _12130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07519__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _12061_/A _12061_/B vssd1 vssd1 vccd1 vccd1 _12061_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07238__B _11184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__A3 _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__A1 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _11012_/A _11012_/B vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10722__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__B2 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ hold37/X hold35/X fanout1/X vssd1 vssd1 vccd1 vccd1 _12963_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11914_ _11983_/A _11914_/B _11914_/C vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _13085_/A hold234/X vssd1 vssd1 vccd1 vccd1 _13188_/D sky130_fd_sc_hd__and2_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__or2_1
XFILLER_0_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ hold269/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11931_/C sky130_fd_sc_hd__or2_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10727_/A _10727_/B vssd1 vssd1 vccd1 vccd1 _10738_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _10658_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10660_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _09808_/B _10708_/B hold277/A vssd1 vssd1 vccd1 vccd1 _10589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12328_ reg1_val[2] curr_PC[2] _12444_/S vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10410__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _12112_/A _12258_/X _12257_/Y vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08382__A2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06819_/A _06819_/B _12221_/A vssd1 vssd1 vccd1 vccd1 _06821_/B sky130_fd_sc_hd__a21o_1
X_06751_ reg1_val[2] _09634_/A vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09470_ _10201_/S _09317_/X _09164_/B vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__o21ai_1
X_06682_ reg2_val[12] _06748_/B vssd1 vssd1 vccd1 vccd1 _06682_/X sky130_fd_sc_hd__and2_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08421_ _08421_/A _08424_/A _08421_/C vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ _08352_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08353_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07303_ _07303_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07304_/B sky130_fd_sc_hd__and2_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08283_ _08272_/X _08283_/B _08283_/C vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _11271_/A _11184_/B _11184_/A vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10464__S _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ _07165_/A _07165_/B vssd1 vssd1 vccd1 vccd1 _07165_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout302_A _06511_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _07186_/A _09309_/S _09495_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07271_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07948__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 _12664_/Y vssd1 vssd1 vccd1 vccd1 _12692_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout212 _06904_/X vssd1 vssd1 vccd1 vccd1 _12280_/A sky130_fd_sc_hd__clkbuf_8
Xfanout223 _12668_/A vssd1 vssd1 vccd1 vccd1 _08755_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__09554__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 _09342_/X vssd1 vssd1 vccd1 vccd1 _12000_/A2 sky130_fd_sc_hd__buf_2
Xfanout234 _11134_/S vssd1 vssd1 vccd1 vccd1 _11033_/A sky130_fd_sc_hd__buf_4
Xfanout289 fanout298/X vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__buf_2
Xfanout267 _12662_/A vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__buf_4
X_09806_ _10208_/B _10077_/C hold239/A vssd1 vssd1 vccd1 vccd1 _09806_/Y sky130_fd_sc_hd__a21oi_1
Xfanout278 _06665_/A2 vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__buf_6
X_07998_ _08165_/A _08165_/B _07993_/Y vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09570__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A1 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _08916_/A _06949_/B vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07581__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__A _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _09737_/A _09737_/B vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10468__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ curr_PC[3] _09669_/B vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__or2_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09599_ _09372_/A _09372_/B _09371_/A vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__o21ai_2
X_08619_ _08623_/A _08623_/B vssd1 vssd1 vccd1 vccd1 _08624_/A sky130_fd_sc_hd__nor2_1
X_11630_ _11448_/A _11620_/X _11621_/Y _11629_/X vssd1 vssd1 vccd1 vccd1 _11630_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07097__C1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11561_ _11662_/B _11561_/B vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10514_/A sky130_fd_sc_hd__and2_1
XANTENNA__10640__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ _11585_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11494_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13231_ _13234_/CLK _13231_/D vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
X_10443_ _10443_/A _10443_/B _10443_/C vssd1 vssd1 vccd1 vccd1 _10444_/B sky130_fd_sc_hd__and3_1
X_13162_ _13169_/CLK hold196/X vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10374_ _10374_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__xnor2_2
X_12113_ _12113_/A _12113_/B _12113_/C vssd1 vssd1 vccd1 vccd1 _12113_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ hold275/X _06858_/B _13092_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold276/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09464__A _09464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12044_ _11976_/B _11975_/Y _12160_/A _12042_/X vssd1 vssd1 vccd1 vccd1 _12045_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08116__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10122__B _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ _07916_/A _12962_/B2 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__o21a_1
XANTENNA__08808__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ hold210/X _12885_/A2 _12885_/B1 _13180_/Q vssd1 vssd1 vccd1 vccd1 hold211/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11828_/A _11828_/B _11828_/C vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__nand3_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _11869_/A _11759_/B vssd1 vssd1 vccd1 vccd1 _11834_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__11423__A2 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10226__A3 _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08543__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08971_/B sky130_fd_sc_hd__xor2_4
XANTENNA__06998__A _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__B _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ _08801_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07925_/B sky130_fd_sc_hd__xnor2_1
X_07852_ _07714_/X _07829_/Y _07850_/B _07960_/A vssd1 vssd1 vccd1 vccd1 _07879_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ reg1_val[27] _07044_/A vssd1 vssd1 vccd1 vccd1 _06803_/Y sky130_fd_sc_hd__nand2_1
X_07783_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07884_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08107__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _11726_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09523_/B sky130_fd_sc_hd__xor2_1
X_06734_ _06734_/A _06734_/B vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09313__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06665_ _06763_/B _06665_/A2 _06646_/A _06663_/X vssd1 vssd1 vccd1 vccd1 _06936_/A
+ sky130_fd_sc_hd__a31oi_4
X_09453_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout252_A _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08454_/B sky130_fd_sc_hd__xnor2_1
X_09384_ _09534_/B _09384_/B vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10870__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06596_ _06596_/A _06596_/B vssd1 vssd1 vccd1 vccd1 _06839_/A sky130_fd_sc_hd__nor2_1
X_08335_ _08335_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07217_ _07565_/B _07217_/B vssd1 vssd1 vccd1 vccd1 _07276_/A sky130_fd_sc_hd__or2_1
X_08197_ _08144_/A _08144_/B _08142_/Y vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__12914__A2 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07069__A _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ reg1_val[24] _07148_/B vssd1 vssd1 vccd1 vccd1 _07152_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08594__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _07079_/A _07079_/B _07079_/C vssd1 vssd1 vccd1 vccd1 _07081_/A sky130_fd_sc_hd__and3_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _12303_/A _10076_/X _10089_/X vssd1 vssd1 vccd1 vccd1 _10091_/D sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07554__B1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _12999_/B _13000_/A _12773_/X vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07306__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ _10992_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10993_/B sky130_fd_sc_hd__nand2_1
X_12731_ _11385_/B _12731_/A2 hold65/X _13111_/A vssd1 vssd1 vccd1 vccd1 _13158_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A hold163/X vssd1 vssd1 vccd1 vccd1 _12663_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11613_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__or2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12593_ _12615_/B _07087_/B _12599_/B vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ curr_PC[19] _11633_/C vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _11739_/A fanout11/X fanout44/X fanout64/X vssd1 vssd1 vccd1 vccd1 _11476_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13217_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ _10274_/B _10290_/B _10272_/Y vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10117__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _13188_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07793__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ curr_PC[9] _10597_/C vssd1 vssd1 vccd1 vccd1 _10357_/X sky130_fd_sc_hd__xor2_1
X_13076_ _13080_/A _13076_/B vssd1 vssd1 vccd1 vccd1 _13246_/D sky130_fd_sc_hd__and2_1
XANTENNA__07707__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12027_ _12102_/B _12027_/B vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__and2b_1
X_12929_ hold141/A _12665_/A _12955_/B1 hold85/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold86/A sky130_fd_sc_hd__o221a_1
XFILLER_0_88_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10852__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07076__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__A1 _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__B1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__B _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08051_ _08565_/B _08715_/A2 _08735_/B1 fanout83/X vssd1 vssd1 vccd1 vccd1 _08052_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07002_ _07002_/A _07002_/B vssd1 vssd1 vccd1 vccd1 _07002_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09222__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09308__S _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _08953_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08956_/A sky130_fd_sc_hd__nor2_1
X_07904_ _08607_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ _07624_/A _07624_/B _07622_/Y vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__o21ai_4
X_07835_ _07839_/A _07839_/B vssd1 vssd1 vccd1 vccd1 _07835_/X sky130_fd_sc_hd__or2_1
X_07766_ _07768_/B _07768_/C _07768_/A vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08448__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06717_ _06717_/A vssd1 vssd1 vccd1 vccd1 _06719_/A sky130_fd_sc_hd__inv_2
X_09505_ reg1_val[2] _09634_/A _12309_/B1 vssd1 vssd1 vccd1 vccd1 _09505_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07697_ _07810_/A _07810_/B _07696_/A vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07071__B _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06648_ _06978_/A vssd1 vssd1 vccd1 vccd1 _07165_/A sky130_fd_sc_hd__inv_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ _06579_/A _11935_/A vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__and2_1
X_09367_ _09366_/B _09367_/B vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__and2b_1
X_09298_ _09074_/X _09076_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09298_/X sky130_fd_sc_hd__mux2_1
XANTENNA_50 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08318_ _08318_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08319_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_72 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 reg1_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08249_ _08249_/A _08249_/B vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08016__A1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12899__B2 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _11240_/Y _11241_/X _11248_/X _11259_/X vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08016__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10211_ _09808_/B _10469_/C hold300/A vssd1 vssd1 vccd1 vccd1 _10211_/Y sky130_fd_sc_hd__a21oi_1
X_11191_ _11462_/A fanout11/X fanout44/X fanout76/X vssd1 vssd1 vccd1 vccd1 _11192_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07527__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _09482_/X _09485_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11874__A2 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12714_ _12714_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12714_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11626__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10975_ _12086_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12645_ reg1_val[29] _12656_/A vssd1 vssd1 vccd1 vccd1 _12646_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12576_ reg1_val[15] _12576_/B vssd1 vssd1 vccd1 vccd1 _12578_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11527_ _11527_/A _11527_/B vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09917__A _10321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08007__B2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08007__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ _11458_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__A _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11390_/A _11390_/B _11390_/C vssd1 vssd1 vccd1 vccd1 _11391_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _10257_/A _10257_/B _10255_/X vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13128_ _13208_/CLK _13128_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07230__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__B2 _12728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13059_/A _13059_/B vssd1 vssd1 vccd1 vccd1 _13059_/Y sky130_fd_sc_hd__xnor2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07172__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07551_ _07661_/A _07661_/B _07661_/C vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12248__A_N _12728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07482_ _07875_/A _07482_/B vssd1 vssd1 vccd1 vccd1 _07484_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07297__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08494__A1 _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _09221_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08103_ _11470_/A _08101_/B _08150_/A vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_114_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _09081_/X _09082_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09083_/X sky130_fd_sc_hd__mux2_1
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ _09986_/A _09986_/B _09986_/C vssd1 vssd1 vccd1 vccd1 _10168_/A sky130_fd_sc_hd__a21o_1
X_08936_ _08936_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__nor2_1
X_08867_ _08864_/A _08864_/B _08868_/B vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09562__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12700__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07818_ _07818_/A _07818_/B vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06709__A_N _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ _09313_/S _08798_/B vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__or2_1
X_07749_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08906__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout30_A _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _11184_/A _10760_/B vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08485__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__B2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10691_ _11238_/A _10690_/X _10689_/X vssd1 vssd1 vccd1 vccd1 _10692_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _09862_/B _09419_/B vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__xnor2_2
X_12430_ _12439_/A _12430_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
XANTENNA__06859__A_N _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _12361_/A _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11241__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _12290_/A _12290_/B _12290_/C vssd1 vssd1 vccd1 vccd1 _12292_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11312_/A _11312_/B vssd1 vssd1 vccd1 vccd1 _11314_/B sky130_fd_sc_hd__xnor2_1
X_11243_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11243_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10347__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07257__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11174_ fanout60/X fanout41/X _08135_/B _12148_/A vssd1 vssd1 vccd1 vccd1 _11175_/B
+ sky130_fd_sc_hd__o22a_1
X_10125_ _10607_/A _10125_/B _10125_/C vssd1 vssd1 vccd1 vccd1 _10126_/C sky130_fd_sc_hd__nand3_1
X_10056_ _09621_/A _09019_/B _09019_/A vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08173__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__B1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10411__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__A2 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10958_ _10957_/A _11296_/A _10957_/C vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10283__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ reg1_val[26] _12656_/A vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__nand2_1
X_10889_ _10738_/A _10738_/B _10748_/X vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11783__A1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ reg1_val[12] _12559_/B vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold106 hold108/X vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07167__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _06982_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__xnor2_4
X_09770_ _10049_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__nor2_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__nand2b_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08655_/A sky130_fd_sc_hd__xnor2_1
X_07603_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__nor2_4
XANTENNA__10321__A _10321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08583_ _08564_/Y _08569_/B _08582_/X vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__o21a_1
X_07534_ _07534_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09321__S _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09204_ _10607_/A _09204_/B vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07396_ _07396_/A _07396_/B vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07690__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09135_ _11238_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09135_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07442__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _12499_/A reg1_val[31] _09092_/S vssd1 vssd1 vccd1 vccd1 _09066_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ _10853_/A _08017_/B vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__nor2_1
X_08919_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _09194_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout78_A fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _11930_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _11930_/X sky130_fd_sc_hd__or2_1
X_09899_ _09737_/A _09737_/B _09735_/Y vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _11852_/Y _11853_/X _11857_/X _11860_/X vssd1 vssd1 vccd1 vccd1 _11861_/X
+ sky130_fd_sc_hd__o211a_1
X_10812_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10812_/Y sky130_fd_sc_hd__nand2_1
X_11792_ _11743_/A _11743_/B _11744_/Y vssd1 vssd1 vccd1 vccd1 _11827_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10743_ _10744_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__and2_1
XANTENNA__08636__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12006__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _10674_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10676_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10017__A1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _12571_/B _12414_/B vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10017__B2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__B1 _12248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ _12517_/B _12344_/B vssd1 vssd1 vccd1 vccd1 _12345_/B sky130_fd_sc_hd__or2_1
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12275_ hold174/A hold233/A _12275_/C vssd1 vssd1 vccd1 vccd1 _12275_/X sky130_fd_sc_hd__or3_1
XFILLER_0_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _11226_/A _11226_/B _11226_/C vssd1 vssd1 vccd1 vccd1 _11227_/B sky130_fd_sc_hd__nand3_1
X_11157_ _11157_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11163_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ _10108_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__xnor2_4
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__or2_1
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08697__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08697__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__A1 _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11185__A2_N fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ _09422_/A _12094_/A _12148_/A _09222_/B2 vssd1 vssd1 vccd1 vccd1 _07251_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07181_ _11794_/A _07187_/B _11883_/A vssd1 vssd1 vccd1 vccd1 _07183_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09377__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10316__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A1 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__C1 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__B2 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__B1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _09767_/A _09767_/B _09765_/X vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__a21o_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09753_ _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__xor2_1
X_06965_ _10156_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__xor2_1
X_08704_ _08704_/A _08704_/B vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__xor2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__C _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ instruction[6] is_load vssd1 vssd1 vccd1 vccd1 _06896_/Y sky130_fd_sc_hd__nor2_1
X_09684_ _09683_/B _09684_/B vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08635_ _08740_/A2 _08737_/A2 _08733_/B1 _08755_/B vssd1 vssd1 vccd1 vccd1 _08636_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08606_/A2 _08782_/B2 _08813_/B1 _08642_/B vssd1 vssd1 vccd1 vccd1 _08567_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ _07533_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__nand2_1
Xfanout12 _07183_/X vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__buf_6
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11444__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout23 _11620_/B vssd1 vssd1 vccd1 vccd1 _11781_/B sky130_fd_sc_hd__buf_4
Xfanout56 _07059_/X vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__buf_4
XFILLER_0_91_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout45 _07391_/B vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__buf_4
XFILLER_0_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout34 _08233_/B vssd1 vssd1 vccd1 vccd1 fanout34/X sky130_fd_sc_hd__clkbuf_8
X_08497_ _08497_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07448_ _07444_/A _07444_/B _07507_/A vssd1 vssd1 vccd1 vccd1 _07468_/B sky130_fd_sc_hd__a21o_1
Xfanout89 _12688_/A vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__buf_8
Xfanout67 _12712_/A vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__clkbuf_8
Xfanout78 fanout79/X vssd1 vssd1 vccd1 vccd1 fanout78/X sky130_fd_sc_hd__clkbuf_8
X_07379_ _07405_/A _07405_/B _07376_/Y vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12706__A _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _09116_/X _09117_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ _10285_/A _10285_/B _10282_/A vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ _09049_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _11914_/C sky130_fd_sc_hd__and2_1
X_12060_ _12058_/Y _12060_/B vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08915__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _11012_/A _11012_/B vssd1 vssd1 vccd1 vccd1 _11159_/A sky130_fd_sc_hd__and2_1
XANTENNA__10722__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ hold37/X _13112_/B _12248_/B _12962_/B2 _12961_/Y vssd1 vssd1 vccd1 vccd1
+ hold38/A sky130_fd_sc_hd__o221a_1
XANTENNA__11057__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ hold233/X _13084_/B2 _13084_/A2 hold174/X vssd1 vssd1 vccd1 vccd1 hold234/A
+ sky130_fd_sc_hd__a22o_1
X_11913_ _11913_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _11913_/Y sky130_fd_sc_hd__nand2_1
X_11844_ _06837_/A _11842_/X _11843_/Y vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__a21o_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11696_/A _11773_/Y _11774_/Y _09156_/B vssd1 vssd1 vccd1 vccd1 _11786_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08300__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10726_ _10727_/A _10727_/B vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__or2_1
XFILLER_0_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ _10776_/B _10657_/B vssd1 vssd1 vccd1 vccd1 _10658_/B sky130_fd_sc_hd__or2_1
X_10588_ hold255/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12327_ _12333_/B _12327_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10410__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10410__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12258_ _12258_/A _12258_/B _12258_/C _12258_/D vssd1 vssd1 vccd1 vccd1 _12258_/X
+ sky130_fd_sc_hd__and4_1
X_11209_ _11092_/A _11092_/B _11095_/A vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__o21bai_1
X_12189_ _12190_/B _12275_/C hold233/A vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12351__A _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _09634_/A reg1_val[2] vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__and2b_1
X_06681_ _10933_/A _06681_/B vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08420_ _08421_/A _08424_/A _08421_/C vssd1 vssd1 vccd1 vccd1 _08422_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__A _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__B1 _10321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ _08272_/X _08281_/Y _08335_/A vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ _08272_/A _08272_/B _08272_/C vssd1 vssd1 vccd1 vccd1 _08283_/C sky130_fd_sc_hd__a21o_1
X_07302_ _11183_/A _11385_/A _07300_/X vssd1 vssd1 vccd1 vccd1 _07302_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _11184_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout128_A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ _06945_/A _06979_/A _06943_/B _07289_/B vssd1 vssd1 vccd1 vccd1 _07165_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12245__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07095_ reg1_val[27] _07095_/B vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout202 _12277_/B1 vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__buf_4
Xfanout213 _06904_/X vssd1 vssd1 vccd1 vccd1 _12238_/C1 sky130_fd_sc_hd__clkbuf_4
Xfanout246 _12304_/B1 vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__buf_4
Xfanout224 _09313_/S vssd1 vssd1 vccd1 vccd1 _09319_/S sky130_fd_sc_hd__clkbuf_8
Xfanout235 _10924_/S vssd1 vssd1 vccd1 vccd1 _11134_/S sky130_fd_sc_hd__buf_4
Xfanout268 _06509_/Y vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__buf_4
X_09805_ hold239/A _10208_/B _10077_/C vssd1 vssd1 vccd1 vccd1 _09805_/X sky130_fd_sc_hd__and3_1
XANTENNA__07581__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _11713_/A vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__buf_8
Xfanout279 _06665_/A2 vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__buf_6
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09570__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ fanout82/X fanout80/X _06940_/A _10099_/A1 vssd1 vssd1 vccd1 vccd1 _06949_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07581__B2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__B _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ _09736_/A _09736_/B vssd1 vssd1 vccd1 vccd1 _09737_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09858__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _10924_/S _12280_/A _09620_/Y _09666_/X vssd1 vssd1 vccd1 vccd1 _09667_/X
+ sky130_fd_sc_hd__a211o_2
X_06879_ instruction[25] _06887_/B vssd1 vssd1 vccd1 vccd1 _06879_/X sky130_fd_sc_hd__or2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08530__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _08625_/A _08625_/B _08617_/A vssd1 vssd1 vccd1 vccd1 _08623_/B sky130_fd_sc_hd__a21oi_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09448_/A _09448_/B _09446_/Y vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08549_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _08560_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07097__B1 _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _11559_/B _11560_/B vssd1 vssd1 vccd1 vccd1 _11561_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout7_A fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ _11068_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10513_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10640__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13031__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13230_/CLK _13230_/D vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _11491_/A _11491_/B _11491_/C vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10640__B2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _10443_/A _10443_/B _10443_/C vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__a21o_1
X_13161_ _13169_/CLK _13161_/D vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_1
X_10373_ _10371_/X _10373_/B vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__nand2b_1
X_13092_ hold265/X _13091_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_1
X_12112_ _12112_/A _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12113_/C sky130_fd_sc_hd__or3_1
X_12043_ _11976_/A _11976_/B _11972_/A _11974_/B _12160_/A vssd1 vssd1 vccd1 vccd1
+ _12107_/B sky130_fd_sc_hd__a311oi_2
XANTENNA__11353__C1 _11350_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10122__C _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12945_ hold122/A _12662_/A _12955_/B1 hold113/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o221a_1
X_12876_ _13062_/A hold169/X vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11827_ _11827_/A _11827_/B vssd1 vssd1 vccd1 vccd1 _11828_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12081__B1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11758_ _11599_/X _11757_/Y _11678_/B vssd1 vssd1 vccd1 vccd1 _11759_/B sky130_fd_sc_hd__a21oi_2
X_10709_ _09808_/B _10820_/B hold261/A vssd1 vssd1 vccd1 vccd1 _10709_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08824__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11689_ _11689_/A _11689_/B vssd1 vssd1 vccd1 vccd1 _11689_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10934__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ _11295_/B2 _08756_/B2 _11297_/A _08782_/A2 vssd1 vssd1 vccd1 vccd1 _07921_/B
+ sky130_fd_sc_hd__o22a_1
X_07851_ _07959_/A _07959_/B _07959_/C vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__o21ai_1
X_06802_ reg1_val[28] _07067_/A vssd1 vssd1 vccd1 vccd1 _06819_/A sky130_fd_sc_hd__nand2_1
X_07782_ _07782_/A _07782_/B _07854_/A vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__nor3_1
X_06733_ reg1_val[5] _06928_/C vssd1 vssd1 vccd1 vccd1 _06734_/B sky130_fd_sc_hd__and2_1
XFILLER_0_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ fanout13/X _07763_/B _12690_/A _07156_/X vssd1 vssd1 vccd1 vccd1 _09522_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06664_ _06763_/B _06665_/A2 _06646_/A _06663_/X vssd1 vssd1 vccd1 vccd1 _06941_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06519__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__xnor2_4
X_06595_ _12297_/A _12264_/A _12221_/A _12175_/A vssd1 vssd1 vccd1 vccd1 _06596_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08403_ _08401_/A _08401_/B _08402_/X vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__o21ba_1
X_09383_ _09383_/A _09383_/B vssd1 vssd1 vccd1 vccd1 _09384_/B sky130_fd_sc_hd__or2_1
XANTENNA__10870__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__B2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_A _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _08280_/A _08280_/B _08280_/C vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08734__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ _08266_/B _08266_/A vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07216_ _07216_/A _07216_/B _07216_/C vssd1 vssd1 vccd1 vccd1 _07217_/B sky130_fd_sc_hd__nor3_1
X_08196_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07069__B _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ _07147_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07147_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12127__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _08276_/A _07078_/B _07078_/C vssd1 vssd1 vccd1 vccd1 _07079_/C sky130_fd_sc_hd__or3_1
XFILLER_0_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07003__B1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__B1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__C1 _12502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout60_A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__B2 _07305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__A1 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _09720_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__nand2_1
X_10991_ _10991_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13241_/CLK sky130_fd_sc_hd__clkbuf_8
X_12730_ hold64/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__or2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ hold23/X hold162/X vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__nand2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11612_ _06837_/D _11610_/X _11611_/Y vssd1 vssd1 vccd1 vccd1 _11612_/X sky130_fd_sc_hd__a21o_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12592_ _12592_/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__or2_1
XFILLER_0_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11543_ _06980_/A _12280_/A _06907_/A _11542_/X vssd1 vssd1 vccd1 vccd1 _11543_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _11474_/A _11474_/B vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11070__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ _13217_/CLK _13213_/D vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _10425_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__xnor2_1
X_13144_ _13188_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10377__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__A1 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10356_ _11153_/A _10597_/C _10355_/Y _10353_/X vssd1 vssd1 vccd1 vccd1 dest_val[8]
+ sky130_fd_sc_hd__o31ai_4
X_13075_ hold292/X _13084_/A2 _13074_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 _13076_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12669__A2 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__B2 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__nand2_1
X_12026_ _12026_/A _12026_/B vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__or2_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ _06961_/B _12692_/B hold142/X vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10852__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ _13170_/Q _12885_/A2 _12885_/B1 hold207/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__A2 _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10604__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _08050_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ _06980_/B _07065_/A _07058_/B1 vssd1 vssd1 vccd1 vccd1 _07002_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09222__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _08952_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__nor2_1
X_08883_ _07653_/A _07653_/B _07654_/Y vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__a21bo_2
X_07903_ _08642_/B fanout93/X _12690_/A _08606_/A2 vssd1 vssd1 vccd1 vccd1 _07904_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout195_A _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _10126_/A _07834_/B vssd1 vssd1 vccd1 vccd1 _07839_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11332__A2 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08733__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _07764_/B _07764_/C _10853_/A vssd1 vssd1 vccd1 vccd1 _07768_/C sky130_fd_sc_hd__a21o_1
X_06716_ reg1_val[7] _07123_/A vssd1 vssd1 vccd1 vccd1 _06717_/A sky130_fd_sc_hd__nor2_1
X_09504_ _09634_/A _12238_/C1 _09150_/Y _09503_/Y vssd1 vssd1 vccd1 vccd1 _09504_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07696_ _07696_/A _07696_/B vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06647_ reg2_val[17] _06700_/B _06657_/B1 _06646_/X vssd1 vssd1 vccd1 vccd1 _06978_/A
+ sky130_fd_sc_hd__a22o_2
XANTENNA__07071__C _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09435_/Y sky130_fd_sc_hd__nor2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06578_ reg1_val[24] _06578_/B vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ _09367_/B _09366_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__and2b_1
X_09297_ _09073_/X _09092_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__mux2_1
XANTENNA_40 reg2_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08317_ _08318_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08317_/X sky130_fd_sc_hd__and2_1
XFILLER_0_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_73 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _08248_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08369_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12714__A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12899__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ hold289/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10469_/C sky130_fd_sc_hd__or2_1
XFILLER_0_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08016__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ _11068_/A _08179_/B vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10359__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__A1 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _11308_/B _11190_/B vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07775__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _11794_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11859__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _11033_/A _10068_/X _10071_/Y _11135_/S vssd1 vssd1 vccd1 vccd1 _10072_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ fanout71/X fanout14/X fanout52/X fanout76/X vssd1 vssd1 vccd1 vccd1 _10975_/B
+ sky130_fd_sc_hd__o22a_1
X_12713_ hold21/X _12720_/B _12712_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__o211a_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10834__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ reg1_val[29] _12656_/A vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12575_ _12578_/B _12575_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
XANTENNA__07463__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06606__B _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _11433_/Y _11437_/B _11435_/B vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08007__A2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _11663_/A fanout7/X fanout5/X fanout76/X vssd1 vssd1 vccd1 vccd1 _11458_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11388_ _11459_/B _11388_/B vssd1 vssd1 vccd1 vccd1 _11390_/C sky130_fd_sc_hd__xnor2_1
X_10408_ _10406_/X _10408_/B vssd1 vssd1 vccd1 vccd1 _10425_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13127_ _13253_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_10339_ _10809_/A _10339_/B vssd1 vssd1 vccd1 vccd1 _10339_/X sky130_fd_sc_hd__or2_1
XANTENNA__11562__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13080_/A hold284/X vssd1 vssd1 vccd1 vccd1 _13242_/D sky130_fd_sc_hd__and2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07518__A1 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _11988_/Y _11989_/X _12008_/X vssd1 vssd1 vccd1 vccd1 _12009_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__07518__B2 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06726__C1 _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ _07660_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _07661_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10825__A1 _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07481_ _09885_/A _07287_/X _07291_/Y _09880_/B2 vssd1 vssd1 vccd1 vccd1 _07482_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _09221_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__and2_1
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _09151_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _09151_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09082_ reg1_val[14] reg1_val[17] _09092_/S vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ _08149_/A _08149_/B _08149_/C vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08033_ _08262_/A _08032_/B _08029_/Y vssd1 vssd1 vccd1 vccd1 _08853_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout110_A _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A _07847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09843__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _10132_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09986_/C sky130_fd_sc_hd__or2_1
X_08935_ _08935_/A _08935_/B vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07363__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _07827_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__nand2b_1
X_08797_ _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__nand2_1
X_07748_ _07819_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12266__B1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07679_ _10156_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08485__A2 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ _10570_/A _10568_/X _10586_/S vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _09727_/A fanout17/X fanout9/X _08798_/B vssd1 vssd1 vccd1 vccd1 _09419_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09349_ _09324_/A _09330_/Y _09333_/Y _09145_/Y _09348_/Y vssd1 vssd1 vccd1 vccd1
+ _09349_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ _12361_/A _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10229__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08922__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ _11312_/A _11312_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__nand2_1
X_12291_ _12290_/A _12290_/B _12290_/C vssd1 vssd1 vccd1 vccd1 _12291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _11129_/Y _11133_/B _11131_/B vssd1 vssd1 vccd1 vccd1 _11246_/A sky130_fd_sc_hd__o21a_1
X_11173_ _11656_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11177_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10124_ _10125_/B _10125_/C _10607_/A vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__a21o_1
X_10055_ _10449_/A _10447_/A _10053_/X _10054_/Y _09061_/X vssd1 vssd1 vccd1 vccd1
+ _10091_/A sky130_fd_sc_hd__a311oi_2
XANTENNA__07273__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__B2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10957_ _10957_/A _11296_/A _10957_/C vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__or3_1
XFILLER_0_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10283__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12627_ reg1_val[26] _12656_/A vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__or2_1
X_10888_ _10778_/A _10778_/B _10777_/A vssd1 vssd1 vccd1 vccd1 _10896_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ reg1_val[12] _12559_/B vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__or2_1
XFILLER_0_53_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12489_ _12496_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__and2_1
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11509_ _11509_/A _11509_/B _11547_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__or3_1
XFILLER_0_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07065_/A _07028_/C _07058_/B1 vssd1 vssd1 vccd1 vccd1 _06983_/B sky130_fd_sc_hd__o21ai_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _08729_/A _08752_/A _08713_/Y vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__a21bo_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08651_/A _08651_/B vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__xnor2_2
X_07602_ _07255_/A _06585_/B _06592_/B _07068_/A _09495_/A vssd1 vssd1 vccd1 vccd1
+ _07604_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08582_ _08589_/A _08589_/B vssd1 vssd1 vccd1 vccd1 _08582_/X sky130_fd_sc_hd__or2_1
X_07533_ _07533_/A _07671_/A _07533_/C vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__and3_1
XANTENNA__07911__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07464_ _07689_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout158_A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12248__B _12248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _10481_/A fanout68/X fanout65/X _07000_/A vssd1 vssd1 vccd1 vccd1 _09204_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ _07395_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _07396_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_91_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09134_ _11696_/A _09130_/Y _09133_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _09134_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07427__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09065_ _11238_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09065_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07358__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ _08430_/B _08715_/A2 _08735_/B1 fanout79/X vssd1 vssd1 vccd1 vccd1 _08017_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12723__A1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10734__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__and2_1
X_08918_ _11271_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09687_/A _09687_/B _09688_/Y vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__o21ai_4
X_08849_ _08370_/A _08370_/B _08848_/X vssd1 vssd1 vccd1 vccd1 _08849_/X sky130_fd_sc_hd__o21a_1
X_11860_ _09293_/A _10340_/Y _10350_/Y _09330_/A _11859_/X vssd1 vssd1 vccd1 vccd1
+ _11860_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09655__A1 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__or2_1
X_11791_ _11713_/A _11788_/X _11789_/Y _11790_/X vssd1 vssd1 vccd1 vccd1 dest_val[22]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10742_ _11656_/A _10742_/B vssd1 vssd1 vccd1 vccd1 _10744_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ _10673_/A _10673_/B vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09407__A1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B2 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07418__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ reg1_val[14] curr_PC[14] _12444_/S vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _12517_/B _12344_/B vssd1 vssd1 vccd1 vccd1 _12354_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12274_ hold301/A _12304_/B1 _12272_/Y _12273_/Y _09810_/A vssd1 vssd1 vccd1 vccd1
+ _12274_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11225_ _11226_/A _11226_/B _11226_/C vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11156_ _11156_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _11157_/B sky130_fd_sc_hd__and2_2
X_10107_ _11654_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__xnor2_4
X_11087_ _11212_/B _11087_/B _11088_/B vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__and3_1
X_10038_ _10038_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08697__A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__B1 _11149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ _11988_/A _11988_/B _09498_/A vssd1 vssd1 vccd1 vccd1 _11989_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11453__A1 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09949__A2 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ reg1_val[28] _07180_/B vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__A _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10964__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__B1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A1 _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07906__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _11636_/S _09819_/Y _09820_/X _09818_/X vssd1 vssd1 vccd1 vccd1 dest_val[4]
+ sky130_fd_sc_hd__a31o_4
XANTENNA__12531__B _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ _09750_/Y _09752_/B vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__and2b_1
X_06964_ fanout79/X _12694_/A _08430_/B _10490_/B2 vssd1 vssd1 vccd1 vccd1 _06965_/B
+ sky130_fd_sc_hd__o22a_1
X_08703_ _08696_/A _08696_/B _08702_/Y vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__o21bai_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06895_ instruction[17] _06890_/X _09135_/B _06527_/X vssd1 vssd1 vccd1 vccd1 _06895_/X
+ sky130_fd_sc_hd__a31o_1
X_09683_ _09684_/B _09683_/B vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08634_ _08634_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _08656_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08755_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _08603_/A sky130_fd_sc_hd__or2_1
X_07516_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout13 _07153_/X vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__buf_8
XFILLER_0_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11163__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout24 _10208_/B vssd1 vssd1 vccd1 vccd1 _11620_/B sky130_fd_sc_hd__buf_4
Xfanout46 _07187_/Y vssd1 vssd1 vccd1 vccd1 _07391_/B sky130_fd_sc_hd__buf_4
XFILLER_0_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08496_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08513_/A sky130_fd_sc_hd__xnor2_1
Xfanout35 _07305_/X vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__buf_8
XFILLER_0_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07447_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__and2_1
Xfanout68 _12712_/A vssd1 vssd1 vccd1 vccd1 fanout68/X sky130_fd_sc_hd__clkbuf_4
Xfanout57 _12716_/A vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout79 _06957_/X vssd1 vssd1 vccd1 vccd1 fanout79/X sky130_fd_sc_hd__buf_8
X_07378_ _07478_/A _07378_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09568__A _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12944__A1 _07131_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ reg1_val[3] reg1_val[28] _09120_/S vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06704__B _06931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ _09048_/A _09048_/B _09048_/C _09048_/D vssd1 vssd1 vccd1 vccd1 _09049_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10955__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout90_A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _11010_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11012_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11380__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ hold60/A _12664_/A rst vssd1 vssd1 vccd1 vccd1 _12961_/Y sky130_fd_sc_hd__a21oi_1
X_12892_ _13085_/A hold238/X vssd1 vssd1 vccd1 vccd1 _13187_/D sky130_fd_sc_hd__and2_1
X_11912_ _12112_/A _11909_/Y _11910_/X _12113_/A vssd1 vssd1 vccd1 vccd1 _11913_/B
+ sky130_fd_sc_hd__o31a_1
X_11843_ _06837_/A _11842_/X _09139_/Y vssd1 vssd1 vccd1 vccd1 _11843_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _12302_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08300__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10725_ _11296_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _12309_/B1 _10586_/X _06699_/B vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ _12326_/A _12326_/B vssd1 vssd1 vccd1 vccd1 _12327_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10410__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ _12290_/B _12257_/B vssd1 vssd1 vccd1 vccd1 _12257_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12188_ hold237/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12275_/C sky130_fd_sc_hd__or2_1
X_11208_ _11089_/B _11096_/B _11087_/X vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__a21o_1
X_11139_ hold267/A _12000_/A2 _11252_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11139_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10152__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A3 _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _10920_/A _06960_/A vssd1 vssd1 vccd1 vccd1 _06681_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08350_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__and2_1
XFILLER_0_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _11271_/A _07301_/B vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ _08272_/A _08272_/B _08272_/C vssd1 vssd1 vccd1 vccd1 _08281_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07232_ reg1_val[17] _07232_/B vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12926__A1 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ _07639_/B _07163_/B vssd1 vssd1 vccd1 vccd1 _07203_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12526__B _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__C fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ reg1_val[26] _07263_/C _07176_/C _07128_/A vssd1 vssd1 vccd1 vccd1 _07095_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout203 _09153_/X vssd1 vssd1 vccd1 vccd1 _12277_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout214 _06890_/X vssd1 vssd1 vccd1 vccd1 _12303_/A sky130_fd_sc_hd__clkbuf_8
Xfanout247 _09342_/X vssd1 vssd1 vccd1 vccd1 _12304_/B1 sky130_fd_sc_hd__buf_4
X_09804_ hold194/A hold247/A _13160_/Q hold189/A vssd1 vssd1 vccd1 vccd1 _10077_/C
+ sky130_fd_sc_hd__or4_2
Xfanout236 _07099_/A vssd1 vssd1 vccd1 vccd1 _10924_/S sky130_fd_sc_hd__clkbuf_4
Xfanout225 _12668_/A vssd1 vssd1 vccd1 vccd1 _09313_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout269 _13070_/B2 vssd1 vssd1 vccd1 vccd1 _12885_/A2 sky130_fd_sc_hd__buf_4
Xfanout258 _06848_/Y vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__buf_4
X_07996_ _07996_/A vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__inv_2
X_06947_ _06978_/B _06944_/Y _06945_/Y _06943_/Y vssd1 vssd1 vccd1 vccd1 _06947_/X
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__07581__A2 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _09736_/A _09736_/B vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09858__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _09145_/Y _09621_/X _09622_/Y _09665_/X vssd1 vssd1 vccd1 vccd1 _09666_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07869__B1 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B2 _07015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06878_ instruction[15] _06850_/Y _06877_/X _12498_/C vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__07371__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08530__A1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _08617_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _08625_/B sky130_fd_sc_hd__nor2_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09441_/A _09440_/B _09438_/Y vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__a21o_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08548_ _08546_/A _08576_/A _08591_/A vssd1 vssd1 vccd1 vccd1 _08560_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07097__A1 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ _08714_/A _08479_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11490_ _11491_/A _11491_/B _11491_/C vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10640__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ fanout64/X fanout37/X _08233_/B _11876_/A vssd1 vssd1 vccd1 vccd1 _10511_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10443_/A _10443_/B _10443_/C vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08046__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13160_ _13169_/CLK _13160_/D vssd1 vssd1 vccd1 vccd1 _13160_/Q sky130_fd_sc_hd__dfxtp_1
X_10372_ _10371_/A _10371_/B _10371_/C vssd1 vssd1 vccd1 vccd1 _10373_/B sky130_fd_sc_hd__a21o_1
X_13091_ _13091_/A _13091_/B vssd1 vssd1 vccd1 vccd1 _13091_/Y sky130_fd_sc_hd__xnor2_1
X_12111_ _12112_/A _12258_/B _12258_/A vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12042_ _11976_/A _11972_/A _11974_/B vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__a21o_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11068__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12944_ _07131_/Y _12962_/B2 hold123/X vssd1 vssd1 vccd1 vccd1 _13213_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12875_ hold168/X _12885_/A2 _12885_/B1 hold210/A vssd1 vssd1 vccd1 vccd1 hold169/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06609__B _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11827_/B _11827_/A vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__and2b_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08285__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11757_ _11757_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ hold277/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10820_/B sky130_fd_sc_hd__or2_1
XFILLER_0_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11688_ _06792_/X _11687_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11689_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09001__A _09001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10639_ _10639_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ reg1_val[31] _07184_/B _12309_/B1 vssd1 vssd1 vccd1 vccd1 _12309_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07456__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07959_/C sky130_fd_sc_hd__xnor2_1
X_06801_ reg1_val[29] _06801_/B vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__nand2_1
X_07781_ _07779_/A _07779_/B _07862_/A vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__o21bai_2
X_06732_ reg1_val[5] _06928_/C vssd1 vssd1 vccd1 vccd1 _06732_/X sky130_fd_sc_hd__or2_1
X_09520_ _09523_/A vssd1 vssd1 vccd1 vccd1 _09520_/Y sky130_fd_sc_hd__inv_2
X_06663_ reg2_val[15] _06748_/B vssd1 vssd1 vccd1 vccd1 _06663_/X sky130_fd_sc_hd__and2_1
X_09451_ _09452_/B _09452_/A vssd1 vssd1 vccd1 vccd1 _09451_/Y sky130_fd_sc_hd__nand2b_1
X_06594_ _12056_/A _12117_/A _11988_/A _11918_/A vssd1 vssd1 vccd1 vccd1 _06596_/A
+ sky130_fd_sc_hd__or4_1
X_08402_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08402_/X sky130_fd_sc_hd__and2b_1
X_09382_ _09383_/A _09383_/B vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10870__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08333_ _09313_/S _08333_/B vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__or2_1
XFILLER_0_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout238_A _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _07216_/A _07216_/B _07216_/C vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__o21a_1
X_08195_ _08195_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _07147_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07146_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07077_ _07078_/B _07078_/C _08276_/A vssd1 vssd1 vccd1 vccd1 _07079_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07003__B2 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A1 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__A1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__B2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _07979_/A _07979_/B vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__nand2_1
X_09718_ _11183_/A _09718_/B vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12835__B1 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout53_A _07112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _10991_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__or2_1
X_09649_ reg1_val[2] _06749_/X _09494_/Y vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__a21o_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ hold162/A vssd1 vssd1 vccd1 vccd1 _12660_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11611_ _06837_/D _11610_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11611_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ _12591_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_38_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07040__S _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11810__B2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11542_ _10450_/A _11514_/Y _11515_/X _11541_/Y vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11810__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11473_ _11473_/A _11473_/B vssd1 vssd1 vccd1 vccd1 _11474_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ _13217_/CLK hold105/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dfxtp_1
X_10424_ _10424_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__xnor2_1
X_13143_ _13254_/CLK _13143_/D vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10377__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__B2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12182__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10355_ curr_PC[7] _10354_/C curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10355_/Y sky130_fd_sc_hd__a21oi_2
X_13074_ hold291/X _13073_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10118_/A _10118_/B _10116_/A vssd1 vssd1 vccd1 vccd1 _10288_/B sky130_fd_sc_hd__a21o_1
X_12025_ _12026_/A _12026_/B vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__and2_1
XANTENNA__11629__A1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ _13204_/Q _12665_/A _12955_/B1 hold141/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold142/A sky130_fd_sc_hd__o221a_1
X_12858_ _13071_/A hold187/X vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10852__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A_N _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _11885_/A _11809_/B vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ hold53/X hold249/X vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__and2b_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__A _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10604__A2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__B2 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07481__A1 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ _07000_/A vssd1 vssd1 vccd1 vccd1 _07000_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09222__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _08952_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08953_/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08882_ _08985_/A _08985_/B _09058_/B _08880_/Y _08881_/A vssd1 vssd1 vccd1 vccd1
+ _08982_/A sky130_fd_sc_hd__a311o_4
X_07902_ _07902_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07967_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11868__A1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _10099_/A1 _10009_/A _09725_/B2 _12702_/A vssd1 vssd1 vccd1 vccd1 _07834_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08733__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _10853_/A _07764_/B _07764_/C vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ hold296/A _09503_/B vssd1 vssd1 vccd1 vccd1 _09503_/Y sky130_fd_sc_hd__xnor2_1
X_06715_ _07123_/A reg1_val[7] vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__and2b_1
X_07695_ _07695_/A _07695_/B _07695_/C vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06646_ _06646_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _06646_/X sky130_fd_sc_hd__or2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09434_ _09434_/A _09434_/B vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06577_ reg1_val[24] _06578_/B vssd1 vssd1 vccd1 vccd1 _06579_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12267__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ _11794_/A _09365_/B vssd1 vssd1 vccd1 vccd1 _09366_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_41 reg2_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _09294_/X _09295_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_30 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _08316_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08318_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 reg2_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _08315_/B _08315_/A vssd1 vssd1 vccd1 vccd1 _08248_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08178_ _08813_/B1 fanout37/X _08233_/B _08737_/A2 vssd1 vssd1 vccd1 vccd1 _08179_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10359__B2 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07129_ _07284_/B _07130_/C reg1_val[22] vssd1 vssd1 vccd1 vccd1 _07132_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07775__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10377_/A1 _07513_/B fanout92/X fanout15/X vssd1 vssd1 vccd1 vccd1 _10141_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10071_ _11033_/A _11033_/B vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09921__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10250__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08488__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _11799_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__xnor2_1
X_12712_ _12712_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12712_/Y sky130_fd_sc_hd__nand2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12643_ _12647_/B _12643_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__nor2_8
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ _12574_/A _12574_/B _12574_/C vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07463__B2 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__A1 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11525_ _11523_/Y _11525_/B vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08660__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09917__C _10320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _11633_/C _11455_/Y _11713_/A _11453_/X vssd1 vssd1 vccd1 vccd1 dest_val[18]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__08390__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11387_ _11387_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__or2_1
X_10407_ _10545_/B _10406_/B _10406_/C vssd1 vssd1 vccd1 vccd1 _10408_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _13234_/CLK _13126_/D vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ _09095_/X _09111_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _10339_/B sky130_fd_sc_hd__mux2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ hold283/X _13084_/A2 _13056_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold284/A
+ sky130_fd_sc_hd__a22o_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12008_ _12008_/A _12008_/B _12008_/C _12008_/D vssd1 vssd1 vccd1 vccd1 _12008_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__08715__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__B2 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10269_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _09979_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07484_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10825__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__B1 _07152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _09151_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _09150_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09081_ reg1_val[15] reg1_val[16] _09092_/S vssd1 vssd1 vccd1 vccd1 _09081_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ _11470_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _08149_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _08029_/Y _08032_/B vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06532__B _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__nor2_1
X_08934_ _08934_/A _08934_/B vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__xnor2_1
X_08865_ _08859_/B _08865_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nand2b_1
X_07816_ _07816_/A _07816_/B vssd1 vssd1 vccd1 vccd1 _07827_/B sky130_fd_sc_hd__xnor2_2
X_08796_ _08792_/A _08792_/C _08792_/B vssd1 vssd1 vccd1 vccd1 _08797_/B sky130_fd_sc_hd__o21ai_1
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07678_ fanout79/X _12688_/A _07304_/Y _08430_/B vssd1 vssd1 vccd1 vccd1 _07679_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06629_ instruction[29] _06637_/B vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__and2_4
XFILLER_0_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ _09417_/A _09417_/B vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__nor2_1
X_09348_ _09334_/Y _09335_/X _09347_/X vssd1 vssd1 vccd1 vccd1 _09348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__B2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11310_ _11310_/A vssd1 vssd1 vccd1 vccd1 _11312_/B sky130_fd_sc_hd__inv_2
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12290_ _12290_/A _12290_/B _12290_/C vssd1 vssd1 vccd1 vccd1 _12290_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _11240_/A _11240_/B _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _11950_/A fanout50/X _07988_/B _12095_/A vssd1 vssd1 vccd1 vccd1 _11173_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _07075_/A _07075_/B _07000_/A vssd1 vssd1 vccd1 vccd1 _10125_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_101_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10054_ _10449_/A _10053_/X _10447_/A vssd1 vssd1 vccd1 vccd1 _10054_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08173__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _12089_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10957_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10887_ _10771_/A _10771_/B _10757_/A vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06617__B _06987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ _12626_/A _12630_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12557_ _12562_/B _12557_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_12488_ reg1_val[26] curr_PC[26] _12495_/S vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11508_ _11506_/X _11508_/B vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _11625_/B _09501_/B _11439_/S vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _13109_/A _13109_/B _13109_/C vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__or3_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _06980_/A _06980_/B vssd1 vssd1 vccd1 vccd1 _07028_/C sky130_fd_sc_hd__or2_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07464__A _07689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08650_ _08651_/B _08651_/A vssd1 vssd1 vccd1 vccd1 _08650_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07372__B1 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06714__A3 _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__C _10321_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _09862_/B _07601_/B vssd1 vssd1 vccd1 vccd1 _07608_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ _08579_/A _08579_/B _08627_/A vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__a21oi_1
X_07532_ _12085_/A _07525_/B _07531_/X vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ _06985_/A _12704_/A _12702_/A _06977_/A vssd1 vssd1 vccd1 vccd1 _07464_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06527__B _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _10252_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _07411_/A _07393_/C _07393_/A vssd1 vssd1 vccd1 vccd1 _07395_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07427__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09133_ _09328_/A _09132_/X _11696_/A vssd1 vssd1 vccd1 vccd1 _09133_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07427__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09064_ _12053_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09064_/Y sky130_fd_sc_hd__nor2_2
X_08015_ _08535_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12723__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10734__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _11654_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__xnor2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ fanout80/X fanout42/X _07239_/A _10099_/A1 vssd1 vssd1 vccd1 vccd1 _08918_/B
+ sky130_fd_sc_hd__o22a_1
X_09897_ _09753_/A _09752_/B _09750_/Y vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__a21o_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _08370_/A _08370_/B _08367_/A vssd1 vssd1 vccd1 vccd1 _08848_/X sky130_fd_sc_hd__a21o_1
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _09007_/A sky130_fd_sc_hd__and2_1
X_10810_ _11135_/S _09656_/X _10809_/X vssd1 vssd1 vccd1 vccd1 _10810_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ curr_PC[22] _11866_/C _06847_/X vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_95_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ _11663_/A fanout50/X _07988_/B _11739_/A vssd1 vssd1 vccd1 vccd1 _10742_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06874__C1 _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12417_/B _12411_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07418__A1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ _10673_/A _10673_/B vssd1 vssd1 vccd1 vccd1 _10672_/X sky130_fd_sc_hd__and2_1
XANTENNA__09407__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07418__B2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ reg1_val[4] curr_PC[4] _12444_/S vssd1 vssd1 vccd1 vccd1 _12344_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _12304_/B1 _12272_/Y hold301/A vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11224_ _11327_/B _11224_/B vssd1 vssd1 vccd1 vccd1 _11226_/C sky130_fd_sc_hd__or2_1
XFILLER_0_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _11155_/A _11159_/B _11160_/A vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__and3_1
X_10106_ _11387_/A _11564_/A fanout38/X fanout71/X vssd1 vssd1 vccd1 vccd1 _10107_/B
+ sky130_fd_sc_hd__o22a_2
X_11086_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__xor2_1
X_10037_ _10038_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11150__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ _11988_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11989__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ _09330_/A _10925_/X _10938_/Y _09120_/S _10936_/X vssd1 vssd1 vccd1 vccd1
+ _10939_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11453__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__A3 _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12365__A _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12609_ reg1_val[22] _12615_/B vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__or2_1
XANTENNA__08606__B1 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10964__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08909__A1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__B2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07906__B _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A2 _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09820_ curr_PC[4] _09957_/C vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__or2_1
XANTENNA__07194__A _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ _06963_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _06963_/Y sky130_fd_sc_hd__xnor2_4
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09751_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__nand2_1
X_08702_ _08707_/A _08731_/A vssd1 vssd1 vccd1 vccd1 _08702_/Y sky130_fd_sc_hd__nor2_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06894_ _09140_/B _09153_/B vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__or2_2
XANTENNA__07345__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09682_ _11794_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout170_A _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _08634_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _08640_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08564_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08564_/Y sky130_fd_sc_hd__inv_2
X_07515_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout25 _12190_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__clkbuf_4
Xfanout47 _07156_/X vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__buf_6
Xfanout14 fanout15/X vssd1 vssd1 vccd1 vccd1 fanout14/X sky130_fd_sc_hd__buf_8
X_08495_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08495_/X sky130_fd_sc_hd__or2_1
Xfanout36 fanout37/X vssd1 vssd1 vccd1 vccd1 fanout36/X sky130_fd_sc_hd__clkbuf_8
Xfanout69 _07014_/Y vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _11955_/A _07446_/B vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout58 _12716_/A vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__buf_4
XFILLER_0_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _07377_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09568__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ reg1_val[2] reg1_val[29] _09120_/S vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09047_ _11838_/B _11838_/C vssd1 vssd1 vccd1 vccd1 _11914_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__A1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__B2 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12722__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__A1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _06732_/X _12309_/B1 _09141_/Y _09926_/A _09948_/X vssd1 vssd1 vccd1 vccd1
+ _09949_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11380__A1 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _07267_/B _12686_/B hold61/X vssd1 vssd1 vccd1 vccd1 _13221_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12891_ hold225/X _13084_/B2 _13084_/A2 hold233/X vssd1 vssd1 vccd1 vccd1 hold238/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07832__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _12112_/A _11910_/X _11909_/Y vssd1 vssd1 vccd1 vccd1 _11913_/A sky130_fd_sc_hd__o21ai_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _06796_/X _11841_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11842_/X sky130_fd_sc_hd__mux2_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11773_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08300__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10724_ _10957_/A fanout7/X fanout5/X _10876_/A1 vssd1 vssd1 vccd1 vccd1 _10725_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10655_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10776_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ _09147_/X _09141_/Y _10586_/S vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__mux2_1
X_12325_ _12326_/A _12326_/B vssd1 vssd1 vccd1 vccd1 _12333_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12699__A1 _11091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__nand3_1
X_12187_ _12187_/A _12187_/B vssd1 vssd1 vccd1 vccd1 _12195_/C sky130_fd_sc_hd__nor2_1
X_11207_ _11319_/B _11207_/B vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__nor2_1
X_11138_ _12000_/A2 _11252_/B hold267/A vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06630__B _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _11184_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11069_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07300_ _09979_/A _11468_/A _07301_/B vssd1 vssd1 vccd1 vccd1 _07300_/X sky130_fd_sc_hd__and3_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08280_ _08280_/A _08280_/B _08280_/C vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__or3_1
XFILLER_0_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08573__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10634__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ reg1_val[13] reg1_val[16] _07091_/B _07091_/C _07050_/A vssd1 vssd1 vccd1
+ vccd1 _07232_/B sky130_fd_sc_hd__o41a_1
XANTENNA__12095__A _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12926__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07163_/B sky130_fd_sc_hd__and2_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08055__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08055__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07802__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ _07263_/C _07176_/C _07128_/A vssd1 vssd1 vccd1 vccd1 _07103_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout204 _09148_/X vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__buf_4
XANTENNA__12542__B _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout226 _08936_/A vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__buf_8
Xfanout237 _06737_/Y vssd1 vssd1 vccd1 vccd1 _11135_/S sky130_fd_sc_hd__clkbuf_8
X_09803_ _11696_/A _09801_/X _09802_/Y _06889_/Y _09796_/Y vssd1 vssd1 vccd1 vccd1
+ _09817_/C sky130_fd_sc_hd__o311a_1
XFILLER_0_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout248 _09151_/X vssd1 vssd1 vccd1 vccd1 _12313_/A1 sky130_fd_sc_hd__buf_4
Xfanout259 _12080_/A vssd1 vssd1 vccd1 vccd1 _12444_/S sky130_fd_sc_hd__clkbuf_8
X_07995_ _08734_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__xnor2_1
X_06946_ _06943_/Y _06945_/Y _06944_/Y _06978_/B vssd1 vssd1 vccd1 vccd1 _06946_/X
+ sky130_fd_sc_hd__o2bb2a_2
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09858__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ instruction[22] _06887_/B vssd1 vssd1 vccd1 vccd1 _06877_/X sky130_fd_sc_hd__or2_1
X_09665_ _09152_/Y _09645_/X _09660_/X _09664_/X vssd1 vssd1 vccd1 vccd1 _09665_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07869__B2 _06961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _08616_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06541__A1 _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08547_ _08590_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__or2_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10625__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _08670_/A2 _08733_/B1 _08735_/A2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08479_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ _07429_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07521_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07099__A _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08046__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10443_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08046__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _10371_/A _10371_/B _10371_/C vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__and3_1
XANTENNA__11050__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _12738_/X _13090_/B vssd1 vssd1 vccd1 vccd1 _13091_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _12110_/A _12110_/B _12110_/C _12110_/D vssd1 vssd1 vccd1 vccd1 _12258_/B
+ sky130_fd_sc_hd__and4_2
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ _12107_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__or2_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12943_ hold103/X _12662_/A _13112_/B hold122/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold123/A sky130_fd_sc_hd__o221a_1
XANTENNA__07562__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12874_ _13071_/A hold183/X vssd1 vssd1 vccd1 vccd1 _13178_/D sky130_fd_sc_hd__and2_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11825_ _11905_/A _11825_/B vssd1 vssd1 vccd1 vccd1 _11827_/B sky130_fd_sc_hd__or2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08285__B2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08285__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ _11871_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _12309_/B1 _10706_/X _06693_/B vssd1 vssd1 vccd1 vccd1 _10707_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ _06837_/D _11609_/X _06628_/A vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10638_ _10639_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10638_/X sky130_fd_sc_hd__and2_1
XFILLER_0_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ _06777_/Y _10568_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12308_ hold128/A _12306_/X _12307_/Y vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__a21o_1
X_12239_ _09135_/Y _09474_/X _09488_/X _09064_/Y _12238_/X vssd1 vssd1 vccd1 vccd1
+ _12240_/C sky130_fd_sc_hd__a221o_1
XANTENNA__13097__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _06800_/A _07255_/A vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__or2_1
X_07780_ _07861_/A _07861_/B vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__nor2_1
X_06731_ reg1_val[5] _06928_/C vssd1 vssd1 vccd1 vccd1 _06734_/A sky130_fd_sc_hd__nor2_1
X_09450_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07720__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06662_ _06660_/Y _06662_/B vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__nand2b_1
X_08401_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__xor2_1
X_06593_ _06591_/X _06593_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ _11654_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09383_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08332_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12537__B _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07214_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07216_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout133_A _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _08193_/A _08193_/B _08195_/A vssd1 vssd1 vccd1 vccd1 _08194_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09225__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout300_A _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ _07303_/A _07109_/A _07109_/B _06730_/B vssd1 vssd1 vccd1 vccd1 _07147_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09776__A1 _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _07075_/A _07075_/B _06828_/A vssd1 vssd1 vccd1 vccd1 _07078_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07787__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11169__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07979_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13088__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06929_ _07109_/A _06932_/C vssd1 vssd1 vccd1 vccd1 _06979_/A sky130_fd_sc_hd__nor2_2
X_09717_ _11297_/A fanout36/X fanout34/X _11387_/A vssd1 vssd1 vccd1 vccd1 _09718_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09700__A1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ hold257/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__and2_1
XFILLER_0_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09700__B2 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12728__A _12728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10099_/A1 fanout36/X fanout34/X _11297_/A vssd1 vssd1 vccd1 vccd1 _09580_/B
+ sky130_fd_sc_hd__o22a_1
X_11610_ _06790_/X _11609_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ reg1_val[18] _12615_/B vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__nand2_1
X_11541_ _11516_/Y _11517_/X _11540_/Y vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11810__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13012__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11472_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11473_/B sky130_fd_sc_hd__and2_1
X_13211_ _13217_/CLK _13211_/D vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__dfxtp_1
X_10423_ _10424_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__nand2b_1
X_13142_ _13241_/CLK _13142_/D vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07557__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10354_ curr_PC[7] curr_PC[8] _10354_/C vssd1 vssd1 vccd1 vccd1 _10597_/C sky130_fd_sc_hd__and3_2
XANTENNA__10377__A2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13073_ _13073_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13073_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ _10285_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12024_ _12102_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12026_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07950__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ _10850_/A _12926_/A2 hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__o21a_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10837__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ hold186/X _12885_/A2 _12885_/B1 _13170_/Q vssd1 vssd1 vccd1 vccd1 hold187/A
+ sky130_fd_sc_hd__a22o_1
X_11808_ fanout55/X fanout8/X fanout6/X fanout58/X vssd1 vssd1 vccd1 vccd1 _11809_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12788_ hold243/X hold76/X vssd1 vssd1 vccd1 vccd1 _12971_/B sky130_fd_sc_hd__nand2b_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _11739_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _11741_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07769__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ _11183_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__xnor2_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__nor2_2
X_07901_ _07969_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09682__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07832_ _07832_/A _07832_/B vssd1 vssd1 vccd1 vccd1 _07839_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08733__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ hold243/A hold249/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09503_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07763_ _08430_/B _07763_/B vssd1 vssd1 vccd1 vccd1 _07764_/C sky130_fd_sc_hd__or2_1
X_06714_ _06763_/B _06646_/A _12537_/B _06713_/X vssd1 vssd1 vccd1 vccd1 _07123_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _07692_/A _07692_/B _07786_/A vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06645_ instruction[0] instruction[1] _06850_/B instruction[27] pred_val vssd1 vssd1
+ vccd1 vccd1 _12507_/B sky130_fd_sc_hd__o311a_4
XANTENNA_fanout250_A _09146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__and2_1
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ fanout15/X _10117_/A _12684_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _09365_/B
+ sky130_fd_sc_hd__o22a_1
X_06576_ reg2_val[24] _06754_/B _06657_/B1 _06574_/X vssd1 vssd1 vccd1 vccd1 _06578_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10056__A1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12982__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09069_/X _09077_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__mux2_1
XANTENNA_31 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 reg1_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 instruction[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 reg2_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 reg2_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08246_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08177_ _08193_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09068__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _07128_/A _07128_/B vssd1 vssd1 vccd1 vccd1 _07130_/C sky130_fd_sc_hd__and2_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ _07059_/A _07059_/B vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _10073_/S _09478_/X _10069_/Y vssd1 vssd1 vccd1 vccd1 _11033_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12730__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__C1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06684__A_N _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__A _08936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ _11663_/A fanout13/X fanout47/X _11739_/A vssd1 vssd1 vccd1 vccd1 _10973_/B
+ sky130_fd_sc_hd__o22a_1
X_12711_ hold13/X _12720_/B _12710_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o211a_1
XFILLER_0_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12642_ _12642_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__and3_2
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12573_ _12574_/A _12574_/B _12574_/C vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07463__A2 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11524_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08660__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ curr_PC[18] _11454_/B _11636_/S vssd1 vssd1 vccd1 vccd1 _11455_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08660__B2 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10545_/B _10406_/B _10406_/C vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _07300_/X _11385_/B _11385_/Y _11183_/A vssd1 vssd1 vccd1 vccd1 _11459_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13125_ _13260_/CLK _13125_/D vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dfxtp_1
X_10337_ _10337_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ hold287/A _13055_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__mux2_1
X_10268_ _10402_/B _10268_/B vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__nor2_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _09293_/A _10075_/Y _10088_/Y _12073_/B2 _12006_/X vssd1 vssd1 vccd1 vccd1
+ _12008_/D sky130_fd_sc_hd__o221a_1
XANTENNA__08715__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _09626_/X _09631_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _10199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07923__B1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12909_ hold131/X _12662_/A _13112_/B hold146/X _13121_/A vssd1 vssd1 vccd1 vccd1
+ hold147/A sky130_fd_sc_hd__o221a_1
XFILLER_0_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08565__B _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _09072_/X _09079_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08100_ _08098_/A _08098_/B _08099_/Y vssd1 vssd1 vccd1 vccd1 _08154_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08031_ _08031_/A _08031_/B vssd1 vssd1 vccd1 vccd1 _08032_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11538__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08954__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09982_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__and2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ _08933_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08934_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11710__A1 _06987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__nand2_1
X_07815_ _07809_/Y _07813_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _07827_/A sky130_fd_sc_hd__o21ba_1
X_08795_ _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__xor2_1
X_07746_ _07746_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__and2_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07677_ _07832_/A _07677_/B vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__xnor2_1
X_09416_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09417_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06628_ _06628_/A _06628_/B vssd1 vssd1 vccd1 vccd1 _06837_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12018__A2 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09347_ _09336_/B _09501_/B _09340_/Y _09346_/X vssd1 vssd1 vccd1 vccd1 _09347_/X
+ sky130_fd_sc_hd__o211a_1
X_06559_ _06560_/B vssd1 vssd1 vccd1 vccd1 _06559_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07445__A2 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _09279_/B _09279_/A vssd1 vssd1 vccd1 vccd1 _09278_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11910__A _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08229_ _08229_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06723__B _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11240_ _11240_/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11240_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11171_/A _11171_/B vssd1 vssd1 vccd1 vccd1 _11206_/A sky130_fd_sc_hd__nand2_1
X_10122_ _10122_/A _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07905__B1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _10321_/C _10053_/B vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__or2_2
XANTENNA__10261__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10955_ _11297_/A fanout11/X fanout44/X _11295_/B2 vssd1 vssd1 vccd1 vccd1 _10956_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12625_ reg1_val[25] _12656_/A vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12965__B1 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ _12556_/A _12556_/B _12556_/C vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06914__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ _11506_/A _11506_/B _11506_/C vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _12487_/A _12487_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _10938_/A _11437_/Y _12125_/S vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _11370_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13108_ _13111_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _13253_/D sky130_fd_sc_hd__and2_1
XANTENNA__11940__A1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _12757_/X _13039_/B vssd1 vssd1 vccd1 vccd1 _13040_/B sky130_fd_sc_hd__nand2b_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07600_ fanout63/X _09727_/A _08798_/B _12094_/A vssd1 vssd1 vccd1 vccd1 _07601_/B
+ sky130_fd_sc_hd__o22a_2
X_08580_ _08626_/A _08626_/B vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__nor2_1
X_07531_ _07666_/A _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07531_/X sky130_fd_sc_hd__or3_1
XANTENNA__07480__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11456__B1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ _10126_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07393_ _07393_/A _07411_/A _07393_/C vssd1 vssd1 vccd1 vccd1 _07395_/A sky130_fd_sc_hd__and3_1
X_09201_ _06977_/A fanout58/X fanout55/X _06985_/A vssd1 vssd1 vccd1 vccd1 _09202_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ _12499_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07427__A2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12545__B _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09821__B1 _09818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ _09464_/A _09465_/A _10320_/A _09061_/X vssd1 vssd1 vccd1 vccd1 _09063_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08014_ fanout83/X _08689_/B1 _09180_/B2 _08565_/B vssd1 vssd1 vccd1 vccd1 _08015_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07060__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09965_ _10359_/B2 _11564_/A fanout38/X _11387_/A vssd1 vssd1 vccd1 vccd1 _09966_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ _08916_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__xnor2_1
X_09896_ _09896_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__xor2_2
X_08847_ _08371_/Y _09001_/A _08847_/C vssd1 vssd1 vccd1 vccd1 _09048_/B sky130_fd_sc_hd__nand3b_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _08776_/A _08776_/C _08776_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08486__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__B _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07115__A1 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _12086_/A _10740_/B vssd1 vssd1 vccd1 vccd1 _10744_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06722__A_N _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ _10671_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10673_/B sky130_fd_sc_hd__xnor2_2
X_12410_ _12410_/A _12410_/B _12410_/C vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11640__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__B1 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12341_ _12347_/B _12341_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ _13105_/A _12272_/B vssd1 vssd1 vccd1 vccd1 _12272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08379__B1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _11223_/A _11223_/B _11223_/C vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _11153_/A _11150_/X _11151_/X _11153_/Y vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__a22o_4
X_10105_ _10105_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__nor2_2
X_11085_ _11085_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11686__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _09893_/A _09890_/X _09892_/A vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__o21a_2
XANTENNA__06909__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08396__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ _11238_/A _06806_/Y _06814_/X _11986_/X vssd1 vssd1 vccd1 vccd1 _11988_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10938_ _10938_/A vssd1 vssd1 vccd1 vccd1 _10938_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ _10868_/A _10868_/B _10868_/C vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08773__A_N _08784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _12620_/B _12608_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XFILLER_0_14_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08606__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08606__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ _12539_/A _12539_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
XFILLER_0_54_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10964__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08909__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06962_ _06963_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__xor2_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09750_ _09751_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09750_/Y sky130_fd_sc_hd__nor2_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ fanout14/X _10370_/A _07763_/B fanout52/X vssd1 vssd1 vccd1 vccd1 _09682_/B
+ sky130_fd_sc_hd__o22a_1
X_08701_ _08730_/B _08730_/C _08730_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__o21ai_2
X_06893_ _09140_/B _09153_/B vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07345__A1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _08714_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _08563_/A _08563_/B vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__xor2_2
X_07514_ _12085_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08845__A1 _09001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10101__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ _10853_/A _08539_/A _08519_/A vssd1 vssd1 vccd1 vccd1 _08496_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout26 _12223_/A vssd1 vssd1 vccd1 vccd1 _12190_/B sky130_fd_sc_hd__buf_4
X_07445_ _07099_/X _07799_/B _07271_/X _07154_/X vssd1 vssd1 vccd1 vccd1 _07446_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout15 _07106_/X vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__buf_6
Xfanout37 _07302_/Y vssd1 vssd1 vccd1 vccd1 fanout37/X sky130_fd_sc_hd__buf_8
Xfanout59 _07049_/X vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout48 fanout49/X vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__buf_6
X_07376_ _07478_/A _07378_/B vssd1 vssd1 vccd1 vccd1 _07376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _09113_/A _09114_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ _09052_/B _09052_/C vssd1 vssd1 vccd1 vccd1 _11838_/C sky130_fd_sc_hd__or2_1
XFILLER_0_5_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07385__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _06928_/C _12238_/C1 _09147_/X _06734_/B _09947_/Y vssd1 vssd1 vccd1 vccd1
+ _09948_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11380__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout76_A fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__xnor2_1
X_12890_ _13080_/A hold226/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__and2_1
X_11910_ _12110_/A _12110_/B _12110_/C vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__and3_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11767_/A _11765_/X _11782_/S vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__a21o_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11691_/Y _11695_/B _11693_/B vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__o21a_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10723_ _12089_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__xnor2_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ _10654_/A _10654_/B vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__xnor2_1
X_10585_ hold203/A _11781_/B _10703_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _10585_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _12333_/A _12324_/B vssd1 vssd1 vccd1 vccd1 _12326_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07272__B1 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12699__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12290_/B sky130_fd_sc_hd__a21o_1
X_12186_ hold293/A _12304_/B1 _12230_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _12187_/B
+ sky130_fd_sc_hd__a31o_1
X_11206_ _11206_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__and2_1
X_11137_ hold273/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__or2_1
XANTENNA__07575__A1 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ _11068_/A _11068_/B vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _07513_/B fanout92/X _12690_/A fanout14/X vssd1 vssd1 vccd1 vccd1 _10020_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10634__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10634__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _10920_/A _07091_/B _07091_/C _07050_/A vssd1 vssd1 vccd1 vccd1 _07233_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12095__B _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09252__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12139__A1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07176_/C sky130_fd_sc_hd__or2_2
XANTENNA__11347__C1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _09137_/Y vssd1 vssd1 vccd1 vccd1 _12309_/B1 sky130_fd_sc_hd__buf_4
Xfanout216 _13112_/B vssd1 vssd1 vccd1 vccd1 _12955_/B1 sky130_fd_sc_hd__buf_4
Xfanout227 _06764_/X vssd1 vssd1 vccd1 vccd1 _09309_/S sky130_fd_sc_hd__buf_8
Xfanout238 _07108_/C vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__clkbuf_8
X_09802_ _09801_/B _09801_/C _09801_/A vssd1 vssd1 vccd1 vccd1 _09802_/Y sky130_fd_sc_hd__a21oi_1
Xfanout249 _09151_/X vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09624__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07994_ _11295_/B2 _08219_/B _08815_/B _11462_/A vssd1 vssd1 vccd1 vccd1 _07995_/B
+ sky130_fd_sc_hd__o22a_1
X_06945_ _06945_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _06945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__nor2_1
X_06876_ instruction[14] _06850_/Y _06875_/X _12498_/C vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__o211a_4
X_09664_ _09664_/A _09664_/B _09663_/X vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__or3b_1
XANTENNA__07869__A2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__B1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ _08613_/A _08613_/B _08654_/A vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__o21bai_1
X_09595_ _09595_/A _09595_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08546_/A _08576_/A vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07097__A3 _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08477_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08496_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10625__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07428_ _10156_/A _07428_/B vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07359_ _12085_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07361_/C sky130_fd_sc_hd__or2_1
XFILLER_0_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08046__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _10370_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _10371_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10534__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ _08621_/X _09029_/B vssd1 vssd1 vccd1 vccd1 _09030_/B sky130_fd_sc_hd__nand2b_1
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ _12040_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__and2_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 hold299/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08939__A _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ _07875_/A _12962_/B2 hold104/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__o21a_1
XANTENNA__07054__S _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ hold182/X _13070_/B2 _13070_/A2 hold168/X vssd1 vssd1 vccd1 vccd1 hold183/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11824_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11825_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_28_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08285__A2 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ _11755_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__and2_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _09147_/X _09141_/Y _10706_/S vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07493__B1 _07304_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11686_ _11838_/A _09045_/A _09044_/X _12179_/A vssd1 vssd1 vccd1 vccd1 _11686_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _11470_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10568_ _06704_/Y _10453_/X _06706_/B vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06922__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12307_ hold128/A _12306_/X _09152_/Y vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__o21ai_1
X_10499_ _10499_/A vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__inv_2
XFILLER_0_121_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07290__A1_N _06931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _06584_/X _09147_/X _12237_/Y _06586_/B _12238_/C1 vssd1 vssd1 vccd1 vccd1
+ _12238_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09942__C1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__and2_1
XANTENNA__13097__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ reg1_val[5] _06730_/B vssd1 vssd1 vccd1 vccd1 _06730_/Y sky130_fd_sc_hd__nand2_1
X_06661_ reg1_val[16] _06978_/B vssd1 vssd1 vccd1 vccd1 _06662_/B sky130_fd_sc_hd__or2_1
XANTENNA__07720__A1 _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _08714_/A _08400_/B vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__xnor2_1
X_06592_ reg1_val[28] _06592_/B vssd1 vssd1 vccd1 vccd1 _06593_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09380_ _10377_/A1 _11564_/A fanout38/X _10490_/B2 vssd1 vssd1 vccd1 vccd1 _09381_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08331_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08264_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07213_ _07214_/B _07214_/A vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout126_A _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09225__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ _07108_/C _07109_/A _07303_/A _06730_/B vssd1 vssd1 vccd1 vccd1 _07147_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__07787__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__B _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ _07075_/A _07075_/B vssd1 vssd1 vccd1 vccd1 _07075_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07787__B2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11169__B _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09862__B _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _08037_/A vssd1 vssd1 vccd1 vccd1 _07980_/A sky130_fd_sc_hd__inv_2
X_06928_ _07123_/A _07158_/A _06928_/C _07108_/C vssd1 vssd1 vccd1 vccd1 _06932_/C
+ sky130_fd_sc_hd__or4_2
X_09716_ _11184_/A _09716_/B vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ hold257/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06859_ _06850_/B instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _06862_/B sky130_fd_sc_hd__and4b_4
XFILLER_0_96_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12728__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08529_ _08577_/A _08527_/X _08524_/X vssd1 vssd1 vccd1 vccd1 _08533_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _06889_/Y _11528_/X _11539_/Y _11522_/X vssd1 vssd1 vccd1 vccd1 _11540_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10529__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout5_A fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13012__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13210_ _13217_/CLK hold118/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ _10542_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__and2_1
X_13141_ _13241_/CLK _13141_/D vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ _10324_/X _10327_/X _10332_/X _10352_/X _11636_/S vssd1 vssd1 vccd1 vccd1
+ _10353_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _12746_/X _13072_/B vssd1 vssd1 vccd1 vccd1 _13073_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ _12023_/A _12023_/B _12023_/C vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__nor3_1
X_10284_ _11183_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07950__A1 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__B2 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ hold42/X _12665_/A _12955_/B1 _13204_/Q _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold43/A sky130_fd_sc_hd__o221a_1
XANTENNA__10837__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ _13071_/A hold204/X vssd1 vssd1 vccd1 vccd1 _13169_/D sky130_fd_sc_hd__and2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11807_ _11732_/A _11732_/B _11724_/A vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ hold76/X hold243/X vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__and2b_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ _11738_/A _11738_/B vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11669_ _11749_/A _11669_/B vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__and2_1
XFILLER_0_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07218__B1 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07769__A1 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08880_ _08881_/B _08880_/B vssd1 vssd1 vccd1 vccd1 _08880_/Y sky130_fd_sc_hd__nor2_1
X_07900_ _07900_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10525__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07831_ _12694_/A _07000_/A fanout93/X _10481_/A vssd1 vssd1 vccd1 vccd1 _07832_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09174__S _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A0 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _09501_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07762_ _10982_/A _06957_/B _09180_/B2 vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06713_ reg2_val[7] _06748_/B vssd1 vssd1 vccd1 vccd1 _06713_/X sky130_fd_sc_hd__and2_1
X_07693_ _07785_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06644_ _11439_/S _06644_/B vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _09432_/A _09432_/B _09432_/C vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__or3_1
X_06575_ reg2_val[24] _06754_/B _06657_/B1 _06574_/X vssd1 vssd1 vccd1 vccd1 _07029_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ _09578_/A _09363_/B vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__or2_1
X_08314_ _08312_/A _08312_/B _08313_/Y vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_32 reg2_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _09067_/X _09070_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__mux2_1
XANTENNA_10 curr_PC[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_21 reg1_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09997__A2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_65 instruction[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 reg2_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ _08244_/B _08244_/C _08244_/A vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_76 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__B1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08176_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08177_/B sky130_fd_sc_hd__nor2_1
X_07127_ _07132_/A _07132_/B vssd1 vssd1 vccd1 vccd1 _07127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _06578_/B _07065_/A _07065_/B _07058_/B1 vssd1 vssd1 vccd1 vccd1 _07059_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__09873__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08489__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10971_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__xor2_1
X_12710_ _12710_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12710_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08936__B _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12642_/B _12642_/C _12642_/A vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__10259__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12572_ _12572_/A _12578_/A vssd1 vssd1 vccd1 vccd1 _12574_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12992__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11523_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08660__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11454_ curr_PC[18] _11454_/B vssd1 vssd1 vccd1 vccd1 _11633_/C sky130_fd_sc_hd__and2_1
XFILLER_0_34_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10406_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ hold159/X _12663_/C _13121_/A vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__o21a_1
X_10336_ _10334_/Y _10336_/B vssd1 vssd1 vccd1 vccd1 _10337_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13055_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13055_/Y sky130_fd_sc_hd__xnor2_1
X_10267_ _10267_/A _10267_/B vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__nor2_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _07059_/A _06905_/Y _11625_/B _06566_/A _12005_/Y vssd1 vssd1 vccd1 vccd1
+ _12006_/X sky130_fd_sc_hd__o221a_1
X_10198_ _09624_/X _09627_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07923__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12908_ _07053_/B _12686_/B hold132/X vssd1 vssd1 vccd1 vccd1 _13195_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11553__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _13160_/Q _12885_/A2 _12885_/B1 hold247/X vssd1 vssd1 vccd1 vccd1 hold248/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09958__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12983__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13246_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09981_ _11183_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__xnor2_1
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09364__B1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _08861_/X _08863_/B vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07814_ _07898_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__nor2_1
X_08794_ _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _08794_/X sky130_fd_sc_hd__and2b_1
X_07745_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07746_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09667__A1 _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 _07304_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _10957_/A _08606_/A2 _07000_/A fanout80/X vssd1 vssd1 vccd1 vccd1 _07677_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__and2_1
X_06627_ reg1_val[20] _06982_/A vssd1 vssd1 vccd1 vccd1 _06628_/B sky130_fd_sc_hd__nor2_1
X_09346_ _12302_/A _09330_/B _09341_/X _09345_/X vssd1 vssd1 vccd1 vccd1 _09346_/X
+ sky130_fd_sc_hd__o211a_1
X_06558_ reg1_val[27] _07064_/B vssd1 vssd1 vccd1 vccd1 _06560_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12974__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _09277_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07388__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08307_/A _08307_/B _08225_/X vssd1 vssd1 vccd1 vccd1 _08229_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _08160_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__B1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _11169_/A _11296_/A _11169_/C vssd1 vssd1 vccd1 vccd1 _11171_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11638__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _10398_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__xnor2_1
X_10052_ _10309_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07905__A1 _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__B1 _11160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _11296_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ _10885_/A _10885_/B vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12624_ _12624_/A _12630_/A vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12965__A1 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12555_ _12556_/A _12556_/B _12556_/C vssd1 vssd1 vccd1 vccd1 _12562_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08094__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ _11506_/A _11506_/B _11506_/C vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__and3_1
XFILLER_0_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _12484_/A _12477_/B _12481_/A _12481_/B vssd1 vssd1 vccd1 vccd1 _12487_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07841__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11437_ _11437_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11437_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_max_cap256_A _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12193__A2 _09637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__A _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _12086_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13107_ hold245/X _06858_/B _13106_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 _13108_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__xor2_2
X_11299_ _12089_/A _11299_/B vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__xor2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13085_/A hold268/X vssd1 vssd1 vccd1 vccd1 _13238_/D sky130_fd_sc_hd__and2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__A2 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__A _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07759_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_89_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07461_ _12706_/A _10009_/A _09725_/B2 fanout77/X vssd1 vssd1 vccd1 vccd1 _07462_/B
+ sky130_fd_sc_hd__o22a_1
X_07392_ _12668_/A _07391_/B _12142_/A vssd1 vssd1 vccd1 vccd1 _07393_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__12405__A0 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ _09200_/A _09200_/B vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12956__A1 _07187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ _12499_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08085__B1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09062_ _09465_/A _10320_/A _09464_/A vssd1 vssd1 vccd1 vccd1 _09062_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09821__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12842__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08013_ _08019_/B _08019_/A vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__A1 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11458__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__B2 _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _11726_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__xnor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08915_ _06940_/A fanout76/X fanout71/X fanout82/X vssd1 vssd1 vccd1 vccd1 _08916_/B
+ sky130_fd_sc_hd__o22a_1
X_09895_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__xor2_2
X_08846_ _08371_/Y _08846_/B vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__nand2b_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _08776_/A _08776_/C _08776_/B vssd1 vssd1 vccd1 vccd1 _08777_/Y sky130_fd_sc_hd__a21oi_1
X_07728_ _07735_/B _07735_/C _07735_/A vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07115__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07659_ _07660_/A _07662_/A _07660_/C vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _10671_/B _10671_/A vssd1 vssd1 vccd1 vccd1 _10670_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _12125_/S _09328_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ _12340_/A _12340_/B _12340_/C vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _09293_/B _12270_/Y _12271_/S vssd1 vssd1 vccd1 vccd1 _12271_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08379__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ _11223_/A _11223_/B _11223_/C vssd1 vssd1 vccd1 vccd1 _11327_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11368__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10359__A2_N _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 _10447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ _11153_/A _11265_/C vssd1 vssd1 vccd1 vccd1 _11153_/Y sky130_fd_sc_hd__nor2_1
X_10104_ _10104_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__nor2_1
X_11084_ _11083_/B _11084_/B vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__nand2b_1
X_10035_ _09852_/A _09852_/B _09850_/Y vssd1 vssd1 vccd1 vccd1 _10038_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__12199__A _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _12053_/A _11986_/B vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _10809_/A _09487_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12938__A1 _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06925__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ reg1_val[20] _12615_/B _12603_/A vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08067__B1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ _10868_/A _10868_/B _10868_/C vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__or3_1
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09803__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08606__A2 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ _11230_/B _10797_/X _10798_/Y vssd1 vssd1 vccd1 vccd1 _10799_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__A _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12536_/Y _12538_/B vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _12469_/A vssd1 vssd1 vccd1 vccd1 _12478_/C sky130_fd_sc_hd__inv_2
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__A _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06961_ _10529_/A _06961_/B vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09971__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _09680_/A _09680_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__xor2_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _09309_/S _10252_/A _08700_/C vssd1 vssd1 vccd1 vccd1 _08730_/C sky130_fd_sc_hd__and3_2
XANTENNA__07345__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ _06892_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08542__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _08670_/A2 _08782_/B2 _08813_/B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08632_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08562_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08588_/B sky130_fd_sc_hd__nor2_1
X_07513_ _12668_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _07514_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10101__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08493_ _08518_/A _08518_/B _08518_/C vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__a21oi_1
X_07444_ _07444_/A _07444_/B vssd1 vssd1 vccd1 vccd1 _07506_/A sky130_fd_sc_hd__xor2_1
Xfanout27 _08983_/Y vssd1 vssd1 vccd1 vccd1 _12223_/A sky130_fd_sc_hd__buf_4
XFILLER_0_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout38 _08135_/B vssd1 vssd1 vccd1 vccd1 fanout38/X sky130_fd_sc_hd__buf_6
Xfanout16 _07074_/X vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__10101__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 _07138_/Y vssd1 vssd1 vccd1 vccd1 fanout49/X sky130_fd_sc_hd__buf_8
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07375_ _07375_/A _07375_/B vssd1 vssd1 vccd1 vccd1 _07378_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06554__B _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ reg1_val[1] reg1_val[30] _09120_/S vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09045_ _09045_/A _09045_/B _09045_/C _11608_/C vssd1 vssd1 vccd1 vccd1 _09052_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11365__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ hold285/A _09945_/X _09946_/Y vssd1 vssd1 vccd1 vccd1 _09947_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09881__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09876_/Y _09878_/B vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__and2b_1
X_08829_ _09009_/A _09009_/B _08803_/X vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__o21a_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A _11840_/B vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__or2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11769_/Y _11771_/B vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08297__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ fanout81/X fanout11/X fanout44/X _11169_/A vssd1 vssd1 vccd1 vccd1 _10723_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _10654_/A _10654_/B vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__and2_1
X_10584_ _11781_/B _10703_/B hold203/A vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _12502_/B _12323_/B vssd1 vssd1 vccd1 vccd1 _12324_/B sky130_fd_sc_hd__or2_1
XANTENNA__07272__A1 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07272__B2 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11356__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ _12290_/A _12254_/B vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _12304_/B1 _12230_/B hold293/A vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08221__B1 _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _11206_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__nor2_1
X_11136_ _11133_/Y _11135_/X _11696_/A vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09721__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _12148_/A fanout37/X _08233_/B _12201_/A vssd1 vssd1 vccd1 vccd1 _11068_/B
+ sky130_fd_sc_hd__o22a_1
X_10018_ _12029_/B _10018_/B vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11969_ _11969_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10634__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07160_ _11955_/A _07160_/B vssd1 vssd1 vccd1 vccd1 _07162_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11044__C1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09966__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _10920_/A _07091_/B _07091_/C _07091_/D vssd1 vssd1 vccd1 vccd1 _07263_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA__09252__A2 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12392__A _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout217 _06857_/Y vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__buf_4
Xfanout228 _09479_/S vssd1 vssd1 vccd1 vccd1 _09633_/S sky130_fd_sc_hd__clkbuf_8
X_09801_ _09801_/A _09801_/B _09801_/C vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__and3_1
Xfanout206 _12113_/A vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__buf_4
Xfanout239 _07108_/C vssd1 vssd1 vccd1 vccd1 _10203_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__11736__A _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_1
X_09732_ _09732_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12311__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06944_ _06979_/A _06943_/B _07289_/B vssd1 vssd1 vccd1 vccd1 _06944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06875_ instruction[21] _06887_/B vssd1 vssd1 vccd1 vccd1 _06875_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout273_A hold177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _06745_/Y _09138_/X _09501_/B _06834_/B _09662_/X vssd1 vssd1 vccd1 vccd1
+ _09663_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09206__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__A1 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08614_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__nor2_1
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09595_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12075__A1 _06890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08590_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08507_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10625__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07427_ _12694_/A _10852_/B2 fanout92/X fanout78/X vssd1 vssd1 vccd1 vccd1 _07428_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07358_ _12085_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07361_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09779__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__A _08784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__S _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ _07289_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _07295_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_33_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _10913_/B _10913_/C vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__nand2_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__buf_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12941_ hold155/A _12665_/A _12955_/B1 hold103/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold104/A sky130_fd_sc_hd__o221a_1
X_12872_ _13062_/A hold180/X vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__and2_1
XANTENNA__08955__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__and2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11813__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ _11755_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10705_ _13170_/Q _11781_/B _10817_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _10705_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A1 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ _11838_/A _09044_/X _09045_/A vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10636_ _11739_/A fanout41/X _08135_/B fanout64/X vssd1 vssd1 vccd1 vccd1 _10637_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08690__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ _10449_/A _09023_/A _09023_/B _12179_/A vssd1 vssd1 vccd1 vccd1 _10567_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06922__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _13189_/Q _12275_/X _12190_/B vssd1 vssd1 vccd1 vccd1 _12306_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10498_ _12086_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__xnor2_1
X_12237_ _06584_/X _09501_/B _09138_/X vssd1 vssd1 vccd1 vccd1 _12237_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10001__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ _12214_/B _12168_/B vssd1 vssd1 vccd1 vccd1 _12258_/C sky130_fd_sc_hd__or2_1
X_12099_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12100_/B sky130_fd_sc_hd__nor2_1
X_11119_ _11230_/C _10909_/B _11230_/D _11232_/A vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__a31o_1
X_06660_ _07233_/A _06945_/A vssd1 vssd1 vccd1 vccd1 _06660_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07720__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ reg1_val[28] _06592_/B vssd1 vssd1 vccd1 vccd1 _06591_/X sky130_fd_sc_hd__and2_1
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08330_ _08741_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08261_ _08261_/A _08261_/B vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07212_ _07082_/A _07081_/B _07081_/A vssd1 vssd1 vccd1 vccd1 _07214_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08192_ _08170_/A _08170_/B _08168_/X vssd1 vssd1 vccd1 vccd1 _08195_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__09225__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _07639_/A _07143_/B vssd1 vssd1 vccd1 vccd1 _07162_/A sky130_fd_sc_hd__or2_1
XFILLER_0_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08433__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _07075_/A _07075_/B vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12850__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07976_ _07976_/A _07976_/B vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10370__A _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06927_ _07099_/A _09634_/A _07186_/A _09309_/S vssd1 vssd1 vccd1 vccd1 _07109_/A
+ sky130_fd_sc_hd__or4_4
X_09715_ fanout78/X fanout74/X fanout68/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _09716_/B
+ sky130_fd_sc_hd__o22a_1
X_09646_ hold296/A hold243/A hold249/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09648_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06858_ hold159/A _06858_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
XFILLER_0_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10846__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ _06641_/Y _06788_/X _11521_/A vssd1 vssd1 vccd1 vccd1 _06790_/B sky130_fd_sc_hd__a21o_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__xor2_1
X_08459_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08459_/X sky130_fd_sc_hd__and2_1
XANTENNA__08672__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _11470_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ _10421_/A _10421_/B _10421_/C vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__or3_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _13251_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_10352_ _12073_/B2 _10340_/Y _10341_/X _06890_/X _10351_/X vssd1 vssd1 vccd1 vccd1
+ _10352_/X sky130_fd_sc_hd__o221a_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08015__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ _13071_/A _13071_/B vssd1 vssd1 vccd1 vccd1 _13245_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12022_ _12023_/A _12023_/B _12023_/C vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__o21a_1
X_10283_ _11663_/A fanout36/X fanout34/X _11739_/A vssd1 vssd1 vccd1 vccd1 _10284_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11376__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12287__A1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _06922_/B _12686_/B hold137/X vssd1 vssd1 vccd1 vccd1 _13203_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__10837__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ hold197/X _12885_/A2 _12885_/B1 hold186/X vssd1 vssd1 vccd1 vccd1 hold204/A
+ sky130_fd_sc_hd__a22o_1
X_12786_ hold296/A hold72/X vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__nand2b_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11806_ _11806_/A _11806_/B vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ _11738_/B _11738_/A vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__and2b_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08663__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ _11668_/A _11668_/B _11668_/C vssd1 vssd1 vccd1 vccd1 _11669_/B sky130_fd_sc_hd__or3_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07218__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ _11600_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11599_/X sky130_fd_sc_hd__a21o_1
X_10619_ _10517_/A _10517_/B _10514_/A vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07769__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06729__B1 _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10525__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07850_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_47_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12278__A1 _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _07832_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__xnor2_1
X_09500_ hold247/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09500_/Y sky130_fd_sc_hd__xnor2_1
X_06712_ _06710_/Y _06712_/B vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09143__A1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07692_ _07692_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08595__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06643_ reg1_val[18] _06980_/B vssd1 vssd1 vccd1 vccd1 _06644_/B sky130_fd_sc_hd__or2_1
X_09431_ _09432_/A _09432_/B _09432_/C vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06574_ _06613_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _06574_/X sky130_fd_sc_hd__or2_1
X_09362_ _09361_/B _09362_/B vssd1 vssd1 vccd1 vccd1 _09363_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07004__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08313_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout236_A _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_11 curr_PC[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg1_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 reg2_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__B _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07939__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08244_/A _08244_/B _08244_/C vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__and3_1
XFILLER_0_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_77 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__and2_1
XFILLER_0_6_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10213__B1 _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06562__B _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ reg1_val[21] _07284_/B _07126_/C vssd1 vssd1 vccd1 vccd1 _07132_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ _08798_/B vssd1 vssd1 vccd1 vccd1 _07057_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09134__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _07959_/A _07959_/B _07959_/C vssd1 vssd1 vccd1 vccd1 _07960_/B sky130_fd_sc_hd__or3_1
X_10970_ _11470_/A _10970_/B vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__xnor2_1
X_09629_ _09625_/X _09628_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _09629_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12640_/A _12640_/B _12640_/C vssd1 vssd1 vccd1 vccd1 _12642_/C sky130_fd_sc_hd__or3_2
XFILLER_0_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ reg1_val[14] _12571_/B vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ _11521_/A _11521_/B _11521_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10452__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12729__C1 _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ _06980_/B _12280_/A _06907_/A _11452_/X vssd1 vssd1 vccd1 vccd1 _11453_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _10403_/B _10403_/C _10403_/A vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__a21oi_1
X_13123_ hold23/X hold162/A _13122_/X _13121_/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o211a_1
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11384_ _11491_/B _11384_/B vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__and2_1
XFILLER_0_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10335_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13054_ _12752_/X _13054_/B vssd1 vssd1 vccd1 vccd1 _13055_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11704__A0 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10266_ _10267_/A _10267_/B vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__and2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12005_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12005_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07384__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07923__A2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06928__A _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ hold110/X _12662_/A _13112_/B hold131/X _13013_/A vssd1 vssd1 vccd1 vccd1
+ hold132/A sky130_fd_sc_hd__o221a_1
XFILLER_0_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _13085_/A hold190/X vssd1 vssd1 vccd1 vccd1 _13160_/D sky130_fd_sc_hd__and2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12769_ hold11/X hold255/X vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__and2b_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12983__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09980_ fanout71/X fanout36/X fanout34/X fanout76/X vssd1 vssd1 vccd1 vccd1 _09981_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07494__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08931_/X sky130_fd_sc_hd__and2_1
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _08861_/A _08866_/A _08861_/C vssd1 vssd1 vccd1 vccd1 _08863_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09364__B2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _07813_/A _07813_/B vssd1 vssd1 vccd1 vccd1 _07898_/B sky130_fd_sc_hd__xor2_1
X_08793_ _08792_/A _08797_/A vssd1 vssd1 vccd1 vccd1 _08795_/B sky130_fd_sc_hd__nand2b_1
X_07744_ _08880_/B _07744_/B vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__and2_2
XFILLER_0_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09667__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07695_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07678__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__B _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ _11625_/A vssd1 vssd1 vccd1 vccd1 _06628_/A sky130_fd_sc_hd__inv_2
X_09414_ _11184_/A _09414_/B vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _12313_/A1 _09343_/X _09344_/Y _06905_/Y _09479_/S vssd1 vssd1 vccd1 vccd1
+ _09345_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ reg1_val[27] _07064_/B vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__and2_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12974__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ _08971_/A _08971_/B _08969_/Y vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _08272_/A _08227_/B vssd1 vssd1 vccd1 vccd1 _08307_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__A _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11934__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _08022_/A _07987_/C _07987_/B vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__A1 _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ _07109_/A _07109_/B vssd1 vssd1 vccd1 vccd1 _08765_/C sky130_fd_sc_hd__and2_1
X_08089_ _08087_/A _08087_/B _08088_/X vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout99_A _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _06977_/A fanout9/X fanout3/X _06985_/A vssd1 vssd1 vccd1 vccd1 _10121_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10051_ _10051_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06708__A3 _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__A2 _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__A1 _10315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _11169_/A fanout7/X fanout5/X fanout81/X vssd1 vssd1 vccd1 vccd1 _10954_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10884_ _10884_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12623_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07579__A _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ _12554_/A _12562_/A vssd1 vssd1 vccd1 vccd1 _12556_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08094__B2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08094__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07841__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _11596_/B _11505_/B vssd1 vssd1 vccd1 vccd1 _11506_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _12485_/A _12485_/B vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__nor2_2
XANTENNA__07841__B2 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ _11345_/A _11342_/Y _11344_/B vssd1 vssd1 vccd1 vccd1 _11437_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_34_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10728__A1 _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__B2 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ fanout64/X fanout14/X fanout52/X _11876_/A vssd1 vssd1 vccd1 vccd1 _11368_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _12832_/C fanout1/X _13104_/Y _13105_/Y vssd1 vssd1 vccd1 vccd1 _13106_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13037_ hold267/X _13084_/A2 _13036_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold268/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09346__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ fanout76/X fanout11/X fanout44/X _11663_/A vssd1 vssd1 vccd1 vccd1 _11299_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _10481_/A _12201_/A fanout9/X _07000_/A vssd1 vssd1 vccd1 vccd1 _10250_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11564__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06658__A _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07460_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07391_ _12668_/A _07391_/B _07391_/C _07391_/D vssd1 vssd1 vccd1 vccd1 _07411_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09130_ _11135_/S _09128_/X _09129_/X vssd1 vssd1 vccd1 vccd1 _09130_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08085__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__B2 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09061_ _09148_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _09061_/X sky130_fd_sc_hd__or2_4
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08012_ _08012_/A _08012_/B vssd1 vssd1 vccd1 vccd1 _08019_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__A _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09585__A1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ _10377_/A1 fanout13/X _07156_/X _10490_/B2 vssd1 vssd1 vccd1 vccd1 _09964_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08914_ _08914_/A _08914_/B vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11144__A1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__and2_1
X_08845_ _09001_/A _08847_/C _08846_/B vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__a21o_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _08776_/A _08776_/B _08776_/C vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__nand3_1
X_07727_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07735_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07660_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08783__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ reg1_val[22] _07028_/B vssd1 vssd1 vccd1 vccd1 _11782_/S sky130_fd_sc_hd__and2_1
X_07589_ _10009_/A _11876_/A _11950_/A _09725_/B2 vssd1 vssd1 vccd1 vccd1 _07590_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09328_ _09328_/A _09328_/B vssd1 vssd1 vccd1 vccd1 _09328_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09812__A2 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout14_A fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__or2_1
XFILLER_0_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12302_/C _12270_/B vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11649__A _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _11327_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11223_/C sky130_fd_sc_hd__or2_1
X_11152_ curr_PC[15] _11152_/B vssd1 vssd1 vccd1 vccd1 _11265_/C sky130_fd_sc_hd__and2_1
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _10104_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__and2_1
X_11083_ _11084_/B _11083_/B vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__nand2b_1
X_10034_ _09838_/A _09838_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11985_ _11935_/A _11916_/X _06579_/A vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10936_ _10931_/Y _10932_/X _10935_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _10936_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07511__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _10867_/A _10867_/B vssd1 vssd1 vccd1 vccd1 _10868_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__06925__B _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ _12604_/Y _12606_/B vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08067__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10798_ _11230_/B _10797_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _10798_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10447__B _10447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ reg1_val[8] _12537_/B vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11071__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ _12468_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _11164_/A _11164_/B _11418_/Y vssd1 vssd1 vccd1 vccd1 _11421_/C sky130_fd_sc_hd__a21o_1
X_12399_ _12559_/B _12400_/B vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07578__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06960_ _06960_/A _06960_/B vssd1 vssd1 vccd1 vccd1 _06960_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11126__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__or2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _08801_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08634_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08542__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _08561_/A _08561_/B vssd1 vssd1 vccd1 vccd1 _08584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07512_ _07916_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10101__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ _10853_/A _08539_/A vssd1 vssd1 vccd1 vccd1 _08518_/C sky130_fd_sc_hd__xnor2_1
X_07443_ _07916_/A _07443_/B vssd1 vssd1 vccd1 vccd1 _07444_/B sky130_fd_sc_hd__xnor2_1
Xfanout17 _07074_/X vssd1 vssd1 vccd1 vccd1 fanout17/X sky130_fd_sc_hd__clkbuf_4
Xfanout28 _11458_/A vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout39 _07291_/Y vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__buf_8
XFILLER_0_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07374_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__nor2_1
X_09113_ _09113_/A vssd1 vssd1 vccd1 vccd1 _09113_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10591__A1_N _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ _11608_/B _11608_/C vssd1 vssd1 vccd1 vccd1 _09044_/X sky130_fd_sc_hd__or2_1
XANTENNA__07281__A2 _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06570__B _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ hold285/A _09945_/X _09150_/Y vssd1 vssd1 vccd1 vccd1 _09946_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13106__A2 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06997__S _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__nand2_1
X_08828_ _08811_/A _08811_/B _09011_/A vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__a21boi_1
X_08759_ _08759_/A _08759_/B _08759_/C vssd1 vssd1 vccd1 vccd1 _08776_/A sky130_fd_sc_hd__or3_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11771_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08297__A1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10721_ _10669_/A _10669_/B _10670_/Y vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__o21ai_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06745__B _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10654_/B sky130_fd_sc_hd__xor2_1
X_10583_ hold197/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10703_/B sky130_fd_sc_hd__or2_1
XFILLER_0_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _12502_/B _12323_/B vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07272__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12253_ _12253_/A _12253_/B _12253_/C vssd1 vssd1 vccd1 vccd1 _12254_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _11319_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11206_/B sky130_fd_sc_hd__or2_1
X_12184_ hold302/A _12184_/B vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11135_ _09167_/Y _11134_/X _11135_/S vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07592__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _11212_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__nand2_1
X_10017_ _12684_/A fanout8/X fanout6/X _10117_/A vssd1 vssd1 vccd1 vccd1 _10018_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09721__A1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06936__A _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _11968_/A _11968_/B vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__and2_1
XANTENNA__06655__B _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _10920_/A curr_PC[13] vssd1 vssd1 vccd1 vccd1 _10921_/A sky130_fd_sc_hd__or2_1
X_11899_ _11899_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07090_ reg1_val[22] reg1_val[23] _12600_/B _07128_/B vssd1 vssd1 vccd1 vccd1 _07091_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11289__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout218 _13070_/A2 vssd1 vssd1 vccd1 vccd1 _12885_/B1 sky130_fd_sc_hd__buf_4
Xfanout229 _06756_/X vssd1 vssd1 vccd1 vccd1 _09479_/S sky130_fd_sc_hd__buf_4
X_09800_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09801_/C sky130_fd_sc_hd__nand2_1
X_07992_ _08801_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__xnor2_4
Xfanout207 _09423_/A vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__buf_12
X_06943_ _06979_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _06943_/Y sky130_fd_sc_hd__nand2_1
X_09731_ _09732_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__and2_1
X_06874_ instruction[13] _06850_/Y _06873_/X _12498_/C vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09662_ _09810_/A _09647_/Y _09648_/X _11625_/B _06747_/B vssd1 vssd1 vccd1 vccd1
+ _09662_/X sky130_fd_sc_hd__o32a_1
XANTENNA__10322__A2 _10447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08653_/B sky130_fd_sc_hd__xnor2_1
X_09593_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__and2_1
XANTENNA__12848__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08544_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11283__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__or2_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _07832_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07357_ fanout15/X _09237_/A _09428_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _07359_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09779__A1 _10320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07254__A2 _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07288_ _07137_/A _07109_/A _06932_/C _07303_/A vssd1 vssd1 vccd1 vccd1 _07295_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ _09027_/A _09027_/B _10800_/B vssd1 vssd1 vccd1 vccd1 _10913_/C sky130_fd_sc_hd__nor3b_1
XANTENNA__11050__A3 _11027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__B1 _07070_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09929_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08301__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ _07286_/B _12686_/B hold156/X vssd1 vssd1 vccd1 vccd1 _13211_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10849__B1 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ hold179/X _13070_/B2 _13070_/A2 hold182/A vssd1 vssd1 vccd1 vccd1 hold180/A
+ sky130_fd_sc_hd__a22o_1
X_11822_ _11822_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__xnor2_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A2 _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _11660_/A _11660_/B _11672_/B _11675_/A vssd1 vssd1 vccd1 vccd1 _11755_/B
+ sky130_fd_sc_hd__a31oi_1
X_10704_ _11781_/B _10817_/B _13170_/Q vssd1 vssd1 vccd1 vccd1 _10704_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11684_ _11683_/A _11683_/B _12113_/A vssd1 vssd1 vccd1 vccd1 _11684_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10635_ _11072_/A _10635_/B vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07587__A _07689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A1 _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12305_ hold126/A _12305_/B vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ _10449_/A _09023_/B _09023_/A vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10497_ fanout81/X fanout14/X fanout52/X _11169_/A vssd1 vssd1 vccd1 vccd1 _10498_/B
+ sky130_fd_sc_hd__o22a_1
X_12236_ hold174/A _12234_/X _12235_/Y vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09942__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _12167_/A _12167_/B _12167_/C vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__and3_1
XANTENNA__10001__A1 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11231_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__08211__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _12146_/B _12098_/B _12099_/B vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__and3_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11049_ _09330_/A _11035_/Y _11036_/X _12303_/A _11048_/X vssd1 vssd1 vccd1 vccd1
+ _11049_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12668__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07181__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ _06592_/B vssd1 vssd1 vccd1 vccd1 _07067_/A sky130_fd_sc_hd__inv_2
XFILLER_0_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08260_ _08261_/A _08261_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07211_ _07354_/A _07354_/B vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__and2b_1
X_08191_ _08109_/A _08110_/B _08186_/B _08187_/Y vssd1 vssd1 vccd1 vccd1 _08196_/A
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__07497__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ _07142_/A _07142_/B vssd1 vssd1 vccd1 vccd1 _07143_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08433__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07073_ _07303_/A _07068_/A _07068_/B _06801_/B vssd1 vssd1 vccd1 vccd1 _07075_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10240__B2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10240__A1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07975_ _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10370__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ _09495_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07289_/B sky130_fd_sc_hd__nand2_2
X_09714_ _09714_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__xor2_2
X_06857_ _12665_/A _12664_/B vssd1 vssd1 vccd1 vccd1 _06857_/Y sky130_fd_sc_hd__nand2_1
X_09645_ hold194/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11482__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06788_ _06787_/A _06787_/B _11431_/A vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11256__B1 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08527_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _08458_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08461_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08672__A1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08672__B2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08389_ _10876_/A1 _09222_/B2 fanout93/X _09422_/A vssd1 vssd1 vccd1 vccd1 _08390_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ _10421_/A _10421_/B _10421_/C vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _11448_/A _10343_/Y _10350_/Y _09124_/S _10349_/X vssd1 vssd1 vccd1 vccd1
+ _10351_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ hold291/X _13070_/A2 _13069_/X _13070_/B2 vssd1 vssd1 vccd1 vccd1 _13071_/B
+ sky130_fd_sc_hd__a22o_1
X_10282_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ _12097_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12023_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12287__A2 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ hold136/X _12665_/A _12955_/B1 hold42/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold137/A sky130_fd_sc_hd__o221a_1
XANTENNA__07870__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12854_ _13071_/A hold198/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__and2_1
XFILLER_0_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12785_ hold72/X hold296/A vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11805_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11806_/B sky130_fd_sc_hd__and2_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11798__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__A1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11736_ _12245_/B _11736_/B vssd1 vssd1 vccd1 vccd1 _11738_/B sky130_fd_sc_hd__xnor2_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08663__B2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _11668_/A _11668_/B _11668_/C vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07218__A2 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11598_ _11600_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10618_ _10535_/A _10535_/B _10532_/A vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10549_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10602_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
XANTENNA__12670__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199_ _13222_/CLK hold121/X vssd1 vssd1 vccd1 vccd1 _13199_/Q sky130_fd_sc_hd__dfxtp_1
X_12219_ _06593_/B _12173_/B _06591_/X vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10525__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07760_ _10377_/A1 _08606_/A2 _06999_/Y _10490_/B2 vssd1 vssd1 vccd1 vccd1 _07761_/B
+ sky130_fd_sc_hd__o22a_1
X_06711_ reg1_val[8] _07137_/A vssd1 vssd1 vccd1 vccd1 _06712_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09143__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07691_ _10126_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__xnor2_1
X_09430_ _12029_/B _09430_/B vssd1 vssd1 vccd1 vccd1 _09432_/C sky130_fd_sc_hd__xnor2_1
X_06642_ reg1_val[18] _06980_/B vssd1 vssd1 vccd1 vccd1 _11439_/S sky130_fd_sc_hd__nand2_1
X_06573_ instruction[34] _06637_/B vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__and2_4
XFILLER_0_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09362_/B _09361_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__and2b_1
X_09292_ _10809_/A _09291_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__o21ai_2
X_08312_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 reg1_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08241_/A _08241_/C _08241_/B vssd1 vssd1 vccd1 vccd1 _08244_/C sky130_fd_sc_hd__o21ai_1
XANTENNA_45 reg2_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 reg2_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 reg2_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _06939_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_67 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__A2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _11470_/A _08174_/B vssd1 vssd1 vccd1 vccd1 _08176_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10213__B2 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07125_ _07284_/B _07126_/C reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07132_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _07056_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07056_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07958_ _07967_/A _07967_/B vssd1 vssd1 vccd1 vccd1 _07958_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08786__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ _12499_/A reg1_val[1] reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07050_/B
+ sky130_fd_sc_hd__or4_2
X_07889_ _07889_/A _07889_/B vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11477__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _09627_/X _09626_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout44_A _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _09559_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ reg1_val[14] _12571_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__or2_1
XFILLER_0_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08645__A1 _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09842__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11521_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06671__A3 _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11452_ _11424_/X _11425_/Y _11428_/Y _09145_/Y _11451_/X vssd1 vssd1 vccd1 vccd1
+ _11452_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11383_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__or2_1
X_10403_ _10403_/A _10403_/B _10403_/C vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__and3_1
X_13122_ hold23/X _12663_/B hold163/A _12664_/A vssd1 vssd1 vccd1 vccd1 _13122_/X
+ sky130_fd_sc_hd__a22o_1
X_10334_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10334_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06959__A1 _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ _13080_/A hold288/X vssd1 vssd1 vccd1 vccd1 _13241_/D sky130_fd_sc_hd__and2_1
XANTENNA__11704__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__A _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _11799_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__xor2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12004_ _06566_/A _09141_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _12005_/B sky130_fd_sc_hd__a21o_1
X_10196_ _10194_/Y _10196_/B vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07384__B2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07384__A1 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__B _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ _09564_/A _12926_/A2 hold111/X vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__o21a_1
XANTENNA__10140__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ hold189/X hold177/X _13084_/A2 _13160_/Q vssd1 vssd1 vccd1 vccd1 hold190/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07105__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12768_ hold277/A hold15/X vssd1 vssd1 vccd1 vccd1 _13014_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_84_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12699_ _11091_/A _12731_/A2 hold48/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13142_/D
+ sky130_fd_sc_hd__o211a_1
X_11719_ _11720_/B _11719_/B vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11943__A1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _06828_/A _11385_/B _07842_/A vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__11297__A _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08861_ _08861_/A _08866_/A _08861_/C vssd1 vssd1 vccd1 vccd1 _08861_/X sky130_fd_sc_hd__and3_1
XANTENNA__09364__A2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08572__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ _08792_/A _08792_/B _08792_/C vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__or3_1
X_07743_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08324__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__and2_1
XFILLER_0_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07678__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06625_ reg1_val[20] _06982_/A vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ _10852_/B2 fanout77/X _11462_/A fanout78/X vssd1 vssd1 vccd1 vccd1 _09414_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12959__B1 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ hold249/A _12304_/B1 hold243/A vssd1 vssd1 vccd1 vccd1 _09344_/Y sky130_fd_sc_hd__a21oi_1
X_06556_ _07064_/B vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _09275_/A _09275_/B vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08226_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08307_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08157_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07108_ _09495_/A _07184_/B _07108_/C vssd1 vssd1 vccd1 vccd1 _07109_/B sky130_fd_sc_hd__and3_1
XANTENNA__09884__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10823__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08088_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ _09420_/A _07039_/B vssd1 vssd1 vccd1 vccd1 _07041_/B sky130_fd_sc_hd__nand2_1
X_10050_ _09777_/A _09777_/B _10049_/X vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10883_ _10883_/A _10883_/B _10883_/C vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__and3_1
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__nand2b_1
X_12553_ reg1_val[11] _12553_/B vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08094__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11504_/A _11504_/B _11504_/C vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__nand3_1
X_12484_ _12484_/A _12484_/B vssd1 vssd1 vccd1 vccd1 _12485_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07841__A2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11435_ _11433_/Y _11435_/B vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10728__A2 _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _12029_/B _11366_/B vssd1 vssd1 vccd1 vccd1 _11370_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _13105_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13105_/Y sky130_fd_sc_hd__nor2_1
X_11297_ _11297_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _11301_/A sky130_fd_sc_hd__nor2_1
X_10317_ _08982_/A _10316_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__a21bo_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13036_ hold273/A _13035_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09346__A2 _09330_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10128_/A _10128_/C _10128_/B vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07357__B2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _10179_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__xor2_4
XANTENNA__10361__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__B fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07390_ _07449_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07391_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08085__A2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10908__B _11230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09060_ _09148_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08011_ _08164_/A _08164_/B _08006_/Y vssd1 vssd1 vccd1 vccd1 _08019_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_25_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07045__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09585__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09962_ _09879_/A _09878_/B _09876_/Y vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__a21oi_2
X_08913_ _08913_/A _08913_/B vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout296_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09893_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09895_/B sky130_fd_sc_hd__xor2_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08472_/Y _09001_/B _09037_/A vssd1 vssd1 vccd1 vccd1 _08847_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ _08759_/A _08759_/B _08759_/C vssd1 vssd1 vccd1 vccd1 _08776_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__06568__B _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07749_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06608_ _06608_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__or2_1
X_07588_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07588_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06539_ _06753_/B _06540_/B vssd1 vssd1 vccd1 vccd1 _06539_/X sky130_fd_sc_hd__and2_2
X_09327_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09328_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10958__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09394_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08209_ _08607_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09189_ _09373_/B _09189_/B vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__or2_2
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07036__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ curr_PC[15] _11152_/B vssd1 vssd1 vccd1 vccd1 _11151_/X sky130_fd_sc_hd__or2_1
X_10102_ _11183_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11082_ _12086_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/B sky130_fd_sc_hd__xnor2_1
X_10033_ _09896_/A _09896_/B _09894_/X vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09135__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__A0 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935_ _06960_/A _12280_/A _10934_/X _06681_/B vssd1 vssd1 vccd1 vccd1 _10935_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07511__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _11470_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10867_/B sky130_fd_sc_hd__xnor2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12605_ reg1_val[21] _12615_/B vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08067__A2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10797_ _11230_/A _10683_/B _11232_/A vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11071__A1 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ reg1_val[8] _12537_/B vssd1 vssd1 vccd1 vccd1 _12536_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11071__B2 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _12452_/B _12460_/B _12484_/A vssd1 vssd1 vccd1 vccd1 _12480_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06941__B _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ reg1_val[12] curr_PC[12] _12444_/S vssd1 vssd1 vccd1 vccd1 _12400_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07578__B2 _08936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__A1 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11349_ _11781_/B _11445_/B hold179/A vssd1 vssd1 vccd1 vccd1 _11349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13019_ _12765_/X _13019_/B vssd1 vssd1 vccd1 vccd1 _13020_/B sky130_fd_sc_hd__nand2b_1
X_06890_ instruction[6] instruction[5] _09148_/A vssd1 vssd1 vccd1 vccd1 _06890_/X
+ sky130_fd_sc_hd__or3_4
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _08560_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08584_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07511_ _09568_/A fanout51/X fanout49/X _09698_/A vssd1 vssd1 vccd1 vccd1 _07512_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10919__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08491_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__nand2b_1
X_07442_ _09698_/A fanout51/X fanout49/X _09885_/A vssd1 vssd1 vccd1 vccd1 _07443_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout29 _12095_/B vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__clkbuf_4
Xfanout18 _07070_/Y vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__buf_6
X_07373_ _08714_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09112_ _12499_/A reg1_val[31] _09124_/S vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09043_ _09043_/A _09043_/B vssd1 vssd1 vccd1 vccd1 _11608_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_115_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__B1 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08766__B1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11365__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ hold294/A _10080_/C _09808_/B vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__o21a_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _09876_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11522__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _09010_/B _09013_/A _09010_/A vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__o21ai_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ _08764_/B _08741_/A _08764_/A vssd1 vssd1 vccd1 vccd1 _08759_/C sky130_fd_sc_hd__mux2_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _07705_/A _07705_/B _07754_/A vssd1 vssd1 vccd1 vccd1 _07723_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08297__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ _08813_/A1 _08715_/A2 _08689_/B1 _08274_/A vssd1 vssd1 vccd1 vccd1 _08690_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _11636_/S _10716_/X _10719_/X vssd1 vssd1 vccd1 vccd1 dest_val[11] sky130_fd_sc_hd__o21ai_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ _10576_/X _10578_/Y _10581_/X _12125_/S vssd1 vssd1 vccd1 vccd1 _10582_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11053__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ reg1_val[1] curr_PC[1] _12444_/S vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08987__A_N _08871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _12253_/A _12253_/B _12253_/C vssd1 vssd1 vccd1 vccd1 _12290_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10083__A1_N _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__and2_1
X_12183_ _12302_/A _12181_/X _12182_/Y _09156_/B vssd1 vssd1 vccd1 vccd1 _12195_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10564__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _10199_/X _10201_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _11134_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07873__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _11065_/A _11065_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__or2_1
X_10016_ _11883_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09721__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__A2 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11968_/A _11968_/B vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07496__B1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ _10917_/A _10917_/B _10917_/Y _09498_/A vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ _11899_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _10850_/B _10850_/C _10850_/A vssd1 vssd1 vccd1 vccd1 _10948_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ _12519_/A _12519_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xor2_4
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout219 _13084_/A2 vssd1 vssd1 vccd1 vccd1 _13070_/A2 sky130_fd_sc_hd__buf_4
X_07991_ _11169_/A _08782_/A2 _08756_/B2 _11297_/A vssd1 vssd1 vccd1 vccd1 _07992_/B
+ sky130_fd_sc_hd__o22a_2
Xfanout208 _07847_/A vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__buf_12
XFILLER_0_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06942_ _07304_/A _07137_/A _06942_/C _06942_/D vssd1 vssd1 vccd1 vccd1 _06943_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09730_ _09730_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10858__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ instruction[20] _06887_/B vssd1 vssd1 vccd1 vccd1 _06873_/X sky130_fd_sc_hd__or2_1
X_09661_ _12125_/S _09637_/X _09642_/Y _09643_/X _06889_/Y vssd1 vssd1 vccd1 vccd1
+ _09664_/B sky130_fd_sc_hd__o221a_1
XANTENNA__10858__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _08643_/A _08643_/B vssd1 vssd1 vccd1 vccd1 _08653_/A sky130_fd_sc_hd__or2_1
X_09592_ _09592_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08543_ _08741_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout259_A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11283__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08474_ _08474_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__and2_1
XANTENNA__11283__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _10099_/A1 _10481_/A _08642_/B _12702_/A vssd1 vssd1 vccd1 vccd1 _07426_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07356_ _07916_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07361_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_18_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07287_ _07291_/A _07291_/B _07875_/A vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06581__B _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09026_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _10800_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11050__A4 _11049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09400__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09928_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout74_A _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _10126_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__xnor2_4
X_12870_ _13062_/A hold185/X vssd1 vssd1 vccd1 vccd1 _13176_/D sky130_fd_sc_hd__and2_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09467__A1 _09617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _11822_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11902_/B sky130_fd_sc_hd__and2b_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11752_ _11828_/B _11752_/B vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__nand2_1
X_10703_ hold203/A _10703_/B vssd1 vssd1 vccd1 vccd1 _10817_/B sky130_fd_sc_hd__or2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10634_ _12095_/A fanout43/X _08333_/B fanout60/X vssd1 vssd1 vccd1 vccd1 _10635_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12304_ hold301/A _12272_/Y _12304_/B1 vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__o21a_1
X_10565_ _10681_/B _10563_/X _10564_/Y vssd1 vssd1 vccd1 vccd1 _10565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12235_ hold174/A _12234_/X _09152_/Y vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09294__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12167_/B _12167_/C _12167_/A vssd1 vssd1 vccd1 vccd1 _12214_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10001__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _11155_/A _11016_/B _11159_/A vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__a21oi_1
X_12097_ _12097_/A _12097_/B vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__xor2_1
X_11048_ _09124_/S _11047_/Y _11045_/Y _11042_/X _11039_/X vssd1 vssd1 vccd1 vccd1
+ _11048_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__07108__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07181__A2 _07187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ _12773_/X _12999_/B vssd1 vssd1 vccd1 vccd1 _13000_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06666__B _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12684__A _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ _10156_/A _07210_/B vssd1 vssd1 vccd1 vccd1 _07354_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07778__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ _08205_/A _08205_/B _08183_/X vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_15_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _07142_/A _07142_/B vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08433__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _06592_/B _07068_/A _07303_/A _06801_/B vssd1 vssd1 vccd1 vccd1 _07075_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__10240__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07974_ _07974_/A _07974_/B _07975_/B vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__and3_1
X_06925_ _09495_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _06925_/X sky130_fd_sc_hd__and2_1
X_09713_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__nand2_1
X_09644_ hold247/A _13160_/Q hold189/A _12190_/B vssd1 vssd1 vccd1 vccd1 _09645_/B
+ sky130_fd_sc_hd__o31a_1
X_06856_ _12664_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _06856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06787_ _06787_/A _06787_/B vssd1 vssd1 vccd1 vccd1 _06787_/X sky130_fd_sc_hd__and2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09575_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11256__A1 _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08526_ _08734_/A _08526_/B vssd1 vssd1 vccd1 vccd1 _08577_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__inv_2
XFILLER_0_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08672__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07408_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10826__B _10826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _08388_/A _08388_/B _08388_/C vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__and3_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07339_ _07339_/A _07339_/B vssd1 vssd1 vccd1 vccd1 _07341_/B sky130_fd_sc_hd__xnor2_1
X_10350_ _10203_/S _10202_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10350_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09009_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__xor2_1
X_10281_ _10281_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10282_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10842__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _12020_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__or2_1
XANTENNA__09408__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _07832_/A _12686_/B hold151/X vssd1 vssd1 vccd1 vccd1 _13202_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12853_ hold200/A _12885_/A2 _12885_/B1 hold197/X vssd1 vssd1 vccd1 vccd1 hold198/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12784_ _12782_/X _12784_/B vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__nand2b_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08982__A _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ _11805_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11806_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11798__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11735_ _11876_/A fanout7/X fanout5/X fanout64/X vssd1 vssd1 vccd1 vccd1 _11736_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09289__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _11666_/A _11666_/B vssd1 vssd1 vccd1 vccd1 _11668_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11597_ _11757_/A _11597_/B vssd1 vssd1 vccd1 vccd1 _11600_/C sky130_fd_sc_hd__or2_1
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__xnor2_2
X_10548_ _10433_/A _10433_/B _10431_/Y vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__a21bo_1
X_13267_ instruction[6] vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
X_12218_ _12258_/D _12218_/B vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09376__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10479_ _10450_/X _10452_/X _10478_/X _10357_/X _11153_/A vssd1 vssd1 vccd1 vccd1
+ dest_val[9] sky130_fd_sc_hd__o32a_4
X_13198_ _13230_/CLK _13198_/D vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08222__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _12148_/A _12245_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06710_ reg1_val[8] _07137_/A vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07690_ _12704_/A _10009_/A _09725_/B2 _12706_/A vssd1 vssd1 vccd1 vccd1 _07691_/B
+ sky130_fd_sc_hd__o22a_1
X_06641_ reg1_val[18] _06991_/A vssd1 vssd1 vccd1 vccd1 _06641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06572_ _12278_/S _06572_/B vssd1 vssd1 vccd1 vccd1 _12264_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08892__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__A1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _11726_/A _09360_/B vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__xor2_1
X_09291_ _11134_/S _09290_/X _09166_/B vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__o21a_1
X_08311_ _08308_/A _08308_/B _08374_/A vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08242_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_46 reg2_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 reg2_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 reg2_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_68 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _08755_/A fanout41/X _08135_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08174_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout124_A _06961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ reg1_val[20] reg1_val[31] _09495_/A vssd1 vssd1 vccd1 vccd1 _07126_/C sky130_fd_sc_hd__and3_1
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07055_ _09727_/A vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09228__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__A1 _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _07981_/A _07981_/B _07956_/A vssd1 vssd1 vccd1 vccd1 _07967_/B sky130_fd_sc_hd__a21oi_2
X_06908_ reg1_val[31] _09495_/A vssd1 vssd1 vccd1 vccd1 _06908_/X sky130_fd_sc_hd__and2_1
XANTENNA__11477__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07888_ _07886_/A _07886_/B _07979_/A vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11477__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06839_ _06839_/A _06839_/B _06839_/C vssd1 vssd1 vccd1 vccd1 _06839_/X sky130_fd_sc_hd__and3_1
X_09627_ _09302_/X _09304_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _11184_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08509_ _08427_/X _08467_/Y _08466_/Y _08465_/A vssd1 vssd1 vccd1 vccd1 _08510_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _11238_/A _06641_/Y _06788_/X _11519_/X vssd1 vssd1 vccd1 vccd1 _11521_/B
+ sky130_fd_sc_hd__a31o_1
X_09489_ _09328_/A _09328_/B _09327_/A vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09842__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09842__B2 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout3_A fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _06889_/Y _11438_/X _11450_/Y _11432_/X vssd1 vssd1 vccd1 vccd1 _11451_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07605__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11491_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10403_/C sky130_fd_sc_hd__or3_1
XFILLER_0_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _13121_/A _13121_/B hold134/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__and3_1
X_10333_ _10197_/A _10194_/Y _10196_/B vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__o21a_1
XANTENNA__06959__A2 _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13052_ hold287/X _13084_/A2 _13051_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold288/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11387__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _11091_/A _07154_/X _07799_/B _06946_/X vssd1 vssd1 vccd1 vccd1 _10265_/B
+ sky130_fd_sc_hd__a22o_1
X_12003_ hold228/A _11620_/B _12067_/B _12002_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1
+ _12008_/C sky130_fd_sc_hd__a311o_1
X_10195_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07384__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ hold152/A _12662_/A _13112_/B hold110/X _13013_/A vssd1 vssd1 vccd1 vccd1
+ hold111/A sky130_fd_sc_hd__o221a_1
XANTENNA__10140__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__B2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ _13085_/A _12836_/B vssd1 vssd1 vccd1 vccd1 _13159_/D sky130_fd_sc_hd__and2_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ hold15/X hold277/A vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ hold47/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11718_ _12086_/A _11718_/B vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11649_ _11649_/A _12029_/B _11649_/C vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__and3_1
XFILLER_0_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07072__A1 _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10482__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11297__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08861_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__09482__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _07811_/A _07811_/B _07811_/C vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__or3_1
XANTENNA__08572__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08791_ _08784_/A _08784_/B _08784_/C vssd1 vssd1 vccd1 vccd1 _08792_/C sky130_fd_sc_hd__a21oi_1
X_07742_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__or2_1
XANTENNA__08324__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ _07808_/A _07808_/B _07669_/Y vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08875__A2 _08986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06624_ reg1_val[20] _07012_/B vssd1 vssd1 vccd1 vccd1 _06792_/A sky130_fd_sc_hd__nand2_1
X_09412_ _09412_/A _09412_/B vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__xnor2_1
X_09343_ hold243/A hold249/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__and3_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06555_ reg2_val[27] _06754_/B _06657_/B1 _06554_/X vssd1 vssd1 vccd1 vccd1 _07064_/B
+ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout241_A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11631__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08127__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08225_ _08272_/A _08227_/B vssd1 vssd1 vccd1 vccd1 _08225_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08156_ _08167_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__or2_1
XANTENNA__11934__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _07303_/A _07109_/A _07108_/C vssd1 vssd1 vccd1 vccd1 _08765_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__A3 _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ _08087_/A _08087_/B vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10392__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _09420_/A _07039_/B vssd1 vssd1 vccd1 vccd1 _07041_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _09048_/A _09048_/B _09048_/C _09048_/D vssd1 vssd1 vccd1 vccd1 _09049_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09512__B1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12621_ _12602_/B _12620_/X _12615_/B _07091_/D vssd1 vssd1 vccd1 vccd1 _12623_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_10882_ _10883_/B _10883_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _10884_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09421__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12552_ reg1_val[11] _12553_/B vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _12484_/A _12484_/B vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__and2_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _11504_/A _11504_/B _11504_/C vssd1 vssd1 vccd1 vccd1 _11596_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11434_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09579__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ fanout77/X fanout7/X fanout5/X fanout71/X vssd1 vssd1 vccd1 vccd1 _11366_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13104_ _13104_/A _13104_/B vssd1 vssd1 vccd1 vccd1 _13104_/Y sky130_fd_sc_hd__nand2_1
X_10316_ _11163_/A _11163_/B vssd1 vssd1 vccd1 vccd1 _10316_/Y sky130_fd_sc_hd__nor2_1
X_11296_ _11296_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__xnor2_1
X_13035_ _13035_/A _13035_/B vssd1 vssd1 vccd1 vccd1 _13035_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ _10157_/A _10157_/B _10153_/Y vssd1 vssd1 vccd1 vccd1 _10257_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07357__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _10179_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10178_/X sky130_fd_sc_hd__and2_1
XANTENNA__10361__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12676__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06955__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _13068_/A _12818_/B _12748_/X vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06674__B _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ _08010_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07045__A1 _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__B2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09961_ _09905_/A _09905_/B _09906_/Y vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__06715__A_N _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08913_/B sky130_fd_sc_hd__and2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09892_/A _09892_/B vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06849__B _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__B2 _06890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08843_/A _08843_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout289_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08774_ _08772_/A _08772_/B _08773_/X vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__a21o_1
X_07725_ _07723_/A _07723_/B _07812_/A vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07656_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07656_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06607_ reg2_val[22] _06754_/B _06539_/X _06606_/X vssd1 vssd1 vccd1 vccd1 _07028_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07587_ _07689_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__xnor2_1
X_06538_ instruction[24] _06665_/A2 _06863_/B instruction[41] _06534_/X vssd1 vssd1
+ vccd1 vccd1 _06540_/B sky130_fd_sc_hd__a221o_1
X_09326_ reg1_val[1] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__or2_1
XANTENNA__11604__A1 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _11654_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ _08606_/A2 _08715_/A2 _08689_/B1 _08642_/B vssd1 vssd1 vccd1 vccd1 _08209_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _09187_/B _09188_/B vssd1 vssd1 vccd1 vccd1 _09189_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07036__A1 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08139_ _11468_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _09145_/Y _11122_/X _11123_/Y _11149_/X _11121_/Y vssd1 vssd1 vccd1 vccd1
+ _11150_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11946__A _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ fanout77/X fanout36/X fanout34/X fanout74/X vssd1 vssd1 vccd1 vccd1 _10102_/B
+ sky130_fd_sc_hd__o22a_1
X_11081_ fanout76/X fanout14/X fanout52/X _11663_/A vssd1 vssd1 vccd1 vccd1 _11082_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10850__A _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _10032_/A _10032_/B vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13243_/CLK sky130_fd_sc_hd__clkbuf_8
X_11983_ _11983_/A _11983_/B _11983_/C vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__and3_1
XANTENNA__07511__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ _10933_/A _09141_/Y _10933_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _10934_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ _11876_/A fanout41/X _08135_/B _11950_/A vssd1 vssd1 vccd1 vccd1 _10866_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ reg1_val[21] _12615_/B vssd1 vssd1 vccd1 vccd1 _12604_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _12534_/A _12531_/Y _12533_/B vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10796_ _11014_/A _10796_/B vssd1 vssd1 vccd1 vccd1 _11230_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09297__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11071__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12466_ _12464_/X _12466_/B vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12397_ _12403_/B _12397_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
XANTENNA__06941__C _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11417_ _11329_/A _11326_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__a21o_1
X_11348_ hold184/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__or2_1
XANTENNA__07578__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11279_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10760__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _13103_/A hold262/X vssd1 vssd1 vccd1 vccd1 _13234_/D sky130_fd_sc_hd__and2_1
XANTENNA__08230__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07510_ _07501_/A _07501_/B _07536_/B vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_77_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ _08490_/A _08490_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__xor2_1
X_07441_ _12085_/A _07441_/B vssd1 vssd1 vccd1 vccd1 _07444_/A sky130_fd_sc_hd__xnor2_1
Xfanout19 _12223_/A vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__buf_4
X_07372_ _06977_/A _12704_/A _12706_/A _06985_/A vssd1 vssd1 vccd1 vccd1 _07373_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09996__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ _09110_/X _09103_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09111_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09042_ _09045_/B _09045_/C vssd1 vssd1 vccd1 vccd1 _11608_/B sky130_fd_sc_hd__or2_1
XANTENNA__07018__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__B2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__B1 _07156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ hold222/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09944_/Y sky130_fd_sc_hd__xnor2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__B1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__xnor2_1
X_08826_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__nor2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _08801_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__xnor2_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07708_ _07753_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__and2_1
XFILLER_0_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08688_ _08688_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__xnor2_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07639_/A _07639_/B _07639_/C vssd1 vssd1 vccd1 vccd1 _07640_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10650_/Y sky130_fd_sc_hd__nand2_1
X_09309_ _09097_/X _09124_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10581_ _09951_/Y _10580_/Y _11135_/S vssd1 vssd1 vccd1 vccd1 _10581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10845__A _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12320_ _12326_/A _12320_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
X_12251_ _12288_/A _12251_/B vssd1 vssd1 vccd1 vccd1 _12253_/C sky130_fd_sc_hd__or2_1
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11202_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__nor2_1
X_12182_ _12302_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10564__A1 _10681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__S _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11133_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/Y sky130_fd_sc_hd__xnor2_1
X_11064_ _11065_/A _11065_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__nand2_1
X_10015_ _12141_/A _10370_/A _07763_/B fanout45/X vssd1 vssd1 vccd1 vccd1 _10016_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07193__B1 _07069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11966_ _11966_/A _11966_/B vssd1 vssd1 vccd1 vccd1 _11968_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07496__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _10917_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10917_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11897_ _11897_/A _11897_/B vssd1 vssd1 vccd1 vccd1 _11899_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ _10847_/A _10847_/B _11271_/A vssd1 vssd1 vccd1 vccd1 _10850_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12241__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _10667_/A _10667_/B _10665_/Y vssd1 vssd1 vccd1 vccd1 _10781_/B sky130_fd_sc_hd__a21bo_1
X_12518_ _12516_/Y _12518_/B vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ _12454_/C _12449_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 _08688_/A vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__buf_12
X_07990_ _08814_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06941_ _06941_/A _06963_/A _06960_/A _07278_/A vssd1 vssd1 vccd1 vccd1 _06942_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_0_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12701__C1 _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _11238_/A _09637_/X _09659_/Y _09136_/B vssd1 vssd1 vccd1 vccd1 _09660_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09173__A1 _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06872_ instruction[12] _06850_/Y _06871_/X _12498_/C vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_08611_ _08814_/A _08611_/B vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10858__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ _09592_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__and2b_1
X_08542_ _08740_/A2 _08735_/A2 _08735_/B1 _08755_/B vssd1 vssd1 vccd1 vccd1 _08543_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07304__A _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11283__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07424_ _07420_/A _07420_/B _07504_/A vssd1 vssd1 vccd1 vccd1 _07434_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout154_A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07355_ fanout51/X _09885_/A _09880_/B2 fanout49/X vssd1 vssd1 vccd1 vccd1 _07356_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06862__B _06862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07286_ _11468_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08135__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09025_ _09025_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12880__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__buf_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _09801_/A _09798_/Y _09801_/C vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__o21a_1
XANTENNA_fanout67_A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _10009_/A fanout9/X fanout3/X _07015_/Y vssd1 vssd1 vccd1 vccd1 _09859_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09079_/X _09094_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__mux2_1
X_08809_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__nor2_1
X_11820_ _11902_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__nor2_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__nand2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _11696_/A _10700_/X _10701_/X _12303_/A vssd1 vssd1 vccd1 vccd1 _10715_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11682_ _12110_/A _11834_/A _11834_/B _09621_/A vssd1 vssd1 vccd1 vccd1 _11683_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10633_ _10767_/B _10633_/B vssd1 vssd1 vccd1 vccd1 _10656_/A sky130_fd_sc_hd__or2_1
XFILLER_0_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _10681_/B _10563_/X _09061_/X vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ _12303_/A _12303_/B _12303_/C vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__or3_1
XFILLER_0_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _10494_/B _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__nand2b_1
X_12234_ hold233/A _12275_/C _12190_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _12165_/A vssd1 vssd1 vccd1 vccd1 _12167_/C sky130_fd_sc_hd__inv_2
X_11116_ _11159_/B _11160_/A vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12096_ _12094_/A _12094_/Y _12096_/S vssd1 vssd1 vccd1 vccd1 _12097_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07166__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _11346_/B vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07108__B _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12998_ _13013_/A _12998_/B vssd1 vssd1 vccd1 vccd1 _13230_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ _11949_/A _11949_/B vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10473__B1 _10470_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__A _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ _07916_/A _07140_/B vssd1 vssd1 vccd1 vccd1 _07142_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07071_ _08384_/B _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _07078_/B sky130_fd_sc_hd__and3_1
XANTENNA__12201__C_N _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__B1 _10321_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__B1 _07156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07973_ _07975_/B _07975_/A vssd1 vssd1 vccd1 vccd1 _07973_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09713_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06924_ _10850_/A _10761_/A _06921_/X vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout271_A hold177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06855_ _06754_/B _06532_/X _09153_/A instruction[4] _06852_/Y vssd1 vssd1 vccd1
+ vccd1 _12664_/B sky130_fd_sc_hd__a221o_1
X_09643_ _09638_/X _09640_/X _09641_/Y _11696_/A vssd1 vssd1 vccd1 vccd1 _09643_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _09574_/A _09574_/B vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__xnor2_1
X_06786_ _06785_/A _06785_/B _11339_/A vssd1 vssd1 vccd1 vccd1 _06787_/B sky130_fd_sc_hd__o21bai_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08219_/B _09180_/B2 _10506_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08526_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11256__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08456_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__xnor2_1
X_07407_ _07407_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _09420_/A _08387_/B _08387_/C vssd1 vssd1 vccd1 vccd1 _08388_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10395__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _07338_/A vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__inv_2
XANTENNA__06592__B _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07269_ _12668_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _07635_/S sky130_fd_sc_hd__or2_1
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09019_/A sky130_fd_sc_hd__xnor2_1
X_10280_ _10281_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11954__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ hold150/X _12665_/A _13112_/B hold136/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold151/A sky130_fd_sc_hd__o221a_1
X_12852_ _13071_/A hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__and2_1
X_12783_ hold257/X hold45/X vssd1 vssd1 vccd1 vccd1 _12784_/B sky130_fd_sc_hd__nand2b_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11803_ _11803_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10455__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11657_/A _11657_/B _11653_/X vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__a21o_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _11665_/A _11665_/B vssd1 vssd1 vccd1 vccd1 _11666_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09860__A2 _07070_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10616_ _10616_/A _10616_/B vssd1 vssd1 vccd1 vccd1 _10617_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11596_ _11596_/A _11596_/B _11596_/C vssd1 vssd1 vccd1 vccd1 _11597_/B sky130_fd_sc_hd__and3_1
XFILLER_0_122_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10547_ _10547_/A _10547_/B vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__xnor2_1
X_10478_ _09156_/B _10464_/X _10477_/X _10456_/X vssd1 vssd1 vccd1 vccd1 _10478_/X
+ sky130_fd_sc_hd__a211o_2
X_13266_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
X_12217_ _12258_/D _12218_/B vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__or2_1
XANTENNA__09376__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ _13230_/CLK _13197_/D vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07387__B1 _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _12148_/A _12245_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__or3_1
XANTENNA__07139__B1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ curr_PC[25] curr_PC[26] _12079_/C vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__and3_1
XANTENNA__12132__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__A_N _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ reg2_val[18] _06700_/B _06657_/B1 _06638_/X vssd1 vssd1 vccd1 vccd1 _06980_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06571_ reg1_val[30] _07255_/A vssd1 vssd1 vccd1 vccd1 _06572_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _10073_/S _09289_/X _09164_/B vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _08373_/B _08310_/B vssd1 vssd1 vccd1 vccd1 _08374_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 instruction[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06665__A2 _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ _08241_/A _08241_/B _08241_/C vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__or3_1
XANTENNA_47 reg2_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 reg2_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_25 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_58 reg2_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08172_ _11072_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07301__B _07301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _07123_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07123_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ _07056_/B _07056_/A _08688_/A vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__B2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _07956_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__nor2_1
X_06907_ _06907_/A vssd1 vssd1 vccd1 vccd1 _06907_/Y sky130_fd_sc_hd__inv_2
X_07887_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__or2_1
XANTENNA__11477__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ _06838_/A _06838_/B vssd1 vssd1 vccd1 vccd1 _06839_/C sky130_fd_sc_hd__nor2_1
X_09626_ _09301_/X _09313_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09626_/X sky130_fd_sc_hd__mux2_1
X_06769_ _09785_/B _09785_/C _06834_/A vssd1 vssd1 vccd1 vccd1 _09924_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ fanout78/X fanout77/X fanout74/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _09558_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _09481_/X _09487_/X _10809_/A vssd1 vssd1 vccd1 vccd1 _09488_/X sky130_fd_sc_hd__mux2_2
X_08508_ _08512_/A _08512_/B _08507_/A vssd1 vssd1 vccd1 vccd1 _08553_/A sky130_fd_sc_hd__a21oi_1
X_08439_ _09564_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09842__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12729__A2 _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _11450_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11450_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07605__A1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__B2 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11656_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10403_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10853__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13120_ hold161/A hold164/A hold100/X hold133/X vssd1 vssd1 vccd1 vccd1 hold134/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _10331_/A _10331_/B _10331_/Y _09498_/A vssd1 vssd1 vccd1 vccd1 _10332_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09419__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ hold298/A _13050_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _11620_/B _12067_/B hold228/A vssd1 vssd1 vccd1 vccd1 _12002_/Y sky130_fd_sc_hd__a21oi_1
X_10263_ _10263_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__xor2_1
X_10194_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12499__B _12499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12904_ _07039_/B _12664_/Y hold153/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__a21boi_1
XANTENNA__06928__D _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__A2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ hold189/X _13084_/A2 fanout2/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 _12836_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06895__A2 _06890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ hold261/X hold70/X vssd1 vssd1 vccd1 vccd1 _13019_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__B2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _08384_/A _12731_/A2 hold63/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13141_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11717_ _12094_/A fanout15/X _07513_/B _07070_/Y vssd1 vssd1 vccd1 vccd1 _11718_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _11723_/B _11648_/B vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11579_ _11579_/A _11579_/B _11577_/Y vssd1 vssd1 vccd1 vccd1 _11580_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08233__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13249_ _13250_/CLK _13249_/D vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09349__B2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ _07810_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _07813_/B sky130_fd_sc_hd__xnor2_1
X_08790_ _08790_/A vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__inv_2
XANTENNA__08572__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _07739_/A _07739_/B _07740_/X vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07808_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09521__B2 _07156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06623_ reg2_val[20] _06700_/B _06657_/B1 _06621_/X vssd1 vssd1 vccd1 vccd1 _06982_/A
+ sky130_fd_sc_hd__a22o_2
X_09411_ _09412_/B vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__inv_2
X_09342_ hold33/A _09495_/A vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__and2_1
XANTENNA__12959__A2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06554_ _06613_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _06554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09273_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08224_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08227_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11919__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ _08204_/A _08204_/B _08145_/X vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ _07106_/A _07106_/B vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ _08734_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ reg1_val[2] _07037_/B vssd1 vssd1 vccd1 vccd1 _07039_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08988_ _08988_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__xnor2_2
X_07939_ _08535_/A _07939_/B vssd1 vssd1 vccd1 vccd1 _07942_/B sky130_fd_sc_hd__xnor2_1
X_10950_ _10950_/A _10950_/B _10950_/C vssd1 vssd1 vccd1 vccd1 _10951_/B sky130_fd_sc_hd__and3_1
X_09609_ _09609_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__xor2_1
X_10881_ _10747_/A _10747_/B _10743_/X vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ _12620_/A _12620_/B _12620_/C _12620_/D vssd1 vssd1 vccd1 vccd1 _12620_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12556_/B _12551_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
X_12482_ reg1_val[25] curr_PC[25] _12495_/S vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11596_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11504_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11433_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11433_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09579__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11386__B2 _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11364_ _12089_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__xnor2_1
X_13103_ _13103_/A hold252/X vssd1 vssd1 vccd1 vccd1 _13252_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _09773_/Y _11163_/B _10311_/X _10314_/Y vssd1 vssd1 vccd1 vccd1 _10315_/X
+ sky130_fd_sc_hd__o211a_1
X_11295_ _11462_/A fanout7/X fanout5/X _11295_/B2 vssd1 vssd1 vccd1 vccd1 _11296_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13034_ _12759_/X _13034_/B vssd1 vssd1 vccd1 vccd1 _13035_/B sky130_fd_sc_hd__nand2b_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _10421_/B _10246_/B vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12303__A _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _10177_/A _10177_/B vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10361__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06955__B _06961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ _12748_/X _12818_/B vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__nand2b_1
X_12749_ hold13/X hold263/X vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12692__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10493__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__A2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09960_ _09910_/A _09910_/B _09908_/X vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__a21oi_4
X_08911_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__nor2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08842_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07307__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08784_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08773_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout184_A _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ _07811_/A _07811_/B _07811_/C vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07657_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09522__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _06613_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _06606_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07586_ _06977_/A fanout68/X fanout65/X _06985_/A vssd1 vssd1 vccd1 vccd1 _07587_/B
+ sky130_fd_sc_hd__o22a_1
X_06537_ instruction[41] _06863_/B _06534_/X vssd1 vssd1 vccd1 vccd1 _06537_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ reg1_val[1] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ fanout92/X _11564_/A fanout38/X _10876_/A1 vssd1 vssd1 vccd1 vccd1 _09257_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09187_ _09188_/B _09187_/B vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08782_/B2 fanout37/X _08233_/B _08813_/B1 vssd1 vssd1 vccd1 vccd1 _08139_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12317__A0 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _10957_/A _08782_/A2 _08756_/B2 fanout81/X vssd1 vssd1 vccd1 vccd1 _08070_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout97_A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _11656_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__xnor2_1
X_11080_ _11296_/A _11080_/B vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _10029_/Y _10031_/B vssd1 vssd1 vccd1 vccd1 _10032_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11982_ _11983_/A _11983_/C _11983_/B vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__a21oi_1
X_10933_ _10933_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _10933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09151__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ _10864_/A _10864_/B vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__nor2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12603_/A _12603_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
X_10795_ _10319_/B _11157_/A _10793_/X _10792_/X _10677_/B vssd1 vssd1 vccd1 vccd1
+ _10796_/B sky130_fd_sc_hd__a2111o_4
XANTENNA__11056__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ _12496_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12466_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12397_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06941__D _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ _12125_/S _11345_/Y _11346_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__and2_1
X_13017_ hold261/X _06858_/B _13016_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold262/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08230__B _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _11184_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__xnor2_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06685__B _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11295__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ _12668_/A fanout15/X _07513_/B _09237_/A vssd1 vssd1 vccd1 vccd1 _07441_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09061__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07371_ _10126_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _09106_/X _09109_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _09041_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _09045_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07018__A2 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ hold239/A _10077_/C _10208_/B vssd1 vssd1 vccd1 vccd1 _09944_/B sky130_fd_sc_hd__o21ai_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09874_/Y sky130_fd_sc_hd__nor2_1
X_08825_ _09564_/A _08820_/X _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09012_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ _08782_/A2 _08782_/B2 _08813_/B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08757_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _11183_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__xnor2_1
X_08687_ _08782_/A2 _08737_/A2 _08733_/B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08688_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10398__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13027__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07639_/A _07639_/B _07639_/C vssd1 vssd1 vccd1 vccd1 _07640_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07569_ _07569_/A _07569_/B _07569_/C vssd1 vssd1 vccd1 vccd1 _07570_/B sky130_fd_sc_hd__or3_1
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _09300_/X _09307_/X _10924_/S vssd1 vssd1 vccd1 vccd1 _09308_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10580_ _10580_/A vssd1 vssd1 vccd1 vccd1 _10580_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10845__B _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _09568_/A fanout8/X _09428_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _09240_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _12250_/A _12250_/B _12250_/C vssd1 vssd1 vccd1 vccd1 _12251_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09954__A1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ reg1_val[28] _12226_/C vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__xor2_1
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ _11032_/A _11032_/B _11030_/B vssd1 vssd1 vccd1 vccd1 _11133_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10861__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__B _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ _11063_/A _11063_/B vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__xor2_1
X_10014_ _10014_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07193__B2 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__A1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__B _08985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11965_ _11965_/A _11965_/B vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07496__A2 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916_ _11238_/A _10915_/X _10914_/X vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__o21ba_1
X_11896_ _11896_/A _11896_/B vssd1 vssd1 vccd1 vccd1 _11897_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ _10847_/A _10847_/B _11271_/A vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08445__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778_ _10778_/A _10778_/B vssd1 vssd1 vccd1 vccd1 _10781_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ reg1_val[4] _12517_/B vssd1 vssd1 vccd1 vccd1 _12518_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ _12455_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12449_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11867__A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12542_/B _12379_/B vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ _06940_/A vssd1 vssd1 vccd1 vccd1 _06940_/Y sky130_fd_sc_hd__inv_2
X_06871_ instruction[19] _06887_/B vssd1 vssd1 vccd1 vccd1 _06871_/X sky130_fd_sc_hd__or2_1
XANTENNA__09173__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__C1 _10711_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _08813_/A1 _09180_/B2 _10506_/A _08274_/A vssd1 vssd1 vccd1 vccd1 _08611_/B
+ sky130_fd_sc_hd__o22a_1
X_09590_ _09590_/A _09590_/B vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11268__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ _08714_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08472_ _09041_/A _09000_/A vssd1 vssd1 vccd1 vccd1 _08472_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08133__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ _07503_/A _07503_/B vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__and2_1
XFILLER_0_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A _07122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _07354_/A _07354_/B vssd1 vssd1 vccd1 vccd1 _07366_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _11468_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08135__B _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _09004_/A _09004_/B _08727_/A vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__a21oi_1
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A1 _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10681__A _10681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 hold302/X vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__buf_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _09926_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09926_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07990__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__xor2_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _06834_/A _09786_/X _09787_/Y vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__o21a_1
X_08808_ _09423_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _08812_/B sky130_fd_sc_hd__xnor2_1
X_08739_ _08763_/A _08763_/B _08738_/X vssd1 vssd1 vccd1 vccd1 _08744_/A sky130_fd_sc_hd__or3b_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11750_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__or2_1
XANTENNA__08124__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10696_/X _10697_/Y _12125_/S vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09872__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__xor2_1
X_10632_ _10632_/A _10632_/B vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__nor2_1
X_10563_ _10681_/A _10449_/C _10449_/A vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _12302_/A _12302_/B _12302_/C vssd1 vssd1 vccd1 vccd1 _12303_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10494_ _10495_/B _10494_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__nand2b_1
X_12233_ hold251/A _12231_/X _12232_/Y vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07938__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _12042_/X _12161_/Y _12163_/Y vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08061__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ _12095_/A _12095_/B _12030_/A vssd1 vssd1 vccd1 vccd1 _12096_/S sky130_fd_sc_hd__or3b_1
X_11115_ _11114_/A _11114_/B _11114_/C vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__a21o_1
X_11046_ _10809_/A _09322_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__B2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__A1 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__C _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ hold300/X _12663_/B _12996_/X _12664_/A vssd1 vssd1 vccd1 vccd1 _12998_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11948_ _11948_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__and2_1
XANTENNA__10473__B2 _10471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ _11879_/A _11879_/B _11879_/C vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__and3_1
XFILLER_0_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07140__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07070_ _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _07070_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11725__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__B2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07972_ _07972_/A _07972_/B vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__xor2_2
X_09711_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__or2_1
X_06923_ _10850_/A _10761_/A _06921_/X vssd1 vssd1 vccd1 vccd1 _06923_/Y sky130_fd_sc_hd__a21oi_1
X_06854_ _06754_/B _06532_/X _09153_/A instruction[4] _06852_/Y vssd1 vssd1 vccd1
+ vccd1 _12665_/B sky130_fd_sc_hd__a221oi_2
XFILLER_0_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09642_ _09640_/X _09641_/Y _09638_/X vssd1 vssd1 vccd1 vccd1 _09642_/Y sky130_fd_sc_hd__a21oi_1
X_06785_ _06785_/A _06785_/B vssd1 vssd1 vccd1 vccd1 _06785_/Y sky130_fd_sc_hd__nor2_1
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08524_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06873__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _08464_/A _08464_/B _08464_/C vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__o21ai_1
X_07406_ _07364_/A _07364_/B _07364_/C vssd1 vssd1 vccd1 vccd1 _07407_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06683__A3 _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08386_ _08387_/B _08387_/C _09420_/A vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07050__A _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ _07337_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07268_/A _12245_/A vssd1 vssd1 vccd1 vccd1 fanout8/A sky130_fd_sc_hd__nand2_2
X_07199_ _07377_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07335_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ _09007_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _10187_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12677__C1 _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__xor2_2
X_12920_ _06996_/B _12686_/B hold158/X vssd1 vssd1 vccd1 vccd1 _13201_/D sky130_fd_sc_hd__a21boi_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ hold241/A _12885_/A2 _12885_/B1 hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11802_ _11879_/B _11802_/B vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__nand2_1
X_12782_ hold45/X hold257/X vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__and2b_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11650_/A _11650_/B _11660_/A vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__a21bo_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11664_ _11665_/A _11665_/B vssd1 vssd1 vccd1 vccd1 _11664_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08056__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10615_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10616_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ _11596_/A _11596_/B _11596_/C vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ _10546_/A _10546_/B vssd1 vssd1 vccd1 vccd1 _10547_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ instruction[15] vssd1 vssd1 vccd1 vccd1 loadstore_dest[4] sky130_fd_sc_hd__buf_12
X_10477_ _09135_/Y _10463_/X _10476_/Y _09064_/Y _10474_/Y vssd1 vssd1 vccd1 vccd1
+ _10477_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _12258_/A _12258_/B _12258_/C _12112_/A vssd1 vssd1 vccd1 vccd1 _12218_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09376__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _13230_/CLK _13196_/D vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07387__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _12208_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ curr_PC[25] _12079_/C curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12078_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11029_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12683__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06974__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06570_ reg1_val[30] _07255_/A vssd1 vssd1 vccd1 vccd1 _12278_/S sky130_fd_sc_hd__and2_1
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08241_/C sky130_fd_sc_hd__and2_1
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 instruction[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 reg2_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 reg2_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08171_ _08733_/B1 fanout43/X _08333_/B _08735_/A2 vssd1 vssd1 vccd1 vccd1 _08172_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_59 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ _07123_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07122_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_55_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07053_ _09423_/A _07053_/B vssd1 vssd1 vccd1 vccd1 _07056_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11174__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07955_ _07955_/A _08027_/A _07955_/C vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__and3_1
XANTENNA__09525__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ instruction[6] instruction[5] _12280_/A vssd1 vssd1 vccd1 vccd1 _06907_/A
+ sky130_fd_sc_hd__a21oi_4
XANTENNA__10134__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09625_ _09623_/X _09624_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__mux2_1
X_07886_ _07886_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10685__A1 _11230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ _06837_/A _11767_/A _11689_/A _06837_/D vssd1 vssd1 vccd1 vccd1 _06838_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__11882__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ _09651_/B _09651_/C _06834_/B vssd1 vssd1 vccd1 vccd1 _09785_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09827__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__xor2_1
X_06699_ _10586_/S _06699_/B vssd1 vssd1 vccd1 vccd1 _10570_/A sky130_fd_sc_hd__nand2_1
X_09487_ _09484_/X _09486_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09487_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08507_ _08507_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07302__A1 _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ _08815_/B fanout93/X _10647_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08439_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _08369_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _08370_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07066__B1 _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _12094_/A fanout50/X _07988_/B _12148_/A vssd1 vssd1 vccd1 vccd1 _11381_/B
+ sky130_fd_sc_hd__o22a_1
X_10400_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10402_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _13050_/A _13050_/B vssd1 vssd1 vccd1 vccd1 _13050_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _10263_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__nor2_1
X_12001_ hold231/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12067_/B sky130_fd_sc_hd__or2_1
XANTENNA__08566__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _10067_/A _10064_/Y _10066_/B vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__o21a_1
X_12903_ hold124/X _12662_/A _13112_/B hold152/X _13013_/A vssd1 vssd1 vccd1 vccd1
+ hold153/A sky130_fd_sc_hd__o221a_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _13109_/A _13109_/B _13109_/C vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__o21bai_1
XANTENNA__09818__B1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ hold70/X hold261/X vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__and2b_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11883_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10979__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ hold62/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__or2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11647_ _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12050__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11578_ _11579_/A _11579_/B _11577_/Y vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10529_ _10529_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10600__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08233__B _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13248_ _13250_/CLK _13248_/D vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _13185_/CLK hold170/X vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06969__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _07821_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_74_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07532__A1 _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09521__A2 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06622_ reg2_val[20] _06700_/B _06657_/B1 _06621_/X vssd1 vssd1 vccd1 vccd1 _07012_/B
+ sky130_fd_sc_hd__a22oi_4
X_09410_ _10529_/A _09410_/B vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__xnor2_2
X_06553_ instruction[37] _06637_/B vssd1 vssd1 vccd1 vccd1 _12559_/B sky130_fd_sc_hd__and2_4
X_09341_ _06759_/Y _09138_/X _11625_/B _06761_/A vssd1 vssd1 vccd1 vccd1 _09341_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09272_ _08960_/A _08960_/B _08958_/X vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08223_ _08223_/A _08223_/B _08223_/C vssd1 vssd1 vccd1 vccd1 _08272_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10954__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _08154_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08204_/B sky130_fd_sc_hd__xnor2_4
X_07105_ _11955_/A _07112_/B _12085_/A vssd1 vssd1 vccd1 vccd1 _07106_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08085_ fanout81/X _08219_/B _08815_/B _11169_/A vssd1 vssd1 vccd1 vccd1 _08086_/B
+ sky130_fd_sc_hd__o22a_1
X_07036_ _12499_/A reg1_val[1] _07050_/A vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07220__B1 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06598__B _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _08871_/Y _08987_/B vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__nand2b_1
X_07938_ fanout83/X _09180_/B2 _10506_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _07939_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07869_ fanout79/X _12684_/A _12686_/A _06961_/Y vssd1 vssd1 vccd1 vccd1 _07870_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _09609_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09608_/X sky130_fd_sc_hd__and2_1
X_10880_ _10880_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout42_A fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ _06977_/A fanout63/X fanout60/X _06985_/A vssd1 vssd1 vccd1 vccd1 _09540_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ _12550_/A _12550_/B _12550_/C vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12481_ _12481_/A _12481_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XANTENNA__10830__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ _11501_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11432_ _11431_/A _11431_/B _11431_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11432_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09579__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__B1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11386__A2 _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ hold251/X _06858_/B _13101_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold252/A
+ sky130_fd_sc_hd__a22o_1
X_11363_ _11663_/A fanout11/X fanout44/X _11739_/A vssd1 vssd1 vccd1 vccd1 _11364_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__nor2_1
X_10314_ _10314_/A vssd1 vssd1 vccd1 vccd1 _10314_/Y sky130_fd_sc_hd__inv_2
X_13033_ _13080_/A hold274/X vssd1 vssd1 vccd1 vccd1 _13237_/D sky130_fd_sc_hd__and2_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10246_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10176_ _10177_/B _10177_/A vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout190 _06971_/X vssd1 vssd1 vccd1 vccd1 _08698_/A sky130_fd_sc_hd__buf_8
XFILLER_0_89_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ hold269/X hold21/X vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12748_ hold21/X hold269/X vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ _07147_/Y _12731_/A2 hold52/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13132_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _10126_/A _08910_/B vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__xnor2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09890_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08841_/A _08841_/B _08841_/C vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__and3_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08772_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__xor2_2
X_07723_ _07723_/A _07723_/B vssd1 vssd1 vccd1 vccd1 _07811_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11837__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _07011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _07655_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07654_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06605_ instruction[32] _06637_/B vssd1 vssd1 vccd1 vccd1 _12532_/B sky130_fd_sc_hd__and2_4
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07585_ _07585_/A _07585_/B vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06536_ instruction[41] _06863_/B _06534_/X vssd1 vssd1 vccd1 vccd1 _06727_/B sky130_fd_sc_hd__a21o_1
X_09324_ _09324_/A vssd1 vssd1 vccd1 vccd1 _09324_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _09255_/A _09255_/B vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10684__A _11230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _08249_/A _08249_/B vssd1 vssd1 vccd1 vccd1 _08206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ _11794_/A _09186_/B vssd1 vssd1 vccd1 vccd1 _09187_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ _08137_/A _08137_/B vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ _08734_/A _08068_/B vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07019_ _08698_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07021_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10030_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__nand2_1
X_11981_ _11980_/A _11980_/B _09061_/X vssd1 vssd1 vccd1 vccd1 _11981_/Y sky130_fd_sc_hd__a21oi_1
X_10932_ hold297/A _12000_/A2 _11037_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _10932_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10859__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07233__A _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10863_ _10863_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ _12620_/A _12602_/B _12602_/C vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__and3_2
X_10794_ _10794_/A _10794_/B _10794_/C vssd1 vssd1 vccd1 vccd1 _11157_/A sky130_fd_sc_hd__and3_1
XANTENNA__11056__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12533_ _12531_/Y _12533_/B vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12464_ _12496_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__and2_1
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12395_ _12396_/A _12396_/B _12396_/C vssd1 vssd1 vccd1 vccd1 _12403_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _11509_/A vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10567__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _12125_/S _11346_/B vssd1 vssd1 vccd1 vccd1 _11346_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ hold277/A _13015_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09185__B1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11277_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06538__A2 _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10852_/B2 fanout63/X fanout55/X fanout78/X vssd1 vssd1 vccd1 vccd1 _10229_/B
+ sky130_fd_sc_hd__o22a_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10159_ _10159_/A _10159_/B _10157_/Y vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09342__B _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11295__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11295__B2 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ fanout77/X _10009_/A _09725_/B2 _12710_/A vssd1 vssd1 vccd1 vccd1 _07371_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09660__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ _09000_/A _09000_/B _08556_/B vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10009__A _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09942_ _12302_/A _09940_/X _09941_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _09942_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout294_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _10529_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__xnor2_1
X_08824_ _09420_/A _09015_/A vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__nor2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10730__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ _08755_/A _08755_/B vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__or2_1
X_07706_ _09880_/B2 fanout37/X fanout34/X _10117_/A vssd1 vssd1 vccd1 vccd1 _07707_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07053__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ _08686_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _08696_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13027__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07639_/C sky130_fd_sc_hd__xnor2_1
X_07568_ _07569_/A _07569_/B _07569_/C vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07988__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ _09306_/X _09303_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__mux2_1
X_06519_ _09495_/A vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__inv_2
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07499_ _07495_/A _07495_/B _07700_/A vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ _08933_/A _08933_/B _08931_/X vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _09130_/Y _09330_/A _12302_/B _09293_/A _09155_/Y vssd1 vssd1 vccd1 vccd1
+ _09169_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _12124_/A _12121_/Y _12123_/B vssd1 vssd1 vccd1 vccd1 _12226_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ _11199_/B _11200_/B vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__and2b_1
X_11131_ _11129_/Y _11131_/B vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_102_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11063_/A _11063_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__nand2_1
X_10013_ _10115_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11964_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _11965_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10915_ _06831_/D _10803_/B _10823_/A vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__o21a_1
X_11895_ _11895_/A _11895_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__nor3_1
X_10846_ _07075_/A _07075_/B _07239_/A vssd1 vssd1 vccd1 vccd1 _10847_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ _10777_/A _10777_/B vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__and2_1
XFILLER_0_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ reg1_val[4] _12517_/B vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _12455_/C _12447_/B vssd1 vssd1 vccd1 vccd1 _12454_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ _12542_/B _12379_/B vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11329_/A _11329_/B _11418_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06870_ instruction[11] _06850_/Y _06869_/X _12498_/C vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12701__A1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08905__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__B1 _10710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__A _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08133__A1 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _08670_/A2 _08737_/A2 _08733_/B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08541_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11268__A1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__B2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08471_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08133__B2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07422_ _11183_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07503_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07601__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07353_ _07349_/A _07349_/B _07439_/A vssd1 vssd1 vccd1 vccd1 _07368_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07284_ reg1_val[20] _07284_/B vssd1 vssd1 vccd1 vccd1 _07286_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _09023_/A _09023_/B vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__or2_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09397__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__12940__A1 _07286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10681__B _10681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _12263_/S _09923_/Y _09924_/X vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__a21bo_1
X_09856_ _09854_/Y _09856_/B vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__nand2b_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _09313_/S _08219_/B _09222_/B2 _09237_/A vssd1 vssd1 vccd1 vccd1 _08808_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _06999_/A _06999_/B vssd1 vssd1 vccd1 vccd1 _06999_/Y sky130_fd_sc_hd__nand2_2
X_09787_ _06834_/A _09786_/X _09498_/A vssd1 vssd1 vccd1 vccd1 _09787_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08124__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _08801_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08738_/X sky130_fd_sc_hd__xor2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__xor2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _09814_/Y _10699_/Y _11135_/S vssd1 vssd1 vccd1 vccd1 _10700_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09872__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11680_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11834_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08607__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10631_ _10632_/A _10632_/B vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _10794_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__xor2_4
X_12301_ _12302_/A _12302_/C _12302_/B vssd1 vssd1 vccd1 vccd1 _12303_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ hold251/A _12231_/X _09150_/Y vssd1 vssd1 vccd1 vccd1 _12232_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ _11799_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08342__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12107_/A _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12163_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__07938__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__B1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12094_ _12094_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12094_/Y sky130_fd_sc_hd__nor2_1
X_11114_ _11114_/A _11114_/B _11114_/C vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__nand3_1
X_11045_ _06963_/A _12280_/A _11044_/X _06675_/B vssd1 vssd1 vccd1 vccd1 _11045_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09560__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ hold289/X _12995_/Y hold246/X vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11947_ _11948_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _11949_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07124__C _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07874__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _11879_/A _11879_/B _11879_/C vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__a21oi_1
X_10829_ _09330_/A _10810_/Y _10828_/Y _09293_/A _10826_/X vssd1 vssd1 vccd1 vccd1
+ _10829_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_55_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12922__A1 _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11489__A1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06922_ _10607_/A _06922_/B vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__and2_1
X_09710_ _10529_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09551__B1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__nand2_1
X_06853_ instruction[5] instruction[6] vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__nand2b_4
X_06784_ _11238_/B _11238_/C _11240_/A vssd1 vssd1 vccd1 vccd1 _06785_/B sky130_fd_sc_hd__a21boi_1
X_09572_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09572_/Y sky130_fd_sc_hd__nor2_1
X_08523_ _08801_/A _08523_/B vssd1 vssd1 vccd1 vccd1 _08528_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout257_A _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__A _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07865__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08464_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__xnor2_1
X_08385_ _06938_/A _06938_/B _06828_/A vssd1 vssd1 vccd1 vccd1 _08387_/C sky130_fd_sc_hd__a21o_1
X_07336_ _07336_/A _07336_/B vssd1 vssd1 vccd1 vccd1 _07343_/A sky130_fd_sc_hd__or2_1
XANTENNA__07617__B1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07267_ _12142_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__nand2_1
X_09006_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__xor2_1
X_07198_ _07198_/A _07198_/B vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08345__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09908_/X sky130_fd_sc_hd__and2_1
XANTENNA__08345__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _09677_/Y _09680_/B _09685_/A vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__a21o_2
X_12850_ _13071_/A hold242/X vssd1 vssd1 vccd1 vccd1 _13166_/D sky130_fd_sc_hd__and2_1
XFILLER_0_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11801_ _11801_/A _11801_/B vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__nand2_1
X_12781_ _12779_/X _12781_/B vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11747_/A sky130_fd_sc_hd__xor2_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07241__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _11663_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _11665_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ _11677_/B _11594_/B vssd1 vssd1 vccd1 vccd1 _11596_/C sky130_fd_sc_hd__or2_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _10545_/A _10545_/B _10545_/C vssd1 vssd1 vccd1 vccd1 _10546_/B sky130_fd_sc_hd__and3_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ instruction[14] vssd1 vssd1 vccd1 vccd1 loadstore_dest[3] sky130_fd_sc_hd__buf_12
X_10476_ _11774_/B vssd1 vssd1 vccd1 vccd1 _10476_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08072__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ _13230_/CLK _13195_/D vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__dfxtp_1
X_12215_ _12256_/B _12215_/B vssd1 vssd1 vccd1 vccd1 _12258_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10107__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__A2 _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _12146_/A _12146_/B _12146_/C vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12322__A _12502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _12047_/Y _12048_/X _12051_/Y _12076_/X vssd1 vssd1 vccd1 vccd1 _12077_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12132__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__or2_1
XANTENNA__11340__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12979_ hold257/X _06858_/B _12978_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold258/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 instruction[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_38 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ _08170_/A _08170_/B vssd1 vssd1 vccd1 vccd1 _08189_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_49 reg2_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _07158_/A _06928_/C _07108_/C _07109_/A _07303_/A vssd1 vssd1 vccd1 vccd1
+ _07123_/B sky130_fd_sc_hd__o41ai_4
XFILLER_0_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07052_ _09423_/A _07053_/B vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__or2_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07954_ _07982_/A _07982_/B _08030_/B _07953_/B _07953_/A vssd1 vssd1 vccd1 vccd1
+ _07981_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06905_ _12115_/A _06905_/B vssd1 vssd1 vccd1 vccd1 _06905_/Y sky130_fd_sc_hd__nand2_8
X_07885_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09524__B1 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__A2 _08986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _09297_/X _09305_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__mux2_1
X_06836_ _11521_/A _11431_/A _11339_/A _11240_/A vssd1 vssd1 vccd1 vccd1 _06838_/A
+ sky130_fd_sc_hd__or4b_1
XANTENNA__10134__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11882__A1 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__B2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ _09495_/B _09495_/C _09501_/A vssd1 vssd1 vccd1 vccd1 _09651_/C sky130_fd_sc_hd__a21boi_1
XFILLER_0_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09827__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09555_/Y sky130_fd_sc_hd__nand2b_1
X_06698_ reg1_val[10] _07296_/A vssd1 vssd1 vccd1 vccd1 _06699_/B sky130_fd_sc_hd__or2_1
X_09486_ _09485_/X _09289_/X _09634_/A vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__and2_1
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07061__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _08440_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08437_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08368_ _08319_/A _08319_/B _08317_/X vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12407__A _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07319_ _09568_/A _07513_/B _09428_/A fanout15/X vssd1 vssd1 vccd1 vccd1 _07320_/B
+ sky130_fd_sc_hd__o22a_1
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08354_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ instruction[7] _10329_/X _10328_/X vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10261_ _11656_/A _10261_/B vssd1 vssd1 vccd1 vccd1 _10263_/B sky130_fd_sc_hd__xor2_1
X_12000_ hold299/A _12000_/A2 _12063_/B _11999_/Y _12313_/A1 vssd1 vssd1 vccd1 vccd1
+ _12008_/B sky130_fd_sc_hd__a311o_1
XANTENNA__08566__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _06830_/D _10190_/X _10191_/Y vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09716__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__B1 _09512_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _08276_/A _12926_/A2 hold125/X vssd1 vssd1 vccd1 vccd1 _13192_/D sky130_fd_sc_hd__o21a_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ _12832_/B _12832_/C hold64/X vssd1 vssd1 vccd1 vccd1 _13109_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ hold259/X hold9/X vssd1 vssd1 vccd1 vccd1 _13024_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11715_ fanout55/X _12141_/A fanout45/X fanout63/X vssd1 vssd1 vccd1 vccd1 _11716_/B
+ sky130_fd_sc_hd__o22a_1
X_12695_ hold9/X _12730_/B _12694_/Y _13103_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__o211a_1
XFILLER_0_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11646_ _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__or2_1
X_11577_ _11468_/A _11468_/B _11473_/A vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10061__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ fanout82/X _12201_/A fanout9/X _08565_/B vssd1 vssd1 vccd1 vccd1 _10529_/B
+ sky130_fd_sc_hd__o22a_1
X_13247_ _13250_/CLK _13247_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10460_/B sky130_fd_sc_hd__nand2_1
X_13178_ _13243_/CLK _13178_/D vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ hold235/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07670_ _07670_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11864__A1 _06601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _06646_/A _12522_/B vssd1 vssd1 vccd1 vccd1 _06621_/X sky130_fd_sc_hd__or2_1
X_09340_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09340_/Y sky130_fd_sc_hd__nand2_1
X_06552_ _06552_/A _06552_/B vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10824__C1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _08945_/A _08945_/B _08943_/Y vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _08734_/A _08222_/B _08222_/C vssd1 vssd1 vccd1 vccd1 _08223_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout122_A _06963_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _08151_/A _08151_/B _08152_/X vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_15_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07104_ _12085_/A _11955_/A _07112_/B vssd1 vssd1 vccd1 vccd1 _07106_/A sky130_fd_sc_hd__nand3b_1
X_08084_ _08801_/A _08084_/B vssd1 vssd1 vccd1 vccd1 _08087_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ reg1_val[1] _07035_/B vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06690__A_N _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06879__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _08986_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _12178_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07220__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _11072_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _07942_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07868_ _07868_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06819_ _06819_/A _06819_/B vssd1 vssd1 vccd1 vccd1 _06819_/X sky130_fd_sc_hd__and2_1
X_07799_ _09309_/S _07799_/B vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__nand2_1
X_09607_ _09607_/A _09607_/B vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_109_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout35_A _07305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _09014_/A _09015_/A _11838_/A _12179_/A _09468_/Y vssd1 vssd1 vccd1 vccd1
+ _09469_/X sky130_fd_sc_hd__a311o_1
X_11500_ _11501_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ _12480_/A _12480_/B _12480_/C _12480_/D vssd1 vssd1 vccd1 vccd1 _12481_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA_fanout1_A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11431_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08787__B2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A1 _06511_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__A2 _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ _11321_/A _11321_/B _11323_/Y vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__o21ai_1
X_13101_ hold293/A _13100_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _10181_/A _10181_/B _10312_/X vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__a21oi_1
X_11293_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11304_/A sky130_fd_sc_hd__and2_1
X_13032_ hold273/X _06858_/B _13031_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold274/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10346__A1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__nor2_1
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10177_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout191 _08714_/A vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__buf_12
Xfanout180 _08607_/A vssd1 vssd1 vccd1 vccd1 _07832_/A sky130_fd_sc_hd__buf_6
XANTENNA__09832__A2_N fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ _13063_/B _13064_/A _12749_/X vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_96_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12747_ hold291/X hold17/X vssd1 vssd1 vccd1 vccd1 _13072_/B sky130_fd_sc_hd__nand2b_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ hold51/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__or2_1
XFILLER_0_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _12313_/A1 _11623_/X _11624_/Y _11628_/X vssd1 vssd1 vccd1 vccd1 _11629_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11782__A0 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07450__A1 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07450__B2 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11534__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__C1 _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08840_ _09032_/B _09033_/A _08587_/X vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08771_ _08770_/Y _08771_/B _08771_/C vssd1 vssd1 vccd1 vccd1 _08784_/A sky130_fd_sc_hd__nand3b_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07722_ _07722_/A _07722_/B _07722_/C vssd1 vssd1 vccd1 vccd1 _07811_/B sky130_fd_sc_hd__and3_1
X_07653_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__xnor2_2
X_06604_ _11858_/S _06604_/B vssd1 vssd1 vccd1 vccd1 _06837_/A sky130_fd_sc_hd__nor2_1
X_09323_ _09308_/X _09322_/X _10809_/A vssd1 vssd1 vccd1 vccd1 _09324_/A sky130_fd_sc_hd__mux2_1
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07585_/B sky130_fd_sc_hd__xnor2_2
X_06535_ instruction[1] _06850_/B instruction[25] pred_val vssd1 vssd1 vccd1 vccd1
+ _06535_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__A_N fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ _09255_/A _09255_/B vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__nand2_1
X_09185_ _07513_/B _10117_/A _09880_/B2 fanout14/X vssd1 vssd1 vccd1 vccd1 _09186_/B
+ sky130_fd_sc_hd__o22a_1
X_08205_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08249_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__B2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _11470_/A _08136_/B vssd1 vssd1 vccd1 vccd1 _08137_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _11169_/A _08219_/B _08815_/B _11297_/A vssd1 vssd1 vccd1 vccd1 _08068_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07018_ _10009_/A _12712_/A _09725_/B2 _12714_/A vssd1 vssd1 vccd1 vccd1 _07019_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10205__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08969_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12420__A _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11980_ _11980_/A _11980_/B vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__or2_1
X_10931_ _12000_/A2 _11037_/B hold297/A vssd1 vssd1 vccd1 vccd1 _10931_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07514__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ _10863_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__and2_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12602_/B _12602_/C _12620_/A vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__a21oi_4
X_10793_ _10677_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10793_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11056__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ reg1_val[7] _12532_/B vssd1 vssd1 vccd1 vccd1 _12533_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10264__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ reg1_val[22] curr_PC[22] _12495_/S vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ _11416_/A _11506_/B _11414_/C vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__and3_1
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _12403_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _12396_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08337__A_N _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__B1 _09146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11345_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11276_ _11390_/B _11276_/B vssd1 vssd1 vccd1 vccd1 _11278_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09709__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _13015_/A _13015_/B vssd1 vssd1 vccd1 vccd1 _13015_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09185__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _10529_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07196__B1 _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_10158_ _10159_/A _10159_/B _10157_/Y vssd1 vssd1 vccd1 vccd1 _10158_/X sky130_fd_sc_hd__o21ba_1
X_10089_ _09330_/A _10075_/Y _10088_/Y _09124_/S _10086_/X vssd1 vssd1 vccd1 vccd1
+ _10089_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12330__A _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11295__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08999__A1 _09001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A2 _09637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__B1 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10009__B fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09941_ _11696_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06529__A3 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ fanout83/X fanout58/X fanout55/X _06940_/A vssd1 vssd1 vccd1 vccd1 _09873_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08823_ _09333_/A _08823_/B vssd1 vssd1 vccd1 vccd1 _09015_/A sky130_fd_sc_hd__nand2b_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ _08753_/A _08753_/B _08753_/C vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07705_ _07705_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__xor2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__or2_1
XANTENNA__08687__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07637_/B vssd1 vssd1 vccd1 vccd1 _07636_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06701__A3 _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ _07567_/A _07567_/B vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07988__B _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09304_/X _09305_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09306_/X sky130_fd_sc_hd__mux2_1
X_06518_ reg1_val[30] vssd1 vssd1 vccd1 vccd1 _06800_/A sky130_fd_sc_hd__inv_2
X_07498_ _07699_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__or2_1
X_09237_ _09237_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10797__A1 _11230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__A_N _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06870__C1 _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09168_/A _09168_/B vssd1 vssd1 vccd1 vccd1 _12302_/B sky130_fd_sc_hd__or2_2
XFILLER_0_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _09097_/X _09098_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09099_/X sky130_fd_sc_hd__mux2_1
X_08119_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__xor2_4
X_11130_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12171__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _11656_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11063_/B sky130_fd_sc_hd__xnor2_1
X_10012_ _10011_/B _10012_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _11965_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07350__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914_ _11238_/A _10914_/B _10914_/C vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__and3_1
X_11894_ _11895_/A _11895_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__o21a_1
X_10845_ _10845_/A _10845_/B _10845_/C vssd1 vssd1 vccd1 vccd1 _10847_/A sky130_fd_sc_hd__and3_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10237__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10776_ _10776_/A _10776_/B _10776_/C vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__or3_1
X_12515_ _12514_/A _12511_/Y _12513_/B vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_35_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ _12496_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ reg1_val[9] curr_PC[9] _12444_/S vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06759__A3 _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07419__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _11328_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11259_ _09064_/Y _11135_/X _11247_/B _09135_/Y _11258_/Y vssd1 vssd1 vccd1 vccd1
+ _11259_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12701__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09634__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08905__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11268__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06993__A _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08470_ _08471_/B _08471_/A vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08133__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07421_ _12684_/A fanout36/X fanout34/X _12686_/A vssd1 vssd1 vccd1 vccd1 _07422_/B
+ sky130_fd_sc_hd__o22a_1
X_07352_ _07438_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07283_ reg1_val[19] _07283_/B vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_5_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__nand2_1
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13188_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09397__A1 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__B2 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__buf_1
XANTENNA__09149__A1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09678__A2_N _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _12263_/S _09924_/B _09924_/C vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__or3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09855_ _09855_/A _09855_/B _09855_/C vssd1 vssd1 vccd1 vccd1 _09856_/B sky130_fd_sc_hd__nand3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06887__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _09420_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08812_/A sky130_fd_sc_hd__xnor2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _09495_/A _09784_/X _09785_/X vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__o21a_1
X_06998_ _10481_/A vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__inv_2
X_08737_ _08756_/B2 _08737_/A2 _08813_/B1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 _08738_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07999__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08668_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08124__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07619_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__and2_1
XANTENNA__09872__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _11799_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _10632_/B sky130_fd_sc_hd__xnor2_1
X_08599_ _08740_/A2 _08733_/B1 _08735_/A2 _08755_/B vssd1 vssd1 vccd1 vccd1 _08600_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__C1 _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A1 _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _10319_/B _10794_/B _10792_/B vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__a21o_2
X_12300_ _12299_/A _12299_/B _09145_/Y vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__o21ai_1
X_10492_ _11295_/B2 fanout47/X _11297_/A fanout13/X vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12231_ hold293/A _12230_/B _12304_/B1 vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07938__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _11873_/A _11873_/B _11907_/Y _11975_/Y _12161_/Y vssd1 vssd1 vccd1 vccd1
+ _12167_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__08060__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__A _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ _12146_/B _12098_/B vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__and2_1
X_11113_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11114_/C sky130_fd_sc_hd__xnor2_1
X_11044_ _11043_/A _09141_/Y _11043_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _11044_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09560__A1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B2 _07056_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _12995_/A _12995_/B vssd1 vssd1 vccd1 vccd1 _12995_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ _12245_/B _11946_/B vssd1 vssd1 vccd1 vccd1 _11948_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07323__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__A1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__B2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _11948_/A _11877_/B vssd1 vssd1 vccd1 vccd1 _11879_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10828_ _10828_/A vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11958__B1 fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10759_ fanout78/X _12201_/A fanout9/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10760_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12429_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08051__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__A1 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _08039_/B _08039_/A vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__nand2b_1
X_06921_ _10529_/A _06939_/A vssd1 vssd1 vccd1 vccd1 _06921_/X sky130_fd_sc_hd__and2_1
XANTENNA__12502__B _12502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11489__A2 _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06852_ instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1 vccd1 _06852_/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09640_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__or2_1
XANTENNA__09551__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06783_ _11124_/B _11124_/C _06831_/A vssd1 vssd1 vccd1 vccd1 _11238_/C sky130_fd_sc_hd__o21ai_1
X_09571_ _11885_/A _09571_/B vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__xnor2_1
X_08522_ _08782_/A2 _08715_/A2 _08689_/B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08523_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10957__B _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07865__B2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__A1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07335_ _07335_/A _07335_/B _07335_/C vssd1 vssd1 vccd1 vccd1 _07336_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_73_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__B2 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10973__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ _12142_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__or2_1
XFILLER_0_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _09005_/A _09005_/B vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07197_ _09423_/A _07197_/B vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12677__A1 _07110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__xor2_2
X_09769_ _09769_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _11801_/A _11801_/B vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__or2_1
X_12780_ hold294/A hold51/X vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ _11803_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__and2_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10860__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08805__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _11593_/A _11593_/B _11593_/C vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__and3_1
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10613_ _10500_/A _10500_/B _10496_/A vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__o21ai_1
X_10544_ _10545_/A _10545_/B _10545_/C vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10475_ _10809_/A _10074_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__o21ai_1
X_13263_ instruction[13] vssd1 vssd1 vccd1 vccd1 loadstore_dest[2] sky130_fd_sc_hd__buf_12
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13194_ _13230_/CLK hold112/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__dfxtp_1
X_12214_ _12214_/A _12214_/B _12214_/C vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__or3_1
XFILLER_0_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _12146_/A _12146_/B _12146_/C vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ _12265_/C1 _12055_/Y _12056_/X _12075_/Y vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__a31o_1
X_11027_ _11026_/A _11026_/B _11026_/Y _09498_/A vssd1 vssd1 vccd1 vccd1 _11027_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__06898__A2 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13093__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ hold296/A _12977_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ hold231/A _11620_/B _12001_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _11930_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 instruction[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07120_ _06928_/C _07108_/C _07109_/A _07303_/A vssd1 vssd1 vccd1 vccd1 _07158_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _07051_/A _07051_/B vssd1 vssd1 vccd1 vccd1 _07053_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07953_ _07953_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06511__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _11238_/A _06905_/B vssd1 vssd1 vccd1 vccd1 _06904_/X sky130_fd_sc_hd__and2_1
X_07884_ _07884_/A _07884_/B vssd1 vssd1 vccd1 vccd1 _07886_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09524__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ _06835_/A _06835_/B _06835_/C vssd1 vssd1 vccd1 vccd1 _06839_/B sky130_fd_sc_hd__and3_1
X_09623_ _09295_/X _09298_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11882__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ _06761_/A _06761_/B _09309_/S _06511_/Y vssd1 vssd1 vccd1 vccd1 _09495_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09827__A2 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ _09979_/A _09554_/B vssd1 vssd1 vccd1 vccd1 _09556_/B sky130_fd_sc_hd__xnor2_1
X_06697_ reg1_val[10] _07296_/A vssd1 vssd1 vccd1 vccd1 _10586_/S sky130_fd_sc_hd__nand2_1
X_09485_ _09118_/X _09122_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08505_ _08513_/A _08513_/B _08495_/X vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08436_ _08814_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08440_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11799__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__nor2_2
X_07318_ _07916_/A _07318_/B vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08298_ _10853_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07249_ _07249_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07261_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09212__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ _11295_/B2 _07988_/B _10359_/B2 fanout50/X vssd1 vssd1 vccd1 vccd1 _10261_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08566__A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _06830_/D _10190_/X _09498_/A vssd1 vssd1 vccd1 vccd1 _10191_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09515__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ hold90/X _12662_/A _13112_/B hold124/X _13013_/A vssd1 vssd1 vccd1 vccd1
+ hold125/A sky130_fd_sc_hd__o221a_1
XANTENNA__07526__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ hold64/X _12832_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__and3_1
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ hold9/X hold259/X vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__and2b_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11153_/A _11710_/X _11711_/X _11713_/Y vssd1 vssd1 vccd1 vccd1 dest_val[21]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__10833__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ _12694_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _12694_/Y sky130_fd_sc_hd__nand2_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11723_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11647_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09179__A _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ _11483_/A _11483_/B _11479_/Y vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10527_ _10527_/A vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13246_ _13246_/CLK _13246_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10458_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10458_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09203__B1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _13246_/CLK hold181/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07765__B1 _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__or2_1
X_12128_ hold302/A _12304_/B1 _12184_/B _12127_/Y _09810_/A vssd1 vssd1 vccd1 vccd1
+ _12128_/X sky130_fd_sc_hd__a311o_1
X_12059_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06620_ instruction[30] _06637_/B vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__and2_4
XFILLER_0_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11864__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ reg1_val[26] _07064_/A vssd1 vssd1 vccd1 vccd1 _06552_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11077__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _08899_/A _08899_/B _08898_/A vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08221_ _08222_/B _08222_/C _08734_/A vssd1 vssd1 vccd1 vccd1 _08223_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _08316_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08152_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07103_ _07103_/A _07103_/B vssd1 vssd1 vccd1 vccd1 _07112_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08083_ _10876_/A1 _08782_/A2 _08756_/B2 _10957_/A vssd1 vssd1 vccd1 vccd1 _08084_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout115_A _06999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ _12501_/A _07035_/B vssd1 vssd1 vccd1 vccd1 _08276_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10462__S _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A1 _07044_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08985_ _08985_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07220__A2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B2 _07069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07936_ _09885_/A fanout43/X _08333_/B _09880_/B2 vssd1 vssd1 vccd1 vccd1 _07937_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09552__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07867_ _07868_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07867_/X sky130_fd_sc_hd__or2_1
X_06818_ _06803_/Y _06817_/X _12175_/A vssd1 vssd1 vccd1 vccd1 _06819_/B sky130_fd_sc_hd__a21o_1
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__nor2_1
X_09606_ _09607_/B _09607_/A vssd1 vssd1 vccd1 vccd1 _09606_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12265__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06749_ _06763_/B _06646_/A _12512_/B _06748_/X vssd1 vssd1 vccd1 vccd1 _06749_/X
+ sky130_fd_sc_hd__a31o_1
X_09537_ _09537_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09538_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09015_/A _11838_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _09468_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout28_A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__B1 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08421_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _09399_/A vssd1 vssd1 vccd1 vccd1 _09406_/A sky130_fd_sc_hd__inv_2
X_11430_ _06787_/X _11429_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07011__S _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _11334_/X _11360_/X _11267_/X vssd1 vssd1 vccd1 vccd1 dest_val[17] sky130_fd_sc_hd__a21oi_4
X_13100_ _13100_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _13100_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11791__A1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__A _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _10048_/A _10048_/B _10181_/A _10181_/B vssd1 vssd1 vccd1 vccd1 _10312_/X
+ sky130_fd_sc_hd__o22a_1
X_11292_ _11399_/B _11292_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__nor2_1
X_13031_ hold297/A _13030_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11543__A1 _06980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__xnor2_1
X_10174_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__nor2_1
Xfanout192 _07689_/A vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__buf_12
Xfanout181 _06917_/Y vssd1 vssd1 vccd1 vccd1 _08607_/A sky130_fd_sc_hd__buf_12
Xfanout170 _09222_/B2 vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__buf_6
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12815_ _13059_/A _12814_/B _12751_/X vssd1 vssd1 vccd1 vccd1 _13064_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10806__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ hold17/X hold291/X vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08806__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ _07110_/Y _12731_/A2 hold46/X _13111_/A vssd1 vssd1 vccd1 vccd1 _13131_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _09293_/A _10700_/X _10713_/Y _09330_/A _11627_/X vssd1 vssd1 vccd1 vccd1
+ _11628_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11782__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09059__D _12299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ _11560_/B _11559_/B vssd1 vssd1 vccd1 vccd1 _11662_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07450__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08541__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ _13230_/CLK _13229_/D vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07157__A _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06996__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _09423_/A _08770_/B vssd1 vssd1 vccd1 vccd1 _08770_/Y sky130_fd_sc_hd__xnor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07721_ _11955_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07722_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11298__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ reg1_val[23] _07028_/A vssd1 vssd1 vccd1 vccd1 _06604_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07583_/X sky130_fd_sc_hd__or2_1
XANTENNA__07910__B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06534_ instruction[1] _06850_/B instruction[25] pred_val vssd1 vssd1 vccd1 vccd1
+ _06534_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09322_ _09315_/X _09321_/X _10924_/S vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09663__B1 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08716__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _11796_/A _09253_/B vssd1 vssd1 vccd1 vccd1 _09255_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ _09373_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09188_/B sky130_fd_sc_hd__or2_1
X_08204_ _08204_/A _08204_/B vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ _12668_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08136_/B sky130_fd_sc_hd__or2_1
XFILLER_0_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ _08077_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ _07028_/A _07017_/B vssd1 vssd1 vccd1 vccd1 _07017_/Y sky130_fd_sc_hd__xnor2_1
X_08968_ _07637_/A _07636_/Y _07640_/A vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__a21oi_2
X_08899_ _08899_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__xor2_4
X_07919_ _09420_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__xnor2_1
X_10930_ hold259/A _10930_/B vssd1 vssd1 vccd1 vccd1 _11037_/B sky130_fd_sc_hd__or2_1
XANTENNA__12238__C1 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12600_ _12615_/B _12600_/B vssd1 vssd1 vccd1 vccd1 _12602_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _11068_/A _10861_/B vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__xnor2_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ _10794_/A _10792_/B _10794_/C vssd1 vssd1 vccd1 vccd1 _10792_/X sky130_fd_sc_hd__and3_1
XANTENNA__10875__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ reg1_val[7] _12532_/B vssd1 vssd1 vccd1 vccd1 _12531_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12148__A _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__A1 _11091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__B2 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ _12468_/B _12462_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11413_ _11506_/B _11414_/C vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ _12553_/B _12393_/B vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11344_ _11342_/Y _11344_/B vssd1 vssd1 vccd1 vccd1 _11345_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11275_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11276_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09709__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ _12767_/X _13014_/B vssd1 vssd1 vccd1 vccd1 _13015_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09185__A2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ _06940_/Y _10845_/A _10845_/B _07044_/Y _10393_/A vssd1 vssd1 vccd1 vccd1
+ _10227_/B sky130_fd_sc_hd__a32o_1
XANTENNA__07196__A1 _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__B2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_10157_ _10157_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__xnor2_1
X_10088_ _10203_/S _10087_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10088_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__12229__C1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ hold7/X _12730_/B _12728_/Y _13111_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o211a_1
XFILLER_0_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10007__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08271__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09940_ _11135_/S _09939_/X _09936_/X vssd1 vssd1 vccd1 vccd1 _09940_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap178 _06943_/B vssd1 vssd1 vccd1 vccd1 _06979_/B sky130_fd_sc_hd__clkbuf_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10191__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _06764_/X _08384_/B _07185_/Y _12499_/A vssd1 vssd1 vccd1 vccd1 _09333_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08753_/A _08753_/B _08753_/C vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__and3_1
XANTENNA__10730__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12240__B _12240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _07875_/A _07704_/B vssd1 vssd1 vccd1 vccd1 _07705_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08684_ _08704_/A _08704_/B vssd1 vssd1 vccd1 vccd1 _08706_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08687__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08687__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _07274_/B _12095_/B _07635_/S vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__mux2_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07567_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08446__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06517_ reg1_val[26] vssd1 vssd1 vccd1 vccd1 _07103_/A sky130_fd_sc_hd__inv_2
X_09305_ _09089_/X _09091_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _08916_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07699_/B sky130_fd_sc_hd__xnor2_1
X_09236_ _09356_/A _09235_/C _09235_/A vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09167_ _09168_/B vssd1 vssd1 vccd1 vccd1 _09167_/Y sky130_fd_sc_hd__inv_2
X_09098_ reg1_val[9] reg1_val[22] _09120_/S vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__mux2_1
X_08118_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _10853_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08050_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout95_A _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ _11876_/A fanout50/X _07988_/B _11950_/A vssd1 vssd1 vccd1 vccd1 _11061_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _10012_/B _10011_/B vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07525__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11962_ _12023_/B _11962_/B vssd1 vssd1 vccd1 vccd1 _11964_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09740__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07350__A1 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11893_ _11964_/B _11893_/B vssd1 vssd1 vccd1 vccd1 _11895_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11682__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ _11232_/A _10913_/B _10913_/C vssd1 vssd1 vccd1 vccd1 _10913_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__07350__B2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10844_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__B2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10237__A1 fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xor2_4
XFILLER_0_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ _10776_/A _10776_/B _10776_/C vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ _12496_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12455_/C sky130_fd_sc_hd__nand2_1
X_12376_ _12382_/B _12376_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XFILLER_0_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ _11327_/A _11327_/B _11327_/C vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10126__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _11250_/Y _11251_/X _11254_/X _11257_/Y vssd1 vssd1 vccd1 vccd1 _11258_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10209_ _10208_/B _10465_/C hold241/A vssd1 vssd1 vccd1 vccd1 _10209_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08905__A2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ _11189_/A _11278_/A _11189_/C vssd1 vssd1 vccd1 vccd1 _11190_/B sky130_fd_sc_hd__or3_1
XANTENNA__09126__S _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09866__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06695__A3 _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ _11468_/A _07351_/B vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11425__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10228__A1 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10228__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07282_ reg1_val[19] _07283_/B vssd1 vssd1 vccd1 vccd1 _07282_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _09022_/B sky130_fd_sc_hd__nor2_1
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__B2 _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09397__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold301/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__buf_1
X_09923_ _06739_/Y _09784_/X _06741_/B vssd1 vssd1 vccd1 vccd1 _09923_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09149__A2 _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09854_ _09855_/A _09855_/B _09855_/C vssd1 vssd1 vccd1 vccd1 _09854_/Y sky130_fd_sc_hd__a21oi_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _06828_/A _09568_/A _08813_/B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 _08806_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _06999_/B _06999_/A _07832_/A vssd1 vssd1 vccd1 vccd1 _06997_/X sky130_fd_sc_hd__mux2_1
X_09785_ _12263_/S _09785_/B _09785_/C vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__or3_1
X_08736_ _08814_/A _08736_/B vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__xnor2_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08662_/A _08662_/B _08686_/A vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__o21ai_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07618_ _11184_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _08601_/A _08601_/B vssd1 vssd1 vccd1 vccd1 _08616_/A sky130_fd_sc_hd__nor2_1
X_07549_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07550_/B sky130_fd_sc_hd__or2_1
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__B1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout10_A _12728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10319_/A _10560_/B vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__and2b_1
X_09219_ _11184_/A _09219_/B vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__xnor2_1
X_10491_ _12089_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ hold293/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12272_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08596__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ _12161_/A vssd1 vssd1 vccd1 vccd1 _12161_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08060__A2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12092_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__or2_1
X_11112_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11226_/B sky130_fd_sc_hd__or2_1
X_11043_ _11043_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11043_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10155__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12695__A2 _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07255__A _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__C1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _12775_/X _12994_/B vssd1 vssd1 vccd1 vccd1 _12995_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07323__A1 _07110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ fanout60/X fanout7/X fanout5/X _12095_/A vssd1 vssd1 vccd1 vccd1 _11946_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11655__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__B2 _07147_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08520__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__A3 _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07874__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ _11876_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08086__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827_ _10809_/A _09636_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11958__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08814__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__B2 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10758_ _10652_/A _10652_/B _10650_/Y vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12428_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__a21o_1
X_10689_ _11238_/A _10689_/B _10689_/C vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__and3_1
XANTENNA__12336__A _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__C1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12359_ _12368_/A _12359_/B vssd1 vssd1 vccd1 vccd1 _12361_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10394__B1 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12135__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12135__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ _10607_/A _06922_/B vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__nor2_1
X_06851_ dest_pred_val _06887_/B _06847_/X vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
XANTENNA__09551__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06782_ _11023_/B _11023_/C _11026_/A vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__a21boi_1
X_09570_ _09885_/A fanout8/X fanout6/X _09698_/A vssd1 vssd1 vccd1 vccd1 _09571_/B
+ sky130_fd_sc_hd__o22a_1
X_08521_ _08814_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08528_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08452_ _08452_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06509__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ _07403_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07865__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout145_A _07137_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _08801_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12071__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07617__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07265_ reg1_val[30] _07265_/B vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09004_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ _12720_/A _09222_/B2 _12718_/A _09422_/A vssd1 vssd1 vccd1 vccd1 _07197_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07250__B1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09906_ _09907_/B _09907_/A vssd1 vssd1 vccd1 vccd1 _09906_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12677__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07075__A _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__nor2_1
X_09768_ _09769_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout58_A _12716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08752_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13016__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11730_/A _11730_/B vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__nand2_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09699_ _09564_/A _09564_/B _09562_/X vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__o21a_2
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11574_/A _11574_/B _11572_/Y vssd1 vssd1 vccd1 vccd1 _11671_/A sky130_fd_sc_hd__o21a_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10860__A1 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10860__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__A1 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _11593_/A _11593_/B _11593_/C vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__and2_1
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08805__B2 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ _10403_/A _10403_/C _10403_/B vssd1 vssd1 vccd1 vccd1 _10545_/C sky130_fd_sc_hd__a21boi_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10474_ _10466_/Y _10467_/X _10473_/X vssd1 vssd1 vccd1 vccd1 _10474_/Y sky130_fd_sc_hd__o21ai_1
X_13262_ instruction[12] vssd1 vssd1 vccd1 vccd1 loadstore_dest[1] sky130_fd_sc_hd__buf_12
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13193_ _13230_/CLK hold154/X vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
X_12213_ _12214_/A _12214_/B _12214_/C vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__o21ai_2
X_12144_ _12245_/B _12144_/B vssd1 vssd1 vccd1 vccd1 _12146_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12075_ _06890_/X _12062_/X _12074_/X vssd1 vssd1 vccd1 vccd1 _12075_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06601__B _06601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11026_ _11026_/A _11026_/B vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06752__C1 _12507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13093__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ _12977_/A _12977_/B vssd1 vssd1 vccd1 vccd1 _12977_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11235__A _11235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11928_ _11620_/B _12001_/B hold231/A vssd1 vssd1 vccd1 vccd1 _11930_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ reg1_val[23] _07028_/A _09138_/X _11858_/X vssd1 vssd1 vccd1 vccd1 _11859_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_18 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07050_ _07050_/A _07050_/B vssd1 vssd1 vccd1 vccd1 _07051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10906__A2 _10796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09375__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _07982_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__nand2_1
X_07883_ _07883_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__or2_1
X_06903_ _09146_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _06905_/B sky130_fd_sc_hd__nor2_2
XANTENNA__09524__A2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ _06834_/A _06834_/B _06834_/C _06834_/D vssd1 vssd1 vccd1 vccd1 _06835_/C
+ sky130_fd_sc_hd__and4_1
X_09622_ _09621_/A _09621_/C _09621_/B vssd1 vssd1 vccd1 vccd1 _09622_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10134__A3 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _11387_/A fanout42/X _07239_/A fanout71/X vssd1 vssd1 vccd1 vccd1 _09554_/B
+ sky130_fd_sc_hd__o22a_1
X_06765_ _06700_/B _06762_/X _06763_/X vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09288__A1 _09617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ _08561_/A _08561_/B _08503_/A vssd1 vssd1 vccd1 vccd1 _08513_/B sky130_fd_sc_hd__o21a_1
X_09484_ _09483_/X _09482_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ _07296_/A reg1_val[10] vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _08274_/A _10957_/A _08813_/A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 _08436_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ _08366_/A _08366_/B vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__and2_1
XFILLER_0_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ _10117_/A fanout49/X _09880_/B2 fanout51/X vssd1 vssd1 vccd1 vccd1 _07318_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10055__C1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ _08430_/B _08737_/A2 _09428_/A fanout79/X vssd1 vssd1 vccd1 vccd1 _08298_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07248_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07179_ _07263_/C _12639_/B _07128_/A vssd1 vssd1 vccd1 vccd1 _07180_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__09212__A1 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__A _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _06772_/Y _10189_/X _12263_/S vssd1 vssd1 vccd1 vccd1 _10190_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09212__B2 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__A0 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A1 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _13013_/A hold91/X vssd1 vssd1 vccd1 vccd1 _13191_/D sky130_fd_sc_hd__and2_1
XANTENNA__07526__B2 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _13104_/A _13104_/B vssd1 vssd1 vccd1 vccd1 _12832_/C sky130_fd_sc_hd__or2_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ hold297/A hold62/X vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__nand2b_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _07277_/X _12731_/A2 hold71/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13139_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A _11866_/C vssd1 vssd1 vccd1 vccd1 _11713_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11643_/B _11644_/B vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11465_/Y _11474_/B _11486_/A vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ _11072_/A _10526_/B vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__xnor2_1
X_13245_ _13246_/CLK _13245_/D vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10457_ _10337_/A _10334_/Y _10336_/B vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09203__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _13243_/CLK _13176_/D vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__dfxtp_1
X_10388_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10545_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12127_ _12304_/B1 _12184_/B hold302/A vssd1 vssd1 vccd1 vccd1 _12127_/Y sky130_fd_sc_hd__a21oi_1
X_12058_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11009_ _11010_/B _11010_/A vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07443__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ reg1_val[26] _07064_/A vssd1 vssd1 vccd1 vccd1 _06552_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11077__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__B2 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ _06938_/A _06938_/B _08815_/B vssd1 vssd1 vccd1 vccd1 _08222_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08274__A _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07102_ reg1_val[25] _07102_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__xnor2_4
X_08082_ _08814_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08087_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07033_ _12499_/A reg1_val[31] _09495_/A vssd1 vssd1 vccd1 vccd1 _07035_/B sky130_fd_sc_hd__and3_4
XFILLER_0_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09309__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__B _09817_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout108_A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11552__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ _12115_/A _12297_/A vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07935_ _07955_/A _08027_/A _07955_/C vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09833__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _11072_/A _07866_/B vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__xor2_1
X_09605_ _09605_/A _09605_/B vssd1 vssd1 vccd1 vccd1 _09607_/B sky130_fd_sc_hd__xnor2_1
X_06817_ _12115_/B _12115_/C _12117_/A vssd1 vssd1 vccd1 vccd1 _06817_/X sky130_fd_sc_hd__a21o_1
X_07797_ _07797_/A _07797_/B _07858_/A vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__nor3_1
X_06748_ reg2_val[2] _06748_/B vssd1 vssd1 vccd1 vccd1 _06748_/X sky130_fd_sc_hd__and2_1
X_09536_ _09534_/A _09534_/B _09537_/B vssd1 vssd1 vccd1 vccd1 _09536_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _09617_/C _09465_/Y _09466_/Y vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12017__B1 _11887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06679_ _10920_/A _06960_/A vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09681__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ _10252_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__xnor2_1
X_08349_ _08350_/A _08349_/B _08349_/C vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11335_/Y _11336_/X _11359_/X vssd1 vssd1 vccd1 vccd1 _11360_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _10311_/A _10311_/B _10049_/X vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_15_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13030_ _13030_/A _13030_/B vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__xnor2_1
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09727__B fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10242_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__and2_1
XANTENNA__11543__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _10039_/A _10039_/B _10037_/Y vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout171 _07041_/Y vssd1 vssd1 vccd1 vccd1 _09222_/B2 sky130_fd_sc_hd__buf_8
Xfanout182 _09136_/Y vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__buf_4
Xfanout160 _09428_/A vssd1 vssd1 vccd1 vccd1 _08813_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11700__C1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout193 _06925_/X vssd1 vssd1 vccd1 vccd1 _07303_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12814_ _12751_/X _12814_/B vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12745_ hold29/X hold292/A vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ hold45/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__or2_1
XFILLER_0_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11627_ _07012_/B _06905_/Y _11626_/X _06628_/B vssd1 vssd1 vccd1 vccd1 _11627_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11232__B _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11558_ _12086_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10509_ _11656_/A _10509_/B vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12344__A _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11489_ _11387_/A _11458_/A _11459_/B _11391_/A vssd1 vssd1 vccd1 vccd1 _11491_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13228_ _13234_/CLK _13228_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12731__A1 _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ _13254_/CLK _13159_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__12192__C1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _09309_/S _07154_/X _07799_/B _07185_/Y vssd1 vssd1 vccd1 vccd1 _07721_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11298__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__B2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07652_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06602_ reg1_val[23] _07028_/A vssd1 vssd1 vccd1 vccd1 _11858_/S sky130_fd_sc_hd__and2_1
X_07582_ _12142_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12247__A0 _12728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__B2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A0 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ _09320_/X _09317_/X _09634_/A vssd1 vssd1 vccd1 vccd1 _09321_/X sky130_fd_sc_hd__mux2_1
X_06533_ instruction[25] _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__and2_2
XFILLER_0_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09252_ fanout51/X _07763_/B _10647_/A fanout49/X vssd1 vssd1 vccd1 vccd1 _09253_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08203_ _08203_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__xnor2_4
X_09183_ _09182_/B _09183_/B vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08134_ _11072_/A _08134_/B vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09828__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08077_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10981__B1 _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07016_ _07028_/B _07065_/A _07028_/C _07028_/D _07058_/B1 vssd1 vssd1 vccd1 vccd1
+ _07017_/B sky130_fd_sc_hd__o41a_1
XANTENNA__07348__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__C1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _07627_/A _07627_/B _07625_/X vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ _08898_/A _08898_/B vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__nor2_2
X_07918_ _08274_/A _11739_/A _08765_/A _11663_/A vssd1 vssd1 vccd1 vccd1 _07919_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08179__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07849_ _07946_/A _07946_/B vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__nor2_1
X_10860_ _12095_/A fanout37/X _08233_/B fanout60/X vssd1 vssd1 vccd1 vccd1 _10861_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout40_A fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _11883_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__xnor2_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10791_ _10791_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__nor2_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ _12529_/A _12526_/Y _12528_/B vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10264__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _12468_/A _12457_/Y _12453_/A vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12148__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11412_ _11412_/A _11412_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11414_/C sky130_fd_sc_hd__or3_1
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12392_ _12553_/B _12393_/B vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08642__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11343_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08090__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__or2_1
XANTENNA__09709__A2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ _13013_/A hold278/X vssd1 vssd1 vccd1 vccd1 _13233_/D sky130_fd_sc_hd__and2_1
XANTENNA__08917__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _10180_/A _10180_/B _10178_/X vssd1 vssd1 vccd1 vccd1 _10308_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07196__A2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__xor2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _11134_/S _09321_/X _09166_/B vssd1 vssd1 vccd1 vccd1 _10087_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07721__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10989_ _10989_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10991_/B sky130_fd_sc_hd__nand2_1
X_12728_ _12728_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _12728_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11452__B2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ hold133/X hold161/X hold164/A hold100/X vssd1 vssd1 vccd1 vccd1 hold162/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07120__A2 _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10007__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A2 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08081__B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08821_ _08821_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__xor2_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__B1 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12521__B _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08752_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _08753_/C sky130_fd_sc_hd__nor2_1
X_07703_ _09698_/A fanout41/X _08135_/B _09885_/A vssd1 vssd1 vccd1 vccd1 _07704_/B
+ sky130_fd_sc_hd__o22a_1
X_08683_ _08683_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout175_A _07015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _08901_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08687__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09322__S _10924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07631__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _07565_/A _07565_/B _07565_/C vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__or3_1
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06516_ reg1_val[22] vssd1 vssd1 vccd1 vccd1 _06608_/A sky130_fd_sc_hd__inv_2
X_09304_ _09085_/X _09088_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09304_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07496_ fanout82/X _12694_/A _10490_/B2 _06940_/A vssd1 vssd1 vccd1 vccd1 _07497_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11153__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _09235_/A _09356_/A _09235_/C vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09166_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09558__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ reg1_val[8] reg1_val[23] _09120_/S vssd1 vssd1 vccd1 vccd1 _09097_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08117_ _08814_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07078__A _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ fanout79/X _08733_/B1 _08735_/A2 _08430_/B vssd1 vssd1 vccd1 vccd1 _08049_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12712__A _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__A0 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__A _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout88_A _07304_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _10126_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__xnor2_1
X_09999_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__nor2_1
X_11961_ _11961_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11962_/B sky130_fd_sc_hd__nor2_1
X_10912_ _11232_/A _10913_/C _10913_/B vssd1 vssd1 vccd1 vccd1 _10912_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07350__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _11892_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__and2_1
XANTENNA__11682__A1 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10843_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__A2 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ _10622_/A _10622_/B _10620_/X vssd1 vssd1 vccd1 vccd1 _10776_/C sky130_fd_sc_hd__a21o_1
X_12513_ _12511_/Y _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12444_ reg1_val[19] curr_PC[19] _12444_/S vssd1 vssd1 vccd1 vccd1 _12446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12934__A1 _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ _12375_/A _12375_/B _12375_/C vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _11326_/A vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__inv_2
XFILLER_0_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _06662_/B _11255_/Y _11256_/X vssd1 vssd1 vccd1 vccd1 _11257_/Y sky130_fd_sc_hd__a21oi_2
X_10208_ hold241/A _10208_/B _10465_/C vssd1 vssd1 vccd1 vccd1 _10208_/X sky130_fd_sc_hd__and3_1
XANTENNA__07716__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _11278_/A _11189_/C _11189_/A vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11238__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _10139_/A _10139_/B vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09866__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10796__B _10796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07350_ _12686_/A fanout36/X _08233_/B _12688_/A vssd1 vssd1 vccd1 vccd1 _07351_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07281_ reg1_val[13] _07091_/B _07091_/C _07088_/B _07128_/A vssd1 vssd1 vccd1 vccd1
+ _07283_/B sky130_fd_sc_hd__o41a_4
X_09020_ _10187_/B _10187_/C vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12516__B _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__A2 _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__B1 _10935_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__clkbuf_2
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09922_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ _09714_/A _09714_/B _09713_/A vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout292_A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _06745_/Y _09650_/Y _06747_/B vssd1 vssd1 vccd1 vccd1 _09784_/X sky130_fd_sc_hd__o21a_1
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__xor2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13102__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06996_ _10252_/A _06996_/B vssd1 vssd1 vccd1 vccd1 _06999_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09841__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _08813_/A1 _08735_/A2 _08735_/B1 _08274_/A vssd1 vssd1 vccd1 vccd1 _08736_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__C1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__nand2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07617_ _10099_/A1 fanout79/X _08430_/B _10359_/B2 vssd1 vssd1 vccd1 vccd1 _07618_/B
+ sky130_fd_sc_hd__o22a_1
X_08597_ _08714_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08601_/B sky130_fd_sc_hd__xnor2_1
X_07548_ _07664_/B _07664_/A vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07479_ fanout43/X _12686_/A _12688_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _07480_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10926__S _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ fanout78/X _11387_/A fanout71/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _09219_/B
+ sky130_fd_sc_hd__o22a_1
X_10490_ _10876_/A1 fanout11/X fanout44/X _10490_/B2 vssd1 vssd1 vccd1 vccd1 _10491_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09149_ _12179_/A _09148_/X _08823_/B vssd1 vssd1 vccd1 vccd1 _09149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ _12160_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08596__A1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__B2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11005_/A _11003_/X _11002_/Y vssd1 vssd1 vccd1 vccd1 _11113_/B sky130_fd_sc_hd__o21a_1
X_12091_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ hold171/A _11781_/B _11140_/B _11041_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1
+ _11042_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10155__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__B1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__B1 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12993_ _13013_/A hold290/X vssd1 vssd1 vccd1 vccd1 _13229_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _11897_/A _11897_/B _11896_/A vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11655__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07271__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11875_ _11726_/A _07150_/Y fanout4/X _11874_/Y vssd1 vssd1 vccd1 vccd1 _11948_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08520__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08520__B2 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ _10826_/A _10826_/B _10826_/C vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__and3_1
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10757_ _10757_/A _10757_/B vssd1 vssd1 vccd1 vccd1 _10771_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10688_/X sky130_fd_sc_hd__or2_1
X_12427_ _12484_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12429_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10137__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _12527_/B _12358_/B vssd1 vssd1 vccd1 vccd1 _12359_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07149__C _07152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__A1 _07075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12289_ _12290_/A _12290_/B _12290_/C vssd1 vssd1 vccd1 vccd1 _12289_/X sky130_fd_sc_hd__and3_1
XANTENNA__08339__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ _11193_/Y _11196_/B _11201_/A vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07446__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ instruction[1] _06850_/B instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06850_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_0_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06781_ _10914_/B _10914_/C _10917_/A vssd1 vssd1 vccd1 vccd1 _11023_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08520_ _08274_/A fanout93/X _10647_/A _08813_/A1 vssd1 vssd1 vccd1 vccd1 _08521_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08451_ _08449_/A _08449_/B _08450_/X vssd1 vssd1 vccd1 vccd1 _08477_/A sky130_fd_sc_hd__o21ba_1
X_07402_ _07403_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07402_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _08782_/A2 _10506_/A _10647_/A _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07333_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08275__B1 _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ reg1_val[28] reg1_val[29] _07263_/C _12639_/B _07128_/A vssd1 vssd1 vccd1
+ vccd1 _07265_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__xnor2_2
X_07195_ _07198_/A _07198_/B vssd1 vssd1 vccd1 vccd1 _07335_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_103_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07250__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07356__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _09905_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07075__B _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09836_/A _09836_/B _09836_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__nor3_1
X_06979_ _06979_/A _06979_/B _06979_/C vssd1 vssd1 vccd1 vccd1 _07065_/A sky130_fd_sc_hd__nand3_4
X_09767_ _09767_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09769_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09571__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11637__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ _09698_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__nor2_2
X_08718_ _08734_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _08751_/B sky130_fd_sc_hd__xnor2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07091__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08649_ _08678_/A _08648_/B _08628_/Y vssd1 vssd1 vccd1 vccd1 _08651_/B sky130_fd_sc_hd__a21oi_2
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11660_/A _11660_/B vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__nand2_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10860__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__A2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ _11677_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11593_/C sky130_fd_sc_hd__or2_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10611_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__or2_1
XFILLER_0_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ instruction[11] vssd1 vssd1 vccd1 vccd1 loadstore_dest[0] sky130_fd_sc_hd__buf_12
XFILLER_0_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10473_ _06704_/Y _10468_/Y _10470_/Y _10471_/X _10472_/X vssd1 vssd1 vccd1 vccd1
+ _10473_/X sky130_fd_sc_hd__o221a_1
X_12212_ _12256_/A _12212_/B vssd1 vssd1 vccd1 vccd1 _12214_/C sky130_fd_sc_hd__and2_1
X_13192_ _13230_/CLK _13192_/D vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ fanout9/A fanout7/X fanout6/X _12201_/A vssd1 vssd1 vccd1 vccd1 _12144_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _12068_/Y _12069_/X _12073_/X _12066_/X vssd1 vssd1 vccd1 vccd1 _12074_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07266__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09518__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _11238_/A _11024_/X _11023_/X vssd1 vssd1 vccd1 vccd1 _11026_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__11628__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ _12785_/X _12976_/B vssd1 vssd1 vccd1 vccd1 _12977_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11927_ hold220/A _11927_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11858_ _09501_/B _11625_/B _11858_/S vssd1 vssd1 vccd1 vccd1 _11858_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _10809_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
X_11789_ curr_PC[22] _11866_/C vssd1 vssd1 vccd1 vccd1 _11789_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_19 reg1_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07951_ _11470_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07982_/B sky130_fd_sc_hd__xnor2_2
X_06902_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__nand2b_4
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _07756_/A _07756_/C _07756_/B vssd1 vssd1 vccd1 vccd1 _07883_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06833_ _10331_/A _09501_/A _09336_/B _06833_/D vssd1 vssd1 vccd1 vccd1 _06834_/D
+ sky130_fd_sc_hd__and4_1
X_09621_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__or3_1
XANTENNA__07904__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06764_ _06700_/B _06762_/X _06763_/X vssd1 vssd1 vccd1 vccd1 _06764_/X sky130_fd_sc_hd__o21a_1
X_09552_ _10529_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__xnor2_1
X_08503_ _08503_/A _08503_/B vssd1 vssd1 vccd1 vccd1 _08561_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout255_A _07842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09102_/X _09106_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__mux2_1
X_06695_ _06763_/B _06613_/A _12553_/B _06694_/X vssd1 vssd1 vccd1 vccd1 _07296_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08434_ _08801_/A _08434_/B vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ _08366_/A _08366_/B vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07316_ _07569_/C _07316_/B vssd1 vssd1 vccd1 vccd1 _07327_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ _08607_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__xnor2_1
X_07247_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07249_/A sky130_fd_sc_hd__or2_1
XFILLER_0_5_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07178_ reg1_val[29] _07178_/B vssd1 vssd1 vccd1 vccd1 _07178_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__09212__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10505__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__B1_N _10315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ curr_PC[4] _09957_/C vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__nand2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _13099_/B _13100_/A _12735_/X vssd1 vssd1 vccd1 vccd1 _13104_/B sky130_fd_sc_hd__a21oi_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ hold62/X hold297/A vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12283__A1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ hold70/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__or2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11712_ curr_PC[21] _11712_/B vssd1 vssd1 vccd1 vccd1 _11866_/C sky130_fd_sc_hd__and2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11644_/B _11643_/B vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ _11574_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_107_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _11950_/A fanout43/X _08333_/B _12095_/A vssd1 vssd1 vccd1 vccd1 _10526_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13244_ _13246_/CLK _13244_/D vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
X_10456_ _06830_/C _10454_/X _10455_/Y vssd1 vssd1 vccd1 vccd1 _10456_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08380__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B1 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13246_/CLK _13175_/D vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12126_ hold265/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12184_/B sky130_fd_sc_hd__or2_1
X_10387_ _10537_/B _10387_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12057_ _11994_/A _11991_/Y _11993_/B vssd1 vssd1 vccd1 vccd1 _12061_/A sky130_fd_sc_hd__o21a_1
X_11008_ _11114_/A _11008_/B vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10150__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ hold56/X _12664_/A _12663_/B hold60/X rst vssd1 vssd1 vccd1 vccd1 hold61/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__08478__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10824__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__B _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__or2_1
XANTENNA__09978__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ reg1_val[24] _07263_/C _07128_/A vssd1 vssd1 vccd1 vccd1 _07102_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _08274_/A _11295_/B2 _08813_/A1 _11297_/A vssd1 vssd1 vccd1 vccd1 _08082_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ _07064_/A _07030_/X _07031_/X _07058_/B1 vssd1 vssd1 vccd1 vccd1 _12720_/A
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__08290__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08983_ _12053_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06964__B1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _08028_/A _08028_/B _07931_/Y vssd1 vssd1 vccd1 vccd1 _07955_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07865_ _09880_/B2 fanout43/X _07239_/A _10117_/A vssd1 vssd1 vccd1 vccd1 _07866_/B
+ sky130_fd_sc_hd__o22a_1
X_09604_ _09604_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09605_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06816_ _06805_/Y _06815_/X _12056_/A vssd1 vssd1 vccd1 vccd1 _12115_/C sky130_fd_sc_hd__a21o_1
X_07796_ _07797_/B _07858_/A _07797_/A vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__o21a_1
X_06747_ _06745_/Y _06747_/B vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__nand2b_2
X_09535_ _09406_/A _09406_/B _09404_/Y vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__a21oi_2
X_06678_ _06960_/A _10920_/A vssd1 vssd1 vccd1 vccd1 _11023_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09466_ _09617_/C _09465_/Y _10450_/A vssd1 vssd1 vccd1 vccd1 _09466_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10276__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12017__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _08417_/A _08417_/B vssd1 vssd1 vccd1 vccd1 _08423_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09681__A2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _06985_/A fanout63/X fanout55/X _06977_/A vssd1 vssd1 vccd1 vccd1 _09398_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _08336_/X _08337_/Y _08328_/Y _08332_/X vssd1 vssd1 vccd1 vccd1 _08349_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ _08280_/A _08280_/B _08280_/C vssd1 vssd1 vccd1 vccd1 _08283_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_22_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ _10310_/A _10311_/A _10311_/B _09777_/A vssd1 vssd1 vccd1 vccd1 _11163_/B
+ sky130_fd_sc_hd__or4b_2
X_11290_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__and2_1
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _12089_/A _10241_/B vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _10172_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10751__A1 _07277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout150 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _06985_/A sky130_fd_sc_hd__buf_6
Xfanout183 _09136_/Y vssd1 vssd1 vccd1 vccd1 _12073_/B2 sky130_fd_sc_hd__buf_2
Xfanout161 _07270_/Y vssd1 vssd1 vccd1 vccd1 _09428_/A sky130_fd_sc_hd__buf_8
Xfanout172 _09422_/A vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__buf_6
Xfanout194 _06925_/X vssd1 vssd1 vccd1 vccd1 _07058_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ hold283/A hold166/X vssd1 vssd1 vccd1 vccd1 _12814_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12744_ hold271/X hold19/X vssd1 vssd1 vccd1 vccd1 _13081_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12675_ _07099_/X _12731_/A2 hold73/X _13111_/A vssd1 vssd1 vccd1 vccd1 _13130_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11626_ _06628_/A _09501_/B _11625_/X _09138_/X vssd1 vssd1 vccd1 vccd1 _11626_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11557_ _11950_/A fanout14/X fanout52/X _12095_/A vssd1 vssd1 vccd1 vccd1 _11558_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _11462_/A fanout50/X _07988_/B fanout76/X vssd1 vssd1 vccd1 vccd1 _10509_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _11372_/A _11372_/B _11371_/A vssd1 vssd1 vccd1 vccd1 _11494_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ _13253_/CLK _13227_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
X_10439_ _10440_/B _10440_/A vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_20_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12731__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _13253_/CLK _13158_/D vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13089_ _13103_/A hold266/X vssd1 vssd1 vccd1 vccd1 _13249_/D sky130_fd_sc_hd__and2_1
X_12109_ _12107_/B _12045_/B _11909_/Y _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1
+ _12110_/D sky130_fd_sc_hd__o2111a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11298__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__B1 _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07650_/Y sky130_fd_sc_hd__nor2_1
X_06601_ reg1_val[23] _06601_/B vssd1 vssd1 vccd1 vccd1 _06798_/A sky130_fd_sc_hd__nand2_1
X_07581_ _09568_/A _07391_/B _09428_/A _12141_/A vssd1 vssd1 vccd1 vccd1 _07582_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07910__A2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06532_ instruction[1] _06850_/B instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06532_/X sky130_fd_sc_hd__or4bb_4
X_09320_ _09318_/X _09319_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09320_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10258__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A2 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _11183_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__xnor2_1
X_08202_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_8_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ _09183_/B _09182_/B vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _08737_/A2 fanout43/X _08333_/B _08733_/B1 vssd1 vssd1 vccd1 vccd1 _08134_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07629__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08101_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07015_/A _07015_/B vssd1 vssd1 vccd1 vccd1 _07015_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08926__A1 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__B2 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _07567_/A _07567_/B _07566_/A vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__o21ai_4
X_08897_ _08897_/A _08897_/B _08897_/C vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__and3_1
X_07917_ _07913_/A _07984_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07362__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ _07848_/A _07848_/B vssd1 vssd1 vccd1 vccd1 _07946_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10497__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07779_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07861_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _09880_/B2 _12141_/A fanout45/X _10117_/A vssd1 vssd1 vccd1 vccd1 _09519_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10249__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout33_A _12248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ _10790_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__and2_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09449_ _09275_/A _09275_/B _09273_/Y vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12496_/A _12460_/B vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12391_ reg1_val[11] curr_PC[11] _12444_/S vssd1 vssd1 vccd1 vccd1 _12393_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11412_/A _11412_/B _11412_/C vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__o21ai_1
X_11342_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08642__B _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12961__A2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08090__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__A1 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ _11468_/A _11273_/B vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10972__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ hold277/X _12663_/B _13011_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold278/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08917__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _11153_/A _10221_/X _10222_/X _10223_/Y vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10724__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__B2 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ fanout78/X fanout58/X fanout55/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _10156_/B
+ sky130_fd_sc_hd__o22a_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _10078_/Y _10079_/X _10085_/Y vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12229__A1 _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10989_/B sky130_fd_sc_hd__or2_1
X_12727_ _07075_/Y _12731_/A2 hold82/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13156_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ hold161/X hold164/X hold100/X vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11609_ _11521_/A _11519_/B _11535_/A vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12589_ reg1_val[18] _12615_/B vssd1 vssd1 vccd1 vccd1 _12591_/A sky130_fd_sc_hd__or2_1
XANTENNA__10412__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08081__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08821_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08820_/X sky130_fd_sc_hd__xor2_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09581__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06800__B _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__and2_1
X_07702_ _09979_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__xnor2_1
X_08682_ _08682_/A _08709_/A vssd1 vssd1 vccd1 vccd1 _08704_/A sky130_fd_sc_hd__xnor2_1
X_07633_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _07634_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout168_A _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _07565_/A _07565_/B _07565_/C vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09303_ _09301_/X _09302_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__mux2_1
X_07495_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06515_ reg1_val[16] vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09234_ _09233_/B _09233_/C _09233_/A vssd1 vssd1 vccd1 vccd1 _09235_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _11033_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08116_ _08274_/A fanout76/X _11462_/A _08813_/A1 vssd1 vssd1 vccd1 vccd1 _08117_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__07359__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ _09080_/X _09095_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09129_/B sky130_fd_sc_hd__mux2_1
X_08047_ _08607_/A _08047_/B vssd1 vssd1 vccd1 vccd1 _08050_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10706__A1 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06710__B _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _10156_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__xor2_4
X_08949_ _10876_/A1 fanout36/X fanout34/X _10490_/B2 vssd1 vssd1 vccd1 vccd1 _08950_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11960_ _11961_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__and2_1
XANTENNA__08918__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _11230_/C _10909_/X _10910_/Y vssd1 vssd1 vccd1 vccd1 _10911_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _11892_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10842_ _12086_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10844_/B sky130_fd_sc_hd__xnor2_1
X_10773_ _10617_/A _10617_/B _10616_/A vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ reg1_val[3] _12512_/B vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _12448_/B _12443_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XFILLER_0_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _12375_/A _12375_/B _12375_/C vssd1 vssd1 vccd1 vccd1 _12382_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07269__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _11327_/A _11327_/B _11327_/C vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11256_ _06978_/B _12280_/A _09147_/X _06660_/Y vssd1 vssd1 vccd1 vccd1 _11256_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06901__A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ hold213/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10465_/C sky130_fd_sc_hd__or2_1
X_11187_ _11187_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11189_/C sky130_fd_sc_hd__and2_1
X_10138_ _10139_/A _10139_/B vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__nand2b_1
X_10069_ _09483_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10069_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09866__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09659__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07280_ _09979_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07294_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12085__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold225 hold237/X vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _11983_/A _09018_/A _09018_/B _12179_/A vssd1 vssd1 vccd1 vccd1 _09922_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__B _12532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__xor2_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09017_/A _09781_/X _09782_/Y vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__o21a_1
X_08803_ _08804_/A _08803_/B _08803_/C vssd1 vssd1 vccd1 vccd1 _08803_/X sky130_fd_sc_hd__or3_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13102__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ _10252_/A _06996_/B vssd1 vssd1 vccd1 vccd1 _06999_/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__xnor2_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__B1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _08665_/A vssd1 vssd1 vccd1 vccd1 _08685_/B sky130_fd_sc_hd__inv_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07616_ _07616_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11164__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _08699_/A2 _08737_/A2 _08813_/B1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 _08597_/B
+ sky130_fd_sc_hd__o22a_1
X_07547_ _07661_/A _07547_/B vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07096__A2 _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09221_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06705__B _06931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _09148_/A instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09148_/X
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _09075_/X _09078_/X _09633_/S vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _11110_/A _11110_/B vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__xnor2_1
X_12090_ _12090_/A vssd1 vssd1 vccd1 vccd1 _12092_/B sky130_fd_sc_hd__inv_2
X_11041_ _11620_/B _11140_/B hold171/A vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10155__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ hold289/X _12663_/B _12991_/X _12664_/A vssd1 vssd1 vccd1 vccd1 hold290/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11943_ _06847_/X _11940_/X _12079_/C _11942_/Y vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__11655__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ _07152_/X fanout4/X _11726_/A vssd1 vssd1 vccd1 vccd1 _11874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08520__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _07278_/A _12280_/A _10824_/X _06687_/B vssd1 vssd1 vccd1 vccd1 _10826_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_55_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08383__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _10756_/A _10756_/B vssd1 vssd1 vccd1 vccd1 _10757_/B sky130_fd_sc_hd__or2_1
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10418__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ _10449_/A _09027_/A _09027_/B _12179_/A vssd1 vssd1 vccd1 vccd1 _10688_/B
+ sky130_fd_sc_hd__a31o_1
X_12426_ reg1_val[16] curr_PC[16] _12444_/S vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _12527_/B _12358_/B vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__A2 _07075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _12288_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12290_/C sky130_fd_sc_hd__xnor2_2
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__nand2_1
X_11239_ _11124_/A _11237_/Y _11238_/Y vssd1 vssd1 vccd1 vccd1 _11240_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__08339__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ _06690_/Y _06779_/X _06831_/D vssd1 vssd1 vccd1 vccd1 _10914_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__07462__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _08500_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08450_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07401_ _07366_/A _07366_/B _07369_/A vssd1 vssd1 vccd1 vccd1 _07403_/B sky130_fd_sc_hd__o21ai_2
X_08381_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08404_/A sky130_fd_sc_hd__or2_1
X_07332_ _07332_/A _07332_/B vssd1 vssd1 vccd1 vccd1 _07333_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12527__B _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07263_ reg1_val[28] reg1_val[29] _07263_/C _12639_/B vssd1 vssd1 vccd1 vccd1 _07574_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07194_ _08276_/A _07194_/B vssd1 vssd1 vccd1 vccd1 _07198_/B sky130_fd_sc_hd__xnor2_2
X_09002_ _09002_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _10913_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout200_A _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07250__A2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _09760_/A _09760_/B _09758_/Y vssd1 vssd1 vccd1 vccd1 _09905_/B sky130_fd_sc_hd__a21boi_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _09836_/A _09836_/B _09836_/C vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__o21a_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06978_ _06978_/A _06978_/B vssd1 vssd1 vccd1 vccd1 _06979_/C sky130_fd_sc_hd__nor2_1
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09767_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11637__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ _08219_/B _08733_/B1 _08735_/A2 _08815_/B vssd1 vssd1 vccd1 vccd1 _08718_/B
+ sky130_fd_sc_hd__o22a_1
X_09697_ _09697_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07091__B _07091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ _08628_/Y _08648_/B vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__nand2b_1
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12718__A _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08579_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08626_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10610_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10238__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ _10408_/B _10425_/B _10406_/X vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__a21oi_1
X_13260_ _13260_/CLK hold160/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10472_ _07289_/A _06905_/Y _11625_/B _06706_/B _12080_/A vssd1 vssd1 vccd1 vccd1
+ _10472_/X sky130_fd_sc_hd__o221a_1
X_12211_ _12211_/A _12211_/B _12211_/C vssd1 vssd1 vccd1 vccd1 _12212_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _13230_/CLK _13191_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07777__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _12142_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__xnor2_1
X_12073_ _09293_/A _09940_/X _09952_/X _12073_/B2 _12072_/Y vssd1 vssd1 vccd1 vccd1
+ _12073_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07266__B _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B2 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__A1 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ _10917_/A _10915_/X _10933_/A vssd1 vssd1 vccd1 vccd1 _11024_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08378__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ _13111_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _13225_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13254_/CLK sky130_fd_sc_hd__clkbuf_8
X_11926_ _12302_/A _10218_/Y _11925_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07701__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ _11857_/A _11857_/B vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _09790_/X _09792_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _07028_/B _12280_/A _06907_/A _11787_/X vssd1 vssd1 vccd1 vccd1 _11788_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10739_ _11295_/B2 fanout52/X _11297_/A fanout14/X vssd1 vssd1 vccd1 vccd1 _10740_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13002__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _12410_/A _12410_/B _12410_/C vssd1 vssd1 vccd1 vccd1 _12417_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07950_ _08782_/B2 fanout41/X _08135_/B _09428_/A vssd1 vssd1 vccd1 vccd1 _07951_/B
+ sky130_fd_sc_hd__o22a_1
X_06901_ _12080_/A _06901_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07881_ _07879_/A _07879_/B _07880_/Y vssd1 vssd1 vccd1 vccd1 _07889_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06832_ _06832_/A _09926_/A vssd1 vssd1 vccd1 vccd1 _06834_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08288__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _11983_/A _10321_/A _09917_/B _09619_/Y _09061_/X vssd1 vssd1 vccd1 vccd1
+ _09620_/Y sky130_fd_sc_hd__a311oi_1
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07192__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ reg2_val[0] _06763_/B vssd1 vssd1 vccd1 vccd1 _06763_/X sky130_fd_sc_hd__or2_2
X_09551_ fanout82/X fanout68/X fanout65/X _06940_/A vssd1 vssd1 vccd1 vccd1 _09552_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08502_ _08502_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__or2_1
X_09482_ _09099_/X _09125_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09482_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06694_ reg2_val[10] _06748_/B vssd1 vssd1 vccd1 vccd1 _06694_/X sky130_fd_sc_hd__and2_1
XFILLER_0_53_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_A _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ _08782_/A2 _09180_/B2 _10506_/A _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08434_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ _08362_/A _08362_/B _08363_/X vssd1 vssd1 vccd1 vccd1 _08366_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07315_ _07315_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07316_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ _08642_/B _08715_/A2 _08735_/B1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 _08296_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07246_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09847__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07177_ reg1_val[28] _07263_/C _12639_/B _07128_/A vssd1 vssd1 vccd1 vccd1 _07178_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10505__B _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09818_ _09780_/Y _09817_/X _11713_/A vssd1 vssd1 vccd1 vccd1 _09818_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout63_A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _09749_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__xnor2_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ hold273/A hold47/X vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__nand2b_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ hold15/X _12692_/B _12690_/Y _13013_/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ curr_PC[21] _11712_/B vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ _12086_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11573_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08661__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10524_ _10374_/A _10373_/B _10371_/X vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13243_ _13243_/CLK _13243_/D vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
X_10455_ _06830_/C _10454_/X _09498_/A vssd1 vssd1 vccd1 vccd1 _10455_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _13246_/CLK hold173/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10349__A2 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07277__A _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12125_ _09815_/X _12124_/Y _12125_/S vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__mux2_1
X_10386_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__and2_1
XFILLER_0_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _12056_/A _12056_/B vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__or2_1
X_11007_ _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11008_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _12142_/A _12686_/B hold57/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12274__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09675__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ hold235/A _13084_/B2 _13084_/A2 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__A _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ _11909_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11909_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11234__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _10920_/A _07091_/B _07091_/C _07091_/D _07128_/A vssd1 vssd1 vccd1 vccd1
+ _07148_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07989__B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__B2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08080_ _08240_/A _08240_/B _08078_/A vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08571__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07065_/A _07065_/B _07065_/C _07064_/A vssd1 vssd1 vccd1 vccd1 _07031_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10606__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07187__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06964__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06964__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ _08982_/A _09461_/A vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _07933_/A _07933_/B vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout198_A _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _08916_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07868_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06815_ _06806_/Y _06814_/X _11988_/A vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__a21o_1
X_09603_ _09603_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__xnor2_2
X_07795_ _07857_/A _07857_/B vssd1 vssd1 vccd1 vccd1 _07858_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_64_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06746_ reg1_val[3] _07099_/A vssd1 vssd1 vccd1 vccd1 _06747_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09534_ _09534_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__nand2_1
X_06677_ _06763_/B _06613_/A _12571_/B _06676_/X vssd1 vssd1 vccd1 vccd1 _06960_/A
+ sky130_fd_sc_hd__a31o_4
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09465_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10276__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10276__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08416_ _08416_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08423_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09396_ _09396_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09418__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08410_/A _08410_/B _08343_/X vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _08734_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08280_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08481__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ _08916_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07243_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ fanout44/X fanout92/X _12690_/A fanout11/X vssd1 vssd1 vccd1 vccd1 _10241_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10171_ _10171_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__xnor2_2
Xfanout140 _09880_/B2 vssd1 vssd1 vccd1 vccd1 _08735_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__10751__A2 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout151 _06984_/Y vssd1 vssd1 vccd1 vccd1 _08699_/A2 sky130_fd_sc_hd__buf_8
Xfanout173 _07040_/X vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__buf_8
Xfanout162 _09237_/A vssd1 vssd1 vccd1 vccd1 _08782_/B2 sky130_fd_sc_hd__buf_6
Xfanout195 _12926_/A2 vssd1 vssd1 vccd1 vccd1 _12962_/B2 sky130_fd_sc_hd__buf_4
Xfanout184 _09293_/A vssd1 vssd1 vccd1 vccd1 _09120_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12812_ _13054_/B _13055_/A _12752_/X vssd1 vssd1 vccd1 vccd1 _13059_/A sky130_fd_sc_hd__a21o_1
X_12743_ hold19/X hold271/X vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11082__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ hold72/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__or2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10019__A1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__B1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11625_ _11625_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06904__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _11662_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11560_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _10507_/A _10507_/B vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13226_ _13253_/CLK _13226_/D vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11487_ _11395_/A _11395_/B _11394_/A vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__xnor2_1
X_13157_ _13254_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10484_/B _10369_/B vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__and2_1
X_13088_ hold265/X _06858_/B _13087_/X _13110_/A2 vssd1 vssd1 vccd1 vccd1 hold266/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06946__B2 _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _12160_/B _12108_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__xnor2_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ _12040_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08699__A1 _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06600_ reg2_val[23] _06754_/B _06657_/B1 _06598_/X vssd1 vssd1 vccd1 vccd1 _07028_/A
+ sky130_fd_sc_hd__a22o_2
X_07580_ _07260_/A _07260_/B _07258_/Y vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__a21oi_2
X_06531_ instruction[1] _06850_/B instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06863_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__11455__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10258__A1 _10377_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _10490_/B2 fanout36/X fanout34/X fanout80/X vssd1 vssd1 vccd1 vccd1 _09251_/B
+ sky130_fd_sc_hd__o22a_1
X_08201_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09181_ _11726_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ _08146_/A _08146_/B _08121_/X vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08063_ _08741_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08065_/B sky130_fd_sc_hd__xnor2_1
X_07014_ _07028_/B _07014_/B vssd1 vssd1 vccd1 vccd1 _07014_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__06533__B _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout113_A _11887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__A2 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08926__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _07641_/A _07640_/A _07640_/B _07644_/A vssd1 vssd1 vccd1 vccd1 _08975_/A
+ sky130_fd_sc_hd__o31ai_2
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07927_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11167__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ _08897_/A _08897_/B _08897_/C vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__a21oi_1
X_07847_ _07847_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10497__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__B2 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__B2 _07110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__A2 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _10126_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06729_ reg2_val[5] _06700_/B _12271_/S vssd1 vssd1 vccd1 vccd1 _06928_/C sky130_fd_sc_hd__a21o_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10249__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ _09427_/A _09427_/B _09425_/Y vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__o21ai_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout26_A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ _09448_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__xor2_1
X_12390_ _12396_/B _12390_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11410_ _11506_/A _11410_/B vssd1 vssd1 vccd1 vccd1 _11412_/C sky130_fd_sc_hd__and2_1
XANTENNA__09811__B1 _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _11246_/A _11243_/Y _11245_/B vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08090__A2 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11272_ fanout9/X fanout36/X fanout34/X fanout3/X vssd1 vssd1 vccd1 vccd1 _11273_/B
+ sky130_fd_sc_hd__o22a_1
X_13011_ hold255/X _13010_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08917__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ curr_PC[7] _10354_/C _11153_/A vssd1 vssd1 vccd1 vccd1 _10223_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10185__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _10154_/A _10154_/B vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__xor2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _06832_/A _09141_/Y _10084_/X vssd1 vssd1 vccd1 vccd1 _10085_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06618__B _06987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10989_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ hold81/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__or2_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ hold164/X hold100/X vssd1 vssd1 vccd1 vccd1 _12657_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ _11838_/A _11608_/B _11608_/C vssd1 vssd1 vccd1 vccd1 _11608_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _12588_/A _12592_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
XANTENNA__10412__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _11533_/Y _11534_/X _11538_/X vssd1 vssd1 vccd1 vccd1 _11539_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__08081__A2 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10156__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10412__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09664__B _09664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ _13217_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 _13209_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12371__A _12537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09581__A2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__B _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08744_/A _08743_/C _08743_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__a21o_1
X_07701_ _07137_/Y fanout43/X _08333_/B _12686_/A vssd1 vssd1 vccd1 vccd1 _07702_/B
+ sky130_fd_sc_hd__o22a_1
X_08681_ _08681_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08706_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10479__B2 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__and2_1
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08296__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _09082_/X _09084_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09302_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07565_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06514_ reg1_val[4] vssd1 vssd1 vccd1 vccd1 _07051_/A sky130_fd_sc_hd__inv_2
XFILLER_0_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07494_ _10156_/A _07494_/B vssd1 vssd1 vccd1 vccd1 _07495_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06855__B1 _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _09233_/A _09233_/B _09233_/C vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__and3_1
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13260_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ _09162_/X _09164_/B vssd1 vssd1 vccd1 vccd1 _09166_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10939__C1 _10936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ _08801_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__xnor2_4
X_09095_ _09094_/X _09087_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09095_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10875__A_N _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ _08606_/A2 _08689_/B1 _09180_/B2 _08642_/B vssd1 vssd1 vccd1 vccd1 _08047_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ fanout78/X fanout64/X fanout58/X _10852_/B2 vssd1 vssd1 vccd1 vccd1 _09998_/B
+ sky130_fd_sc_hd__o22a_2
X_08948_ _11796_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _08952_/A sky130_fd_sc_hd__xnor2_1
X_08879_ _08985_/A _08985_/B _08880_/B vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _11230_/C _10909_/X _09061_/X vssd1 vssd1 vccd1 vccd1 _10910_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06689__A3 _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _11964_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__or2_1
XANTENNA__06744__A_N _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _11295_/B2 fanout14/X fanout52/X _11462_/A vssd1 vssd1 vccd1 vccd1 _10842_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _10658_/A _10658_/B _10659_/X vssd1 vssd1 vccd1 vccd1 _10783_/A sky130_fd_sc_hd__o21ba_1
X_12511_ reg1_val[3] _12512_/B vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13051__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12454_/A _12454_/B _12455_/B vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08599__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12382_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12375_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07269__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11324_ _11324_/A _11324_/B vssd1 vssd1 vccd1 vccd1 _11327_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ _06660_/Y _09501_/B _09138_/X vssd1 vssd1 vccd1 vccd1 _11255_/Y sky130_fd_sc_hd__o21ai_1
X_10206_ _12125_/S _10204_/A _10205_/X _09156_/B vssd1 vssd1 vccd1 vccd1 _10220_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07285__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11187_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__nor2_1
X_10137_ _11799_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10139_/B sky130_fd_sc_hd__xor2_1
X_10068_ _09476_/X _09479_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _10068_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12083__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ _11649_/A _12731_/A2 hold167/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13147_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10397__B1 _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09920_ _11983_/A _09018_/B _09018_/A vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12689__A2 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10149__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__xor2_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ reg1_val[10] _06994_/B vssd1 vssd1 vccd1 vccd1 _06996_/B sky130_fd_sc_hd__xor2_1
X_09782_ _09017_/A _09781_/X _12179_/A vssd1 vssd1 vccd1 vccd1 _09782_/Y sky130_fd_sc_hd__a21oi_1
X_08802_ _08803_/B _08803_/C vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__nor2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08733_ _08219_/B _08737_/A2 _08733_/B1 _08815_/B vssd1 vssd1 vccd1 vccd1 _08734_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08664_ _08734_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__xnor2_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _07615_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11164__B _11164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _08801_/A _08595_/B vssd1 vssd1 vccd1 vccd1 _08601_/A sky130_fd_sc_hd__xnor2_1
X_07546_ _07546_/A _07546_/B _07546_/C vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07477_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _09217_/B vssd1 vssd1 vccd1 vccd1 _09216_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09147_ instruction[4] instruction[6] instruction[5] instruction[3] vssd1 vssd1 vccd1
+ vccd1 _09147_/X sky130_fd_sc_hd__and4bb_4
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _09076_/X _09077_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09078_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _08031_/A _08031_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07005__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ hold216/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11140_/B sky130_fd_sc_hd__or2_1
XANTENNA__07556__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B2 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ hold285/X _12990_/Y hold246/X vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12301__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ curr_PC[24] _11941_/B _11636_/S vssd1 vssd1 vccd1 vccd1 _11942_/Y sky130_fd_sc_hd__o21ai_1
X_11873_ _11873_/A _11873_/B vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12065__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10824_ _10823_/A _09141_/Y _10823_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _10824_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ _10756_/A _10756_/B vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10686_ _10449_/A _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__a21oi_1
X_12425_ _12429_/B _12425_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XANTENNA__10379__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ reg1_val[6] curr_PC[6] _12444_/S vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07244__B1 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ _11168_/A _11168_/B _11171_/A vssd1 vssd1 vccd1 vccd1 _11314_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ _12029_/B fanout4/X _12250_/B vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11238_ _11238_/A _11238_/B _11238_/C vssd1 vssd1 vccd1 vccd1 _11238_/Y sky130_fd_sc_hd__nand3_1
X_11169_ _11169_/A _11296_/A _11169_/C vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__or3_1
XFILLER_0_93_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07400_ _07343_/A _07343_/B _07340_/X vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__o21a_1
X_08380_ _10853_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07331_ _07332_/A _07332_/B vssd1 vssd1 vccd1 vccd1 _07333_/A sky130_fd_sc_hd__and2_1
XFILLER_0_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10609__A _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _07262_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _07275_/A sky130_fd_sc_hd__xnor2_1
X_07193_ _07044_/Y _08384_/B _07069_/X _12499_/A vssd1 vssd1 vccd1 vccd1 _07194_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ _09001_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _09903_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__xnor2_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09834_ _09834_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09836_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08735__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06977_ _06977_/A vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__inv_2
X_09765_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__and2_1
XANTENNA__11175__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _08814_/A _08716_/B vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__xnor2_1
X_09696_ _09697_/B _09697_/A vssd1 vssd1 vccd1 vccd1 _09836_/B sky130_fd_sc_hd__and2b_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _08647_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__nand2_1
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__A1 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__B2 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08578_/A vssd1 vssd1 vccd1 vccd1 _08626_/A sky130_fd_sc_hd__inv_2
XANTENNA__08484__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__B _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07529_ _09420_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07758_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ _10540_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__xor2_1
X_10471_ hold255/A _09808_/B _10588_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ _12211_/A _12211_/B _12211_/C vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ _13254_/CLK hold130/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07777__A1 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__B2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _12141_/A fanout4/X vssd1 vssd1 vccd1 vccd1 _12142_/B sky130_fd_sc_hd__nor2_1
X_12072_ _06552_/B _12070_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12072_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09518__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _11238_/A _11023_/B _11023_/C vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__and3_1
XANTENNA__08659__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__B1 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12974_ hold296/X _12663_/B _12973_/X _12664_/A vssd1 vssd1 vccd1 vccd1 _12975_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11925_ _12302_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__B2 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A1 _07137_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ hold220/A _11620_/B _11927_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _11857_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10807_/Y sky130_fd_sc_hd__nand2_1
X_11787_ _11761_/Y _11762_/X _11763_/X _11764_/Y _11786_/X vssd1 vssd1 vccd1 vccd1
+ _11787_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__B2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ _10738_/A _10738_/B vssd1 vssd1 vccd1 vccd1 _10749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13002__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _12417_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12410_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10669_ _10669_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12339_ _12340_/A _12340_/B _12340_/C vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06900_ _09495_/A is_load _06613_/A _06897_/X vssd1 vssd1 vccd1 vccd1 _06901_/B sky130_fd_sc_hd__a22o_2
XANTENNA__08717__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _07902_/B _07902_/A vssd1 vssd1 vccd1 vccd1 _07880_/Y sky130_fd_sc_hd__nand2b_1
X_06831_ _06831_/A _11026_/A _10917_/A _06831_/D vssd1 vssd1 vccd1 vccd1 _06835_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__12277__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ _06512_/Y _06532_/X _06535_/Y _12502_/B vssd1 vssd1 vccd1 vccd1 _06762_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09550_ _09550_/A _09550_/B vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__xnor2_2
X_09481_ _09477_/X _09480_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08501_ _08501_/A vssd1 vssd1 vccd1 vccd1 _08561_/A sky130_fd_sc_hd__inv_2
X_06693_ _10706_/S _06693_/B vssd1 vssd1 vccd1 vccd1 _10692_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _08497_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08452_/A sky130_fd_sc_hd__or2_1
XFILLER_0_86_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ _08419_/B _08419_/A vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07314_ _07315_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07569_/C sky130_fd_sc_hd__nor2_1
X_08294_ _08272_/X _08353_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08294_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__A2 _10447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ _10156_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07248_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07176_ reg1_val[26] reg1_val[27] _07176_/C vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__or3_4
XFILLER_0_42_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _11124_/A vssd1 vssd1 vccd1 vccd1 _12263_/S sky130_fd_sc_hd__buf_4
XANTENNA__10515__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A _09817_/B _09817_/C _09816_/X vssd1 vssd1 vccd1 vccd1 _09817_/X
+ sky130_fd_sc_hd__or4b_1
X_09748_ _09748_/A _09748_/B vssd1 vssd1 vccd1 vccd1 _09749_/B sky130_fd_sc_hd__xor2_2
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09133__B1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ _06987_/A _12280_/A _06907_/A _11709_/X vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__a22o_1
X_09679_ _11726_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__xor2_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12690_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _12690_/Y sky130_fd_sc_hd__nand2_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ fanout63/X fanout15/X _07513_/B fanout60/X vssd1 vssd1 vccd1 vccd1 _11642_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11572_/Y sky130_fd_sc_hd__nand2_1
X_10523_ _10523_/A _10523_/B vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _13243_/CLK _13242_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10454_ _06775_/Y _10453_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09739__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13243_/CLK _13173_/D vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08947__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _12124_/A _12124_/B vssd1 vssd1 vccd1 vccd1 _12124_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12055_ _12056_/A _12056_/B vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07293__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _06508_/Y _12664_/A _12663_/B hold56/X rst vssd1 vssd1 vccd1 vccd1 hold57/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09675__B2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12888_ _13080_/A hold236/X vssd1 vssd1 vccd1 vccd1 _13185_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07686__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ _11873_/A _11873_/B _11907_/Y vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_114_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ _11838_/A _11838_/C _11838_/B vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09978__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07989__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ _07065_/A _07065_/B _07065_/C _07058_/B1 vssd1 vssd1 vccd1 vccd1 _07030_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07187__B _07187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06964__A2 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_11_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07932_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _08028_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11718__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ fanout82/X _12688_/A _12690_/A _06939_/X vssd1 vssd1 vccd1 vccd1 _07864_/B
+ sky130_fd_sc_hd__o22a_1
X_06814_ _06798_/A _06798_/B _11918_/A vssd1 vssd1 vccd1 vccd1 _06814_/X sky130_fd_sc_hd__a21o_1
X_09602_ _09600_/A _09600_/B _09603_/B vssd1 vssd1 vccd1 vccd1 _09602_/Y sky130_fd_sc_hd__a21oi_1
X_07794_ _11468_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07857_/B sky130_fd_sc_hd__xnor2_1
X_09533_ _09412_/A _09411_/Y _09417_/A vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__a21o_1
X_06745_ reg1_val[3] _07099_/A vssd1 vssd1 vccd1 vccd1 _06745_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout260_A _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ reg2_val[13] _06748_/B vssd1 vssd1 vccd1 vccd1 _06676_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _09464_/A _10320_/A _09617_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10276__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _08412_/A _08475_/A _08414_/X _08416_/A vssd1 vssd1 vccd1 vccd1 _08427_/B
+ sky130_fd_sc_hd__o211ai_2
X_09395_ _09395_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09418__A1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__A3 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ _08535_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__B2 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08277_ _12694_/A _08219_/B _09222_/B2 _10957_/A vssd1 vssd1 vccd1 vccd1 _08278_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07228_ _08565_/B _12704_/A _12702_/A fanout82/X vssd1 vssd1 vccd1 vccd1 _07229_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12725__A1 _07069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _07147_/Y _07154_/X _07799_/B _07157_/X vssd1 vssd1 vccd1 vccd1 _07160_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _10168_/A _10168_/B _10171_/B vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__a21o_1
Xfanout130 _08565_/B vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__clkbuf_8
Xfanout152 _08670_/A2 vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__buf_6
Xfanout141 _07158_/Y vssd1 vssd1 vccd1 vccd1 _09880_/B2 sky130_fd_sc_hd__buf_8
Xfanout163 _07186_/Y vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__buf_8
Xfanout174 _09725_/B2 vssd1 vssd1 vccd1 vccd1 _08755_/B sky130_fd_sc_hd__buf_6
Xfanout196 _12731_/A2 vssd1 vssd1 vccd1 vccd1 _12926_/A2 sky130_fd_sc_hd__buf_2
Xfanout185 _09293_/A vssd1 vssd1 vccd1 vccd1 _09124_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__11161__B1 _11157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__B _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12811_ _13049_/A _13050_/A _13049_/B vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ _12740_/X _12742_/B vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _07271_/X _12962_/B2 hold77/X _12970_/A vssd1 vssd1 vccd1 vccd1 _13129_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09409__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ _11623_/B _11698_/B hold263/A vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11555_ _11554_/B _11555_/B vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11486_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__and2_1
X_10506_ _10506_/A _11296_/A _10507_/A vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or3_1
X_13225_ _13253_/CLK _13225_/D vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
X_10437_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__and2_1
XANTENNA__12192__A2 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _13251_/CLK _13156_/D vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06920__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10368_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10369_/B sky130_fd_sc_hd__or2_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13087_ hold299/A _13086_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__mux2_1
X_12107_ _12107_/A _12107_/B vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__nor2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10300_/B _10300_/A vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09345__B1 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _11970_/A _11970_/B _11969_/A vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08699__A2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _06530_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11273__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10258__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _12684_/A _07153_/X fanout47/X _09180_/B2 vssd1 vssd1 vccd1 vccd1 _09181_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08146_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_16_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07831__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ _10876_/A1 _08755_/B fanout93/X _08740_/A2 vssd1 vssd1 vccd1 vccd1 _08063_/B
+ sky130_fd_sc_hd__o22a_1
X_07013_ _07065_/A _07028_/C _07028_/D _07303_/A vssd1 vssd1 vccd1 vccd1 _07014_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout106_A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ _08964_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _08977_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07915_ _12668_/A fanout51/X fanout49/X _08782_/B2 vssd1 vssd1 vccd1 vccd1 _07916_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12978__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A0 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08897_/C sky130_fd_sc_hd__or2_1
XANTENNA__06976__S _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ fanout77/X _07040_/X _07041_/Y _12710_/A vssd1 vssd1 vccd1 vccd1 _07847_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10497__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _12704_/A _09725_/B2 _12702_/A _10009_/A vssd1 vssd1 vccd1 vccd1 _07778_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06728_ reg2_val[5] _06700_/B _12271_/S vssd1 vssd1 vccd1 vccd1 _06730_/B sky130_fd_sc_hd__a21oi_2
X_09516_ _09450_/A _09450_/B _09451_/Y vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10249__A2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09447_ _09447_/A _09447_/B vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06659_ _07233_/A _06978_/B vssd1 vssd1 vccd1 vccd1 _06785_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12726__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__A1 _06737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12946__A1 _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _08740_/A2 _09180_/B2 _10506_/A _08755_/B vssd1 vssd1 vccd1 vccd1 _08330_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout19_A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06724__B _07158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _11339_/A _11339_/B _09498_/A vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ _13010_/A _13010_/B vssd1 vssd1 vccd1 vccd1 _13010_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11271_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ curr_PC[7] _10354_/C vssd1 vssd1 vccd1 vccd1 _10222_/X sky130_fd_sc_hd__or2_1
XANTENNA__10185__A1 _10447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10154_/A _10154_/B vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__nand2b_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_10084_ _06723_/Y _09138_/X _11625_/B _06725_/B _10083_/X vssd1 vssd1 vccd1 vccd1
+ _10084_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _10986_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12725_ _07069_/X _12731_/A2 hold50/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13155_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09498__A _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ _12656_/A _12656_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
XANTENNA__06915__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _11838_/A _11608_/B _11608_/C vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__a21o_1
X_12587_ reg1_val[17] _12615_/B vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06634__B _06980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10412__A2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ _09293_/A _10810_/Y _11531_/X _11537_/X vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11469_ fanout9/A fanout41/X _08135_/B fanout3/X vssd1 vssd1 vccd1 vccd1 _11470_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _13208_/CLK _13208_/D vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _13251_/CLK _13139_/D vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11373__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__C _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__nand2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08680_ _08680_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__xnor2_2
X_07631_ _07875_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _07633_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07562_ _11955_/A _07562_/B vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__xnor2_2
X_06513_ reg1_val[1] vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__inv_2
XFILLER_0_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09301_ _09081_/X _09108_/X _09309_/S vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__mux2_1
X_07493_ _10852_/B2 fanout92/X _07304_/Y fanout78/X vssd1 vssd1 vccd1 vccd1 _07494_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ _09432_/A _09231_/B _09223_/Y vssd1 vssd1 vccd1 vccd1 _09233_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12928__A1 _06961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _10073_/S _09165_/B vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11450__B _11450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12546__B _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08057__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06696__A_N _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ fanout81/X _08782_/A2 _08756_/B2 _11169_/A vssd1 vssd1 vccd1 vccd1 _08115_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _09090_/X _09093_/X _09479_/S vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08045_ _09055_/A _08988_/A vssd1 vssd1 vccd1 vccd1 _08045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09557__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09996_ _10607_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__xor2_4
X_08947_ fanout51/X _09180_/B2 _10506_/A fanout49/X vssd1 vssd1 vccd1 vccd1 _08948_/B
+ sky130_fd_sc_hd__o22a_1
X_08878_ _07897_/Y _08986_/B _09057_/B _08876_/Y _08877_/A vssd1 vssd1 vccd1 vccd1
+ _08985_/B sky130_fd_sc_hd__a311o_4
XANTENNA__07391__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11625__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07829_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11419__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _10840_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _10771_/A _10771_/B vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _12509_/A _12506_/Y _12508_/B vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_54_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12441_ _12454_/B _12455_/B _12454_/A vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08048__B1 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08599__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ _12537_/B _12372_/B vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08950__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ _11324_/B _11324_/A vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ hold253/A _12000_/A2 _11354_/B _11253_/Y _12313_/A1 vssd1 vssd1 vccd1 vccd1
+ _11254_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ _12302_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10205_/X sky130_fd_sc_hd__or2_1
XANTENNA__08220__B1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__B _07286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ _07237_/A fanout3/X _11184_/X _11271_/A vssd1 vssd1 vccd1 vccd1 _11187_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _08384_/A _07154_/X _07799_/B _11091_/A vssd1 vssd1 vccd1 vccd1 _10137_/B
+ sky130_fd_sc_hd__a22o_1
X_10067_ _10067_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10067_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11535__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__B1 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12083__B2 _12148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__A1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10969_ _11950_/A fanout41/X _08135_/B _12095_/A vssd1 vssd1 vccd1 vccd1 _10970_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ hold166/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__or2_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11551__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__B1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12639_ _12656_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09787__B1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 hold216/X vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10149__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__nor2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _07050_/A _06993_/B vssd1 vssd1 vccd1 vccd1 _06994_/B sky130_fd_sc_hd__nand2_1
X_09781_ _11983_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__and2_1
X_08801_ _08801_/A _08810_/A vssd1 vssd1 vccd1 vccd1 _08803_/C sky130_fd_sc_hd__and2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11726__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ _08732_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__xnor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__A2 _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _08815_/B _08715_/A2 _08735_/B1 _08219_/B vssd1 vssd1 vccd1 vccd1 _08664_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout173_A _07040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ _10529_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07616_/B sky130_fd_sc_hd__xnor2_1
X_08594_ _08756_/B2 _08715_/A2 _08735_/B1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 _08595_/B
+ sky130_fd_sc_hd__o22a_1
X_07545_ _07543_/A _07543_/B _07746_/A vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__09630__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09215_ _10529_/A _09215_/B vssd1 vssd1 vccd1 vccd1 _09217_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ _09146_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__or2_2
XANTENNA__08770__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ reg1_val[4] reg1_val[27] _09092_/S vssd1 vssd1 vccd1 vccd1 _09077_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08028_ _08028_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08031_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_A _11235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A2 _07137_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _09979_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__xnor2_1
X_12990_ _12990_/A _12990_/B vssd1 vssd1 vccd1 vccd1 _12990_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ curr_PC[24] _11941_/B vssd1 vssd1 vccd1 vccd1 _12079_/C sky130_fd_sc_hd__and2_2
X_11872_ _11678_/B _11757_/Y _11869_/Y _11871_/Y _11869_/C vssd1 vssd1 vccd1 vccd1
+ _11873_/B sky130_fd_sc_hd__o311a_1
X_10823_ _10823_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _10823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ _10890_/B _10754_/B vssd1 vssd1 vccd1 vccd1 _10756_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10685_ _11230_/A _10684_/B _09061_/X vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__a21o_1
X_12424_ _12424_/A _12424_/B _12424_/C vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10379__A1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _12361_/B _12355_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XANTENNA__07244__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__B2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07296__A _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _11396_/B _11306_/B vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12286_ _12257_/Y _12258_/X _12112_/A vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11237_ _06831_/A _11125_/X _11143_/S vssd1 vssd1 vccd1 vccd1 _11237_/Y sky130_fd_sc_hd__o21ai_1
X_11168_ _11168_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11169_/C sky130_fd_sc_hd__xnor2_1
X_10119_ _10003_/A _10003_/B _09999_/Y vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__a21o_1
X_11099_ _10952_/A _10952_/B _10951_/A vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10450__A _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _07330_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07332_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07261_ _07261_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _07262_/B sky130_fd_sc_hd__xnor2_2
X_09000_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _11426_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_116_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07192_ _09862_/B _07192_/B vssd1 vssd1 vccd1 vccd1 _07198_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12840__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _09902_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_67_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _11726_/A _09833_/B vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08735__B2 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _06984_/A _06984_/B _10398_/A vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10360__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12986__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ _08274_/A _08715_/A2 _08735_/B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 _08716_/B
+ sky130_fd_sc_hd__o22a_1
X_09695_ _09836_/A _09695_/B vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__or2_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__A _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08646_ _08652_/A _08652_/B _08641_/A vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__07171__B1 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__A2 _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__xnor2_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07528_ _06828_/A _12718_/A _08765_/A _12716_/A vssd1 vssd1 vccd1 vccd1 _07529_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07459_ _07457_/Y _07524_/B _07454_/Y vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ _09808_/B _10588_/B hold255/A vssd1 vssd1 vccd1 vccd1 _10470_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _10203_/S _09129_/B vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__A2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__C1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _12094_/A _12096_/S _12097_/B _12097_/A vssd1 vssd1 vccd1 vccd1 _12155_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08005__A _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12071_ _06552_/A _09148_/X _12280_/A _07064_/A vssd1 vssd1 vccd1 vccd1 _12071_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07844__A _09862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__or2_1
XANTENNA__11366__A _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ hold243/X _12972_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11924_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07701__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _11620_/B _11927_/B hold220/A vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__a21oi_1
X_11786_ _11786_/A _11786_/B _11786_/C _11778_/X vssd1 vssd1 vccd1 vccd1 _11786_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10806_ _06831_/D _10803_/X _10804_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _10807_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10737_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10738_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12565_/B _12407_/B vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__or2_1
X_10668_ _10547_/A _10547_/B _10546_/A vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__B1 _10220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _11153_/A _10832_/C _10599_/C vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__or3_1
X_12338_ _12347_/A _12338_/B vssd1 vssd1 vccd1 vccd1 _12340_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12269_ reg1_val[30] _12269_/B vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08717__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B1 _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ _10692_/A _10570_/A _06830_/C _06830_/D vssd1 vssd1 vccd1 vccd1 _06835_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06761_ _06761_/A _06761_/B vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06743__A3 _12517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ _09479_/X _09478_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__mux2_1
X_06692_ reg1_val[11] _07304_/A vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__or2_1
X_08500_ _08500_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08431_ _10853_/A _08431_/B vssd1 vssd1 vccd1 vccd1 _08497_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07313_ _07875_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07315_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08293_ _08291_/A _08291_/B _08292_/Y vssd1 vssd1 vccd1 vccd1 _08304_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07244_ fanout80/X fanout78/X _08430_/B _10099_/A1 vssd1 vssd1 vccd1 vccd1 _07245_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ _07173_/Y _07375_/B _07170_/Y vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06967__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout301 _06828_/A vssd1 vssd1 vccd1 vccd1 _08274_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10515__B2 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__A1 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__B1 _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09330_/A _09796_/B _09815_/X _09120_/S _09813_/X vssd1 vssd1 vccd1 vccd1
+ _09816_/X sky130_fd_sc_hd__o221a_1
X_06959_ _07278_/A _07304_/A _07303_/B _07303_/A vssd1 vssd1 vccd1 vccd1 _06960_/B
+ sky130_fd_sc_hd__o31a_1
X_09747_ _09748_/A _09748_/B vssd1 vssd1 vccd1 vccd1 _09747_/Y sky130_fd_sc_hd__nor2_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _07153_/X _12690_/A _07277_/X _07799_/B vssd1 vssd1 vccd1 vccd1 _09679_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08782_/A2 _08735_/A2 _08735_/B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 _08630_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11640_ _11885_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11644_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _11649_/C _11571_/B vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ _10522_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10523_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13241_ _13241_/CLK _13241_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
X_10453_ _06710_/Y _10329_/X _06712_/B vssd1 vssd1 vccd1 vccd1 _10453_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10265__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _13185_/CLK _13172_/D vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08947__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10384_ _10384_/A _10384_/B vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__xnor2_1
X_12123_ _12121_/Y _12123_/B vssd1 vssd1 vccd1 vccd1 _12124_/B sky130_fd_sc_hd__nand2b_1
X_12054_ _12115_/A _06805_/Y _06815_/X _12053_/X vssd1 vssd1 vccd1 vccd1 _12056_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _11005_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__xnor2_1
X_12956_ _07187_/B _12962_/B2 hold139/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__o21a_1
XANTENNA__09675__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ hold228/X _13084_/B2 _13070_/A2 hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07686__A1 _06983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__B2 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11907_ _11909_/B vssd1 vssd1 vccd1 vccd1 _11907_/Y sky130_fd_sc_hd__inv_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11838_ _11838_/A _11838_/B _11838_/C vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__and3_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08635__B1 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07989__A2 _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08938__B2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__A1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A1 _06963_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10745__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07931_ _07933_/A _07933_/B vssd1 vssd1 vccd1 vccd1 _07931_/Y sky130_fd_sc_hd__nand2_1
X_07862_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11170__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ _08983_/B _06812_/Y _06799_/X instruction[6] _06545_/A vssd1 vssd1 vccd1
+ vccd1 _06813_/X sky130_fd_sc_hd__a2111o_1
X_09601_ _09437_/A _09437_/B _09435_/Y vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__a21oi_2
X_07793_ _09885_/A fanout37/X fanout34/X _09880_/B2 vssd1 vssd1 vccd1 vccd1 _07794_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__xnor2_1
X_06744_ _07099_/A reg1_val[3] vssd1 vssd1 vccd1 vccd1 _09785_/B sky130_fd_sc_hd__and2b_1
XANTENNA__06828__A _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06675_ _11043_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__nand2_2
X_09463_ _09771_/B _09463_/B vssd1 vssd1 vccd1 vccd1 _09617_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09204__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__B1_N _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _08350_/B _08376_/X _08394_/X _08405_/X vssd1 vssd1 vccd1 vccd1 _08414_/X
+ sky130_fd_sc_hd__a211o_1
X_09394_ _09394_/A _09394_/B _09394_/C vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__and3_1
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08345_ fanout83/X _08737_/A2 _08733_/B1 _08565_/B vssd1 vssd1 vccd1 vccd1 _08346_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09418__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ _08276_/A _08276_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07227_ _07227_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07262_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__A2 _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _07158_/A _07158_/B vssd1 vssd1 vccd1 vccd1 _07158_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11933__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07089_ reg1_val[20] reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07128_/B sky130_fd_sc_hd__or2_1
Xfanout120 _06992_/X vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__buf_6
Xfanout131 _06939_/X vssd1 vssd1 vccd1 vccd1 _08565_/B sky130_fd_sc_hd__buf_8
Xfanout153 _06976_/X vssd1 vssd1 vccd1 vccd1 _08670_/A2 sky130_fd_sc_hd__buf_8
XANTENNA__11697__C1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _09885_/A vssd1 vssd1 vccd1 vccd1 _08735_/A2 sky130_fd_sc_hd__buf_6
Xfanout164 _09568_/A vssd1 vssd1 vccd1 vccd1 _08737_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout175 _07015_/Y vssd1 vssd1 vccd1 vccd1 _09725_/B2 sky130_fd_sc_hd__buf_8
Xfanout197 _12665_/Y vssd1 vssd1 vccd1 vccd1 _12731_/A2 sky130_fd_sc_hd__buf_4
Xfanout186 _09065_/Y vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__buf_4
X_12810_ hold3/X hold298/A vssd1 vssd1 vccd1 vccd1 _13049_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12741_ hold299/X hold31/X vssd1 vssd1 vccd1 vccd1 _12742_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06876__C1 _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ hold76/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ hold263/A _11623_/B _11698_/B vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__and3_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09409__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12964__A2 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _11555_/B _11554_/B vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _11485_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__nand2_1
X_10505_ _10506_/A _11296_/A vssd1 vssd1 vccd1 vccd1 _10507_/B sky130_fd_sc_hd__nor2_1
X_13224_ _13253_/CLK _13224_/D vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12177__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10438_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _13251_/CLK _13155_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10723__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06920__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13086_ _13086_/A _13086_/B vssd1 vssd1 vccd1 vccd1 _13086_/Y sky130_fd_sc_hd__xnor2_1
X_12106_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__nand2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09345__B2 _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ _12104_/B _12037_/B vssd1 vssd1 vccd1 vccd1 _12040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08847__B _09001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ hold116/X _12665_/A _12955_/B1 hold155/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold156/A sky130_fd_sc_hd__o221a_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12385__A _12546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08608__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07831__A1 _12694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__B2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08061_ _08714_/A _08061_/B vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07012_ _07012_/A _07012_/B vssd1 vssd1 vccd1 vccd1 _07028_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08963_ _08961_/Y _08963_/B vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__and2b_1
X_07914_ _07913_/B _07913_/C _07913_/A vssd1 vssd1 vccd1 vccd1 _07927_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07347__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A1 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ _08893_/B _08894_/B vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ _07848_/A _07848_/B vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__nor2_1
X_07776_ _08688_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__xnor2_2
X_06727_ _06754_/B _06727_/B _12527_/B vssd1 vssd1 vccd1 vccd1 _06727_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07153__S _11726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ _11153_/A _09669_/B _09514_/Y _09512_/X vssd1 vssd1 vccd1 vccd1 dest_val[2]
+ sky130_fd_sc_hd__o31ai_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ _09444_/A _09444_/B _09447_/B vssd1 vssd1 vccd1 vccd1 _09446_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09869__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _06978_/B vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__inv_2
XFILLER_0_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06589_ reg2_val[28] _06748_/B _06539_/X _06588_/X vssd1 vssd1 vccd1 vccd1 _06592_/B
+ sky130_fd_sc_hd__a22o_4
X_09377_ _11183_/A _09377_/B vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__xnor2_1
X_08328_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08328_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08259_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08261_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__or2_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06740__B _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__B1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _09145_/Y _10187_/Y _10188_/X _10220_/X _10186_/Y vssd1 vssd1 vccd1 vccd1
+ _10221_/X sky130_fd_sc_hd__a311o_1
X_10152_ _11271_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__xnor2_1
X_10083_ _07158_/A _12238_/C1 _10081_/Y _10082_/X vssd1 vssd1 vccd1 vccd1 _10083_/X
+ sky130_fd_sc_hd__o2bb2a_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08948__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ hold49/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__B1 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _11094_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ reg1_val[31] _12655_/B vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ _11834_/A _11604_/X _11605_/Y vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__a21oi_1
X_12586_ _12584_/B _12592_/A vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07299__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11537_ _06636_/B _11536_/X _10828_/Y _09330_/A vssd1 vssd1 vccd1 vccd1 _11537_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06931__A _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11468_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13207_ _13208_/CLK _13207_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11373__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__nor2_1
X_10419_ _10419_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10421_/C sky130_fd_sc_hd__xor2_1
X_13138_ _13234_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11373__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13069_ hold269/X _13068_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10479__A3 _10478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ fanout41/X _12688_/A _12690_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _07631_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11284__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ _07123_/Y _07799_/B _07157_/X _07154_/X vssd1 vssd1 vccd1 vccd1 _07562_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06512_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06512_/Y sky130_fd_sc_hd__inv_2
X_09300_ _09296_/X _09299_/X _10201_/S vssd1 vssd1 vccd1 vccd1 _09300_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10636__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ _07832_/A _07492_/B vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _09432_/A _09231_/B _09223_/Y vssd1 vssd1 vccd1 vccd1 _09233_/B sky130_fd_sc_hd__or3b_1
XANTENNA__12928__A2 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _09630_/S _09165_/B _09161_/A vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08057__A1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__B2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__A1 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08113_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09093_ _09091_/X _09092_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09093_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ _08988_/A vssd1 vssd1 vccd1 vccd1 _08044_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07937__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09557__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09995_ _07000_/Y _10845_/A _10845_/B _07044_/Y _10122_/A vssd1 vssd1 vccd1 vccd1
+ _09996_/B sky130_fd_sc_hd__a32o_1
X_08946_ _07560_/B _07563_/B _07560_/A vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__08768__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _08877_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__nor2_2
XANTENNA__07391__B _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07828_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11419__A2 _11164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _07759_/A _07759_/B vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout31_A _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _10770_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10771_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _09698_/A fanout8/X fanout6/X _09568_/A vssd1 vssd1 vccd1 vccd1 _09430_/B
+ sky130_fd_sc_hd__o22a_1
X_12440_ _12427_/B _12432_/B _12496_/A vssd1 vssd1 vccd1 vccd1 _12455_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08048__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08008__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08599__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12537_/B _12372_/B vssd1 vssd1 vccd1 vccd1 _12382_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07847__A _07847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _11216_/A _11216_/B _11217_/X vssd1 vssd1 vccd1 vccd1 _11324_/B sky130_fd_sc_hd__o21ba_1
X_11253_ _12000_/A2 _11354_/B hold253/A vssd1 vssd1 vccd1 vccd1 _11253_/Y sky130_fd_sc_hd__a21oi_1
X_10204_ _10204_/A vssd1 vssd1 vccd1 vccd1 _10204_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08220__A1 _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11184_/A _11184_/B fanout3/X vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__or3_1
XANTENNA__12304__B1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _11883_/A _10135_/B vssd1 vssd1 vccd1 vccd1 _10139_/A sky130_fd_sc_hd__xnor2_1
X_10066_ _10064_/Y _10066_/B vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07582__A _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06727__C_N _12527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06926__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12083__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _10968_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__nor2_1
X_12707_ hold1/X _12720_/B _12706_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
XANTENNA__10094__B2 _10091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12638_ _12638_/A _12647_/A vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10899_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13032__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12574_/B _12569_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09539__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10149__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08800_ _08810_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _06991_/A _06990_/X _06991_/Y _07065_/A vssd1 vssd1 vccd1 vccd1 _06992_/X
+ sky130_fd_sc_hd__a22o_1
X_09780_ _10320_/B _09778_/X _09779_/Y vssd1 vssd1 vccd1 vccd1 _09780_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _08731_/A _08731_/B vssd1 vssd1 vccd1 vccd1 _08732_/B sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__A3 _09147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ _08662_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__xor2_1
X_07613_ fanout82/X _11387_/A _11462_/A _06940_/A vssd1 vssd1 vccd1 vccd1 _07614_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12838__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout166_A _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__xnor2_1
X_07544_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07746_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _07475_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07549_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ fanout82/X fanout76/X fanout74/X _06940_/A vssd1 vssd1 vccd1 vccd1 _09215_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09778__A1 _10321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _09146_/A _09153_/A vssd1 vssd1 vccd1 vccd1 _09145_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__07789__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ reg1_val[5] reg1_val[26] _09092_/S vssd1 vssd1 vccd1 vccd1 _09076_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08031_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ fanout74/X fanout42/X _07239_/A fanout68/X vssd1 vssd1 vccd1 vccd1 _09979_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06531__B_N _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _09862_/B _08929_/B vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ _12179_/A _11914_/X _11915_/Y _11939_/X _11913_/Y vssd1 vssd1 vccd1 vccd1
+ _11940_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_98_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _11871_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11871_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12065__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10822_ hold259/A _09808_/B _10930_/B _10821_/Y _09810_/A vssd1 vssd1 vccd1 vccd1
+ _10826_/B sky130_fd_sc_hd__a311o_1
XANTENNA__09466__B1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__A _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _10890_/A _10751_/Y _10606_/Y _10612_/A vssd1 vssd1 vccd1 vccd1 _10754_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10684_ _11230_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10684_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09218__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _12424_/A _12424_/B _12424_/C vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12222__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__A2 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12354_/A _12354_/B _12354_/C vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07244__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _11304_/A _11304_/B _11304_/C vssd1 vssd1 vccd1 vccd1 _11306_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12285_ _07255_/A _06905_/Y _12261_/X _12284_/X _12080_/A vssd1 vssd1 vccd1 vccd1
+ dest_val[30] sky130_fd_sc_hd__o221a_4
X_11236_ _11236_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11236_/Y sky130_fd_sc_hd__xnor2_1
X_11167_ _11296_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10731__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11098_ _11000_/A _11000_/B _10998_/Y vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10049_ _10049_/A _10310_/A vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07261_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07191_ _12714_/A _09727_/A _08798_/B _12716_/A vssd1 vssd1 vccd1 vccd1 _07192_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12393__A _12553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09901_ _09902_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ _10876_/A1 fanout47/X _07277_/X _07154_/X vssd1 vssd1 vccd1 vccd1 _09833_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08735__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09764_/B _09764_/A vssd1 vssd1 vccd1 vccd1 _09763_/Y sky130_fd_sc_hd__nand2b_1
X_06975_ _08698_/A _06975_/B vssd1 vssd1 vccd1 vccd1 _06984_/B sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__xnor2_1
X_09694_ _09694_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__and2_1
XANTENNA__07171__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _08644_/Y _08607_/A _08683_/A vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07171__B2 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__nor2_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _09423_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11255__B1 _09138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ _07458_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07524_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07389_ _07389_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07449_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ _09111_/X _09127_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _12267_/A _12223_/B _12223_/C _12299_/A vssd1 vssd1 vccd1 vccd1 _10320_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_0_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _06552_/A _09141_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__a21o_1
X_11021_ _10449_/A _09031_/A _09031_/B _12179_/A vssd1 vssd1 vccd1 vccd1 _11022_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10533__A2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ _12972_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12972_/Y sky130_fd_sc_hd__xnor2_1
X_11923_ _11921_/Y _11923_/B vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__and2b_1
X_11854_ hold191/A _11854_/B vssd1 vssd1 vccd1 vccd1 _11927_/B sky130_fd_sc_hd__or2_1
X_10805_ _10803_/X _10804_/Y _06831_/D vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11785_ _09152_/Y _11780_/X _11781_/Y _11784_/X vssd1 vssd1 vccd1 vccd1 _11786_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08111__B1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10883_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _10667_/A _10667_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__xnor2_2
X_12406_ _12565_/B _12407_/B vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06947__A1_N _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10598_ curr_PC[9] _10597_/C curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10599_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10221__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ _12512_/B _12337_/B vssd1 vssd1 vccd1 vccd1 _12338_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12268_ reg1_val[30] _12269_/B vssd1 vssd1 vccd1 vccd1 _12302_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08178__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11327_/A sky130_fd_sc_hd__and2_1
X_12199_ _12245_/B _12199_/B vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06760_ _06753_/B _06537_/Y _12507_/B _06754_/X reg1_val[1] vssd1 vssd1 vccd1 vccd1
+ _06761_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09678__B1 _07277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ reg1_val[11] _07304_/A vssd1 vssd1 vccd1 vccd1 _10706_/S sky130_fd_sc_hd__nand2_1
XANTENNA__07770__A _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08430_ _08755_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08431_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06900__A1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__A1 _07028_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _08359_/A _08359_/B _08360_/Y vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ _11564_/A _12686_/A fanout38/X _12688_/A vssd1 vssd1 vccd1 vccd1 _07313_/B
+ sky130_fd_sc_hd__o22a_1
X_08292_ _08352_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08292_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ _07243_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07010__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _07174_/A _07174_/B vssd1 vssd1 vccd1 vccd1 _07375_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12062__S _12271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12570__B _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _06511_/Y vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09815_ _11135_/S _09814_/Y _09168_/A vssd1 vssd1 vccd1 vccd1 _09815_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10515__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__A1 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06958_ _07304_/A _07303_/B _07303_/A vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__o21a_2
X_09746_ _09574_/A _09574_/B _09572_/Y vssd1 vssd1 vccd1 vccd1 _09748_/B sky130_fd_sc_hd__a21oi_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ _09680_/A vssd1 vssd1 vccd1 vccd1 _09677_/Y sky130_fd_sc_hd__inv_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__A1 _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ instruction[6] instruction[5] _09148_/A vssd1 vssd1 vccd1 vccd1 _06889_/Y
+ sky130_fd_sc_hd__nor3_4
XANTENNA__08341__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ _08647_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _08628_/Y sky130_fd_sc_hd__nor2_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08559_ _08841_/C _08559_/B vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__and2_1
X_11570_ _11649_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout8_A fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ _10522_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__and2_1
X_13240_ _13241_/CLK _13240_/D vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10452_ _11232_/A _09022_/A _09022_/B _09145_/Y _10451_/Y vssd1 vssd1 vccd1 vccd1
+ _10452_/X sky130_fd_sc_hd__o311a_1
X_13171_ _13185_/CLK hold209/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06958__A1 _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A2 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ _10384_/A _10384_/B vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12122_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__nand2_1
X_12053_ _12053_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__and2_1
XANTENNA__07907__B1 _08741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__xnor2_1
X_12955_ hold138/X _12662_/A _12955_/B1 _13219_/Q _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold139/A sky130_fd_sc_hd__o221a_1
XANTENNA__07590__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _11976_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11909_/B sky130_fd_sc_hd__and2_1
X_12886_ _13071_/A hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07686__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11837_ _12110_/B _11836_/B _09061_/X vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__a21o_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11767_/A _11767_/B _11767_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _11786_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08635__A1 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09832__B1 _07277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08635__B2 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _11153_/A _10719_/B _10719_/C vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__or3_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _11623_/B _11776_/B hold269/A vssd1 vssd1 vccd1 vccd1 _11699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08399__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__A2 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07610__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07930_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07933_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07861_ _07861_/A _07861_/B vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__and2_1
X_06812_ _12264_/A _06811_/X _06823_/A vssd1 vssd1 vccd1 vccd1 _06812_/Y sky130_fd_sc_hd__o21ai_1
X_07792_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07857_/A sky130_fd_sc_hd__xnor2_1
X_09600_ _09600_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11170__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06743_ _06763_/B _06646_/A _12517_/B _06742_/X vssd1 vssd1 vccd1 vccd1 _07099_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ _09532_/B _09532_/A vssd1 vssd1 vccd1 vccd1 _09531_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__06828__B _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06674_ reg1_val[14] _06963_/A vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _08982_/A _09774_/A _09460_/Y vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__a21o_2
XANTENNA__12846__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08413_ _08474_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__nor2_1
X_09393_ _09394_/A _09394_/B _09394_/C vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout246_A _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08344_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08410_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12565__B _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08276_/B _08276_/C _08276_/A vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10366__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ _07227_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07569_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_15_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13185_/CLK sky130_fd_sc_hd__clkbuf_8
X_07157_ _07158_/A _07158_/B vssd1 vssd1 vccd1 vccd1 _07157_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07088_ reg1_val[19] _07088_/B vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__or2_1
Xfanout121 _10957_/A vssd1 vssd1 vccd1 vccd1 _10490_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout110 _11956_/A vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout165 _07098_/Y vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__buf_8
Xfanout143 _07146_/X vssd1 vssd1 vccd1 vccd1 _09885_/A sky130_fd_sc_hd__buf_8
Xfanout154 _10156_/A vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__buf_8
Xfanout132 _12686_/A vssd1 vssd1 vccd1 vccd1 _09180_/B2 sky130_fd_sc_hd__buf_8
Xfanout198 _12730_/B vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__buf_4
XANTENNA__11925__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _09064_/Y vssd1 vssd1 vccd1 vccd1 _09092_/S sky130_fd_sc_hd__clkbuf_8
Xfanout176 _07011_/X vssd1 vssd1 vccd1 vccd1 _08740_/A2 sky130_fd_sc_hd__buf_6
X_09729_ _09730_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09855_/C sky130_fd_sc_hd__nor2_1
XANTENNA__06738__B _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11136__S _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ hold31/X hold281/X vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _07185_/Y _12962_/B2 hold54/X _12970_/A vssd1 vssd1 vccd1 vccd1 _13128_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11653__A_N _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ hold283/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11698_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11553_ _11799_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11484_ _11485_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__or2_1
X_10504_ _10504_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__xnor2_1
X_13223_ _13253_/CLK _13223_/D vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10435_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10435_/Y sky130_fd_sc_hd__nand2b_1
X_13154_ _13251_/CLK _13154_/D vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_12105_ _12104_/A _12104_/B _12104_/C vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__a21o_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ _11656_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__xnor2_1
X_13085_ _13085_/A hold282/X vssd1 vssd1 vccd1 vccd1 _13248_/D sky130_fd_sc_hd__and2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10297_/A _10297_/B vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__xor2_1
X_12036_ _12036_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ _11068_/A _12962_/B2 hold117/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__o21a_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ hold184/X _13070_/B2 _13070_/A2 hold179/X vssd1 vssd1 vccd1 vccd1 hold185/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11570__A _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A1 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08608__B2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07292__B1 _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__A2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _08670_/A2 _10506_/A _10647_/A _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08061_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07011_ _07015_/B _07015_/A _08698_/A vssd1 vssd1 vccd1 vccd1 _07011_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10914__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ _08962_/A _08962_/B vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07913_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__nand3_2
X_08893_ _08894_/B _08893_/B vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__and2b_1
XANTENNA_fanout196_A _12731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__B2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07844_ _09862_/B _07844_/B vssd1 vssd1 vccd1 vccd1 _07848_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07775_ _12706_/A _09727_/A _08798_/B fanout77/X vssd1 vssd1 vccd1 vccd1 _07776_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09215__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06726_ _06512_/Y _06532_/X _06535_/Y _12527_/B _06753_/B vssd1 vssd1 vccd1 vccd1
+ _06726_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09514_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09514_/Y sky130_fd_sc_hd__a21oi_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06657_ reg2_val[16] _06700_/B _06657_/B1 _06656_/Y vssd1 vssd1 vccd1 vccd1 _06978_/B
+ sky130_fd_sc_hd__a22o_2
X_09445_ _09264_/A _09264_/B _09262_/Y vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__a21oi_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06588_ _06613_/A _12565_/B vssd1 vssd1 vccd1 vccd1 _06588_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09376_ fanout80/X fanout36/X fanout34/X _10099_/A1 vssd1 vssd1 vccd1 vccd1 _09377_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08327_ _08688_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08258_ _08259_/B _08259_/A vssd1 vssd1 vccd1 vccd1 _08857_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09885__A _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07209_ fanout80/X _08430_/B _10490_/B2 fanout79/X vssd1 vssd1 vccd1 vccd1 _07210_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _10220_/A _10220_/B _10219_/X vssd1 vssd1 vccd1 vccd1 _10220_/X sky130_fd_sc_hd__or3b_2
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08189_ _08189_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07586__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__B2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _11739_/A fanout42/X _07239_/A fanout64/X vssd1 vssd1 vccd1 vccd1 _10152_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ hold289/A _09808_/B _10210_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _10082_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _10983_/B _10983_/C _10983_/A vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__o21a_1
X_12723_ _07044_/Y _12731_/A2 hold96/X _13103_/A vssd1 vssd1 vccd1 vccd1 _13154_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10645__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12654_ _12651_/A _12653_/B _12651_/B vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _11834_/A _11604_/X _10450_/A vssd1 vssd1 vccd1 vccd1 _11605_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07299__B _07301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12585_ _12585_/A _12585_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xnor2_4
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ _11535_/A _09141_/Y _11535_/Y _12309_/B1 vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13206_ _13208_/CLK hold87/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06931__B _06931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ _11656_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11398_ _11177_/A _11177_/B _11280_/B _11279_/A vssd1 vssd1 vccd1 vccd1 _11401_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ _11271_/A _10418_/B vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__xnor2_1
X_13137_ _13234_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_10349_ _06712_/B _11625_/B _10344_/Y _06710_/Y _10348_/X vssd1 vssd1 vccd1 vccd1
+ _10349_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11373__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__B1_N _11883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13068_/Y sky130_fd_sc_hd__xnor2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _12020_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12097_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08858__B _08858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06659__A _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ _07560_/A _07560_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06511_ _12499_/A vssd1 vssd1 vccd1 vccd1 _06511_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10636__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07491_ fanout80/X _08606_/A2 _08642_/B _10099_/A1 vssd1 vssd1 vccd1 vccd1 _07492_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _09432_/A _09231_/B _09223_/Y vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__nor3b_1
XANTENNA__10636__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _09161_/A vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08057__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ reg1_val[8] reg1_val[23] _09092_/S vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__mux2_1
X_08112_ _08734_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08988_/A sky130_fd_sc_hd__or2_2
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout209_A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout111_A _11887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09557__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _09994_/A _09994_/B vssd1 vssd1 vccd1 vccd1 _10028_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12313__A1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__B _08768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__xnor2_1
X_08876_ _08877_/B _08876_/B vssd1 vssd1 vccd1 vccd1 _08876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07827_ _07827_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07892_/B sky130_fd_sc_hd__xnor2_2
X_07758_ _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07759_/B sky130_fd_sc_hd__and2_1
X_06709_ _07137_/A reg1_val[8] vssd1 vssd1 vccd1 vccd1 _06775_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08784__A _08784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _07689_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ _09428_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__A2 _08733_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ fanout13/X _10370_/A _07763_/B fanout47/X vssd1 vssd1 vccd1 vccd1 _09360_/B
+ sky130_fd_sc_hd__o22ai_1
X_12370_ reg1_val[8] curr_PC[8] _12495_/S vssd1 vssd1 vccd1 vccd1 _12372_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07256__B1 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11324_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06751__B _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ hold267/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _10200_/X _10202_/X _10203_/S vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08756__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08220__A2 _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _07183_/A _07183_/B _07763_/B _10647_/A fanout45/X vssd1 vssd1 vccd1 vccd1
+ _10135_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10065_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06534__A2 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06926__B _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A2 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10729__A _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ _10967_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12706_ _12706_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12706_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _10898_/A _10898_/B vssd1 vssd1 vccd1 vccd1 _10899_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12637_ reg1_val[28] _12656_/A vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__and2_1
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13032__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12663__B _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__A _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ _12568_/A _12568_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12569_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_11519_ _12053_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__and2_1
XANTENNA__06661__B _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ _12499_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _06991_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__nor2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08730_ _08730_/A _08730_/B _08730_/C vssd1 vssd1 vccd1 vccd1 _08731_/B sky130_fd_sc_hd__or3_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _08814_/A _08661_/B vssd1 vssd1 vccd1 vccd1 _08662_/B sky130_fd_sc_hd__xnor2_1
X_07612_ _07616_/A vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__inv_2
XFILLER_0_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08592_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__nor2_1
X_07543_ _07543_/A _07543_/B vssd1 vssd1 vccd1 vccd1 _07745_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10085__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _07475_/B _07475_/A vssd1 vssd1 vccd1 vccd1 _07474_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _09979_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12854__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _12309_/B1 _09143_/X _06829_/B vssd1 vssd1 vccd1 vccd1 _09155_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12231__B1 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07789__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09075_ _09073_/X _09074_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06571__B _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__clkbuf_8
X_08026_ _08026_/A _08026_/B _08026_/C vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__or3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07683__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09977_ _09831_/B _09834_/B _09831_/A vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__12837__A2 hold177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12298__B1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _07057_/Y _10845_/A _10845_/B _09224_/A _07044_/Y vssd1 vssd1 vccd1 vccd1
+ _08929_/B sky130_fd_sc_hd__a32o_1
X_08859_ _08865_/B _08859_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11870_ _11600_/A _11600_/B _11600_/C _11681_/A _11869_/Y vssd1 vssd1 vccd1 vccd1
+ _11873_/A sky130_fd_sc_hd__a2111o_1
X_10821_ _12304_/B1 _10930_/B hold259/A vssd1 vssd1 vccd1 vccd1 _10821_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09466__A1 _09617_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06746__B _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752_ _10606_/Y _10612_/A _10890_/A _10751_/Y vssd1 vssd1 vccd1 vccd1 _10890_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12422_ _12429_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _12424_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11025__A1 _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__B2 _10852_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ _11232_/A _10683_/B vssd1 vssd1 vccd1 vccd1 _10684_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12353_ _12354_/A _12354_/B _12354_/C vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10284__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ _09145_/Y _12267_/Y _12283_/Y _12265_/X vssd1 vssd1 vccd1 vccd1 _12284_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _11304_/A _11304_/B _11304_/C vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__or3_1
X_11235_ _11235_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11295_/B2 fanout7/X fanout5/X _11297_/A vssd1 vssd1 vccd1 vccd1 _11167_/B
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13230_/CLK sky130_fd_sc_hd__clkbuf_8
X_10117_ _10117_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__nor2_1
X_11097_ _10993_/A _10993_/B _10992_/A vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__o21a_1
X_10048_ _10048_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06937__A _06938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _12000_/A2 _12063_/B hold299/A vssd1 vssd1 vccd1 vccd1 _11999_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11264__A1 _11713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10472__C1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07190_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ _09749_/A _09749_/B _09747_/Y vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _09831_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__nor2_1
X_06974_ _08698_/A _06975_/B vssd1 vssd1 vccd1 vccd1 _06984_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07943__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__xnor2_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _10398_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08713_/Y sky130_fd_sc_hd__nand2_1
X_09693_ _09694_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06847__A _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08644_ _08683_/B vssd1 vssd1 vccd1 vccd1 _08644_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07171__A2 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09223__A _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08575_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__and2_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _12712_/A _09422_/A _09222_/B2 _12714_/A vssd1 vssd1 vccd1 vccd1 _07527_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _07524_/A vssd1 vssd1 vccd1 vccd1 _07457_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _09423_/A _07388_/B vssd1 vssd1 vccd1 vccd1 _07449_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ _09126_/X _09119_/X _10073_/S vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _08009_/A vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ _10449_/A _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11191__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12971_ _12787_/X _12971_/B vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__nand2b_1
X_11922_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11663__A _11663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ hold292/A _11623_/B _11851_/X _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11853_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10804_ _06690_/Y _06779_/X _11124_/A vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10279__A _11654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11784_ _09064_/Y _10463_/X _10476_/Y _09135_/Y _11783_/Y vssd1 vssd1 vccd1 vccd1
+ _11784_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08111__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08111__B2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _11068_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10666_ _10666_/A _10666_/B vssd1 vssd1 vccd1 vccd1 _10667_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10206__C1 _09156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _10920_/A curr_PC[13] _12444_/S vssd1 vssd1 vccd1 vccd1 _12407_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ curr_PC[9] curr_PC[10] _10597_/C vssd1 vssd1 vccd1 vccd1 _10832_/C sky130_fd_sc_hd__and3_1
X_12336_ _12512_/B _12337_/B vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12267_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08178__A1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__A _11656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12198_ fanout9/A fanout5/X fanout4/X fanout7/X vssd1 vssd1 vccd1 vccd1 _12199_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08178__B2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__xnor2_1
X_11149_ _06889_/Y _11136_/X _11148_/X _11128_/X vssd1 vssd1 vccd1 vccd1 _11149_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11182__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09678__B2 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _07304_/A reg1_val[11] vssd1 vssd1 vccd1 vccd1 _06690_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10693__C1 _09498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08360_ _08372_/B _08372_/A vssd1 vssd1 vccd1 vccd1 _08360_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07311_ _11468_/A _07311_/B vssd1 vssd1 vccd1 vccd1 _07315_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11788__A2 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07242_ _07243_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07572_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07173_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__B1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout303 reg1_val[13] vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__buf_8
X_09814_ _11134_/S _09635_/Y _09166_/B vssd1 vssd1 vccd1 vccd1 _09814_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07392__A2 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06957_ _10982_/A _06957_/B vssd1 vssd1 vccd1 vccd1 _06957_/X sky130_fd_sc_hd__and2_1
X_09745_ _09877_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__nand2_1
X_06888_ instruction[22] _06850_/Y _06887_/X _06637_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__o211a_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09676_ _11883_/A _09676_/B vssd1 vssd1 vccd1 vccd1 _09680_/A sky130_fd_sc_hd__xnor2_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__B2 _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ _08627_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _08647_/B sky130_fd_sc_hd__or2_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11228__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07509_ _07730_/A _07730_/B _07505_/X vssd1 vssd1 vccd1 vccd1 _07536_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ _08734_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09099__S _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10451_ _11232_/A _09022_/B _09022_/A vssd1 vssd1 vccd1 vccd1 _10451_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10739__B1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _13185_/CLK hold188/X vssd1 vssd1 vccd1 vccd1 _13170_/Q sky130_fd_sc_hd__dfxtp_1
X_10382_ _12086_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _12005_/A _11986_/B _06566_/A vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__09357__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11003_/A _11003_/B _11004_/A vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__and3_1
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12954_ _12085_/A _12962_/B2 hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__o21a_1
XFILLER_0_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11905_ _11905_/A _11905_/B _11905_/C vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__or3_1
X_12885_ hold231/A _12885_/A2 _12885_/B1 hold228/X vssd1 vssd1 vccd1 vccd1 hold229/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _12110_/B _11836_/B vssd1 vssd1 vccd1 vccd1 _11836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08635__A2 _08737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07843__B1 _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__B _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__B2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ curr_PC[11] _10832_/C vssd1 vssd1 vccd1 vccd1 _10719_/C sky130_fd_sc_hd__and2_1
X_11698_ hold263/A _11698_/B vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08399__A1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ _12089_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__B2 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _12499_/B _12319_/B vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__or2_1
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ _07961_/A _07961_/B _07856_/Y vssd1 vssd1 vccd1 vccd1 _07879_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12399__A _12559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ _12221_/A _06810_/X _06821_/A vssd1 vssd1 vccd1 vccd1 _06811_/X sky130_fd_sc_hd__o21a_1
X_07791_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__and2_1
X_06742_ reg2_val[3] _06748_/B vssd1 vssd1 vccd1 vccd1 _06742_/X sky130_fd_sc_hd__and2_1
X_09530_ _09530_/A _09530_/B vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__xnor2_1
X_09461_ _09461_/A _09461_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__and2_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08874__A2 _08871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ reg1_val[14] _06963_/A vssd1 vssd1 vccd1 vccd1 _11043_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08412_ _08412_/A _08412_/B vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ _09211_/A _09208_/X _09210_/A vssd1 vssd1 vccd1 vccd1 _09394_/C sky130_fd_sc_hd__o21a_1
XANTENNA__12958__A1 _12142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08343_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08343_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13023__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout239_A _07108_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08274_ _08274_/A _11169_/A vssd1 vssd1 vccd1 vccd1 _08276_/C sky130_fd_sc_hd__nor2_1
XANTENNA__10647__A _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B1 _08135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ _07225_/A _07225_/B vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08117__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__A2 _12304_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _07156_/A _07156_/B vssd1 vssd1 vccd1 vccd1 _07156_/X sky130_fd_sc_hd__or2_4
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ reg1_val[18] _07087_/B vssd1 vssd1 vccd1 vccd1 _07088_/B sky130_fd_sc_hd__or2_1
XANTENNA__11478__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A _12086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout122 _06963_/Y vssd1 vssd1 vccd1 vccd1 _10957_/A sky130_fd_sc_hd__buf_8
Xfanout111 _11887_/A vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__buf_8
Xfanout100 _12702_/A vssd1 vssd1 vccd1 vccd1 _10359_/B2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11697__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout144 _08689_/B1 vssd1 vssd1 vccd1 vccd1 _12684_/A sky130_fd_sc_hd__buf_8
Xfanout155 _10853_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__buf_12
Xfanout133 _12686_/A vssd1 vssd1 vccd1 vccd1 _10370_/A sky130_fd_sc_hd__clkbuf_4
Xfanout177 _07011_/X vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__buf_6
Xfanout199 _12664_/Y vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__buf_4
XANTENNA__07691__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout188 _08698_/A vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__clkbuf_16
Xfanout166 _08798_/B vssd1 vssd1 vccd1 vccd1 _08756_/B2 sky130_fd_sc_hd__buf_6
X_07989_ _08274_/A _11663_/A _08813_/A1 fanout76/X vssd1 vssd1 vccd1 vccd1 _07990_/B
+ sky130_fd_sc_hd__o22a_2
X_09728_ _09862_/B _09728_/B vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout54_A _12718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _11238_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _09659_/Y sky130_fd_sc_hd__nand2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ hold53/X _12692_/B vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11781_/B _11701_/B hold210/A vssd1 vssd1 vccd1 vccd1 _11621_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _07044_/Y _07154_/X _07799_/B _07069_/X vssd1 vssd1 vccd1 vccd1 _11553_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11483_ _11483_/A _11483_/B vssd1 vssd1 vccd1 vccd1 _11485_/B sky130_fd_sc_hd__xnor2_1
X_10503_ _11296_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__xnor2_1
X_13222_ _13222_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07866__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10434_ _10434_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__xor2_1
X_13153_ _13250_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10365_ _11295_/B2 fanout50/X _07988_/B _11462_/A vssd1 vssd1 vccd1 vccd1 _10366_/B
+ sky130_fd_sc_hd__o22a_1
X_12104_ _12104_/A _12104_/B _12104_/C vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__nand3_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13084_ hold281/X _13084_/A2 _13083_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 hold282/A
+ sky130_fd_sc_hd__a22o_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10297_/A _10297_/B vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ _12036_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12104_/B sky130_fd_sc_hd__or2_1
XANTENNA__08002__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A _13111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ _13209_/Q _12665_/A _12955_/B1 hold116/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold117/A sky130_fd_sc_hd__o221a_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10112__A1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__B2 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ _13062_/A hold219/X vssd1 vssd1 vccd1 vccd1 _13175_/D sky130_fd_sc_hd__and2_1
XANTENNA__11860__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12666__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _11819_/A _11819_/B _11819_/C vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__nor3_1
XANTENNA__11570__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12799_ _12994_/B _12995_/A _12775_/X vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__a21o_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08608__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07292__A1 _12684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__B2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07010_ _08688_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07015_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06680__A _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07776__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08961_ _08962_/A _08962_/B vssd1 vssd1 vccd1 vccd1 _08961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07912_ _07909_/B _07909_/C _07909_/A vssd1 vssd1 vccd1 vccd1 _07913_/C sky130_fd_sc_hd__a21o_1
X_08892_ _12085_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08893_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07347__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _12704_/A _09727_/A _08798_/B _12706_/A vssd1 vssd1 vccd1 vccd1 _07844_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09741__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08400__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _10252_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__xnor2_2
X_06725_ _06723_/Y _06725_/B vssd1 vssd1 vccd1 vccd1 _06832_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__and3_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06656_ _06727_/B _12501_/B vssd1 vssd1 vccd1 vccd1 _06656_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__nand2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12576__B _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06587_ instruction[38] _06637_/B vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__and2_4
XFILLER_0_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06574__B _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09375_ _11796_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__xnor2_1
X_08326_ _08756_/B2 fanout93/X _12690_/A _09727_/A vssd1 vssd1 vccd1 vccd1 _08327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ _08257_/A _08257_/B vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09885__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06590__A _06592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ _08916_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07354_/A sky130_fd_sc_hd__xnor2_2
X_08188_ _08188_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07139_ _10117_/A fanout51/X _12684_/A fanout49/X vssd1 vssd1 vccd1 vccd1 _07140_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11367__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _10529_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _09808_/B _10210_/B hold289/A vssd1 vssd1 vccd1 vccd1 _10081_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12316__C1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10983_ _10983_/A _10983_/B _10983_/C vssd1 vssd1 vccd1 vccd1 _11094_/A sky130_fd_sc_hd__nor3_2
X_12722_ hold95/X _12730_/B vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12653_ _12653_/A _12653_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ _12110_/A _11834_/B _11232_/A vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__a21o_1
X_12584_ _12584_/A _12584_/B _12585_/B vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__or3_1
XFILLER_0_25_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11535_ _11535_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13205_ _13217_/CLK hold143/X vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__dfxtp_1
X_11466_ _12148_/A fanout50/X _07988_/B _12201_/A vssd1 vssd1 vccd1 vccd1 _11467_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11397_ _11303_/A _11303_/B _11302_/A vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__o21ai_1
X_10417_ _11876_/A fanout42/X _07239_/A _11950_/A vssd1 vssd1 vccd1 vccd1 _10418_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13136_ _13260_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_10348_ _07137_/A _12238_/C1 _10346_/Y _10347_/X vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13071_/A hold270/X vssd1 vssd1 vccd1 vccd1 _13244_/D sky130_fd_sc_hd__and2_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _11654_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__xnor2_1
X_12018_ _07106_/A fanout4/X _12017_/Y vssd1 vssd1 vccd1 vccd1 _12020_/B sky130_fd_sc_hd__o21a_1
XANTENNA__06659__B _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07490_ _07501_/A _07490_/B vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06510_ instruction[3] vssd1 vssd1 vccd1 vccd1 _06892_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10636__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _09113_/Y _09165_/B _09309_/S vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__mux2_1
X_09091_ reg1_val[9] reg1_val[22] _09092_/S vssd1 vssd1 vccd1 vccd1 _09091_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08111_ _11295_/B2 _08815_/B _11297_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08112_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _08042_/A _08042_/B _08042_/C vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12010__B2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _09991_/X _09993_/B vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07953__B _07953_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__C _08768_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _07897_/Y _08986_/B _08876_/B vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__10324__A1 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ _07826_/A _07826_/B vssd1 vssd1 vccd1 vccd1 _07892_/A sky130_fd_sc_hd__nor2_2
X_07757_ _07756_/B _07756_/C _07756_/A vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06708_ _06763_/B _06646_/A _12542_/B _06707_/X vssd1 vssd1 vccd1 vccd1 _07137_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ _10099_/A1 _08670_/A2 _06984_/Y _12702_/A vssd1 vssd1 vccd1 vccd1 _07689_/B
+ sky130_fd_sc_hd__o22a_1
X_06639_ reg2_val[18] _06700_/B _06657_/B1 _06638_/X vssd1 vssd1 vccd1 vccd1 _06991_/A
+ sky130_fd_sc_hd__a22oi_2
X_09427_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09358_ _11883_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _09362_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07256__B2 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__A1 _08765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08309_ _08309_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _09115_/X _09158_/B _09630_/S vssd1 vssd1 vccd1 vccd1 _09289_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11320_ _11412_/B _11320_/B vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__or2_1
XANTENNA__10260__B1 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11251_ hold184/A _11781_/B _11348_/B _11448_/A vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__a31o_1
X_10202_ _10201_/X _09166_/A _11134_/S vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08756__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ _12201_/A fanout36/X fanout34/X fanout9/X vssd1 vssd1 vccd1 vccd1 _11183_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11760__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _10275_/A _10132_/C _10132_/A vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10563__A1 _10681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10064_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11385__B _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ _10967_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__and2_1
X_12705_ hold3/X _12720_/B _12704_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
XANTENNA__13105__B fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10897_ _10898_/B _10898_/A vssd1 vssd1 vccd1 vccd1 _10897_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07103__B _07103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12636_ reg1_val[28] _12656_/A vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06942__B _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _12568_/A _12568_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11518_ _11431_/A _11429_/X _11439_/S vssd1 vssd1 vccd1 vccd1 _11519_/B sky130_fd_sc_hd__a21bo_1
X_12498_ reg1_val[0] instruction[25] _12498_/C vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__and3_4
XANTENNA__08215__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _11443_/Y _11444_/X _11448_/X vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13119_ hold133/X _12663_/B _12660_/Y _12664_/A vssd1 vssd1 vccd1 vccd1 _13121_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _06979_/A _06979_/B _06979_/C _07289_/B vssd1 vssd1 vccd1 vccd1 _06990_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08813_/A1 _08689_/B1 _09180_/B2 _08274_/A vssd1 vssd1 vccd1 vccd1 _08661_/B
+ sky130_fd_sc_hd__o22a_1
X_07611_ _11271_/A _07611_/B vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08591_ _08591_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__nand2_1
X_07542_ _07542_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _07745_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07473_ _07473_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _10099_/A1 fanout42/X _07239_/A _10359_/B2 vssd1 vssd1 vccd1 vccd1 _09213_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10490__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _12265_/C1 _09141_/Y _08823_/B vssd1 vssd1 vccd1 vccd1 _09143_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout221_A _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07789__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__B1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ reg1_val[6] reg1_val[25] _09092_/S vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08125__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout2 hold246/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__clkbuf_8
X_08025_ _08034_/B _08034_/A vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07410__A1 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12298__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _09564_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__xnor2_2
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__xnor2_1
X_07809_ _07813_/A vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__inv_2
X_08789_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__nor2_1
X_10820_ hold261/A _10820_/B vssd1 vssd1 vccd1 vccd1 _10930_/B sky130_fd_sc_hd__or2_1
XANTENNA__11258__C1 _11257_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12110__A _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _07277_/X _12029_/B _10638_/X _10644_/A vssd1 vssd1 vccd1 vccd1 _10751_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ _12576_/B _12421_/B vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09218__A2 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ _10449_/C _11231_/B vssd1 vssd1 vccd1 vccd1 _10683_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12352_ _12361_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12354_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06988__B1 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12283_ _12303_/A _12271_/X _12282_/X vssd1 vssd1 vccd1 vccd1 _12283_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11981__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _11303_/A _11303_/B vssd1 vssd1 vccd1 vccd1 _11304_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11234_ _11233_/A _11233_/B _10450_/A vssd1 vssd1 vccd1 vccd1 _11234_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13087__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11069__A_N _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _11073_/A _11073_/B _11069_/X vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__a21oi_2
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__nor2_1
X_11096_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _10048_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__nor2_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06937__B _06938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ hold271/A _11998_/B vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07114__A _12085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ _10950_/A _10950_/B _10950_/C vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10472__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10348__A1_N _07137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12619_ _12619_/A _12624_/A vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12690__A _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09475__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__nor2_1
X_06973_ reg1_val[8] _06973_/B vssd1 vssd1 vccd1 vccd1 _06975_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07943__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ _09604_/A _09604_/B _09602_/Y vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__a21oi_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__xnor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _09550_/A _09549_/B _09549_/A vssd1 vssd1 vccd1 vccd1 _09694_/B sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout171_A _07041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _08643_/A _08643_/B vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _08605_/A _08605_/B vssd1 vssd1 vccd1 vccd1 _08579_/A sky130_fd_sc_hd__nor2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _12085_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11255__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07456_ _09423_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07524_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07387_ _09422_/A _12716_/A _12718_/A _09222_/B2 vssd1 vssd1 vccd1 vccd1 _07388_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10215__B1 _09148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ _09122_/X _09125_/X _09479_/S vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _12223_/C sky130_fd_sc_hd__xor2_4
XANTENNA__09620__A2 _10321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _08714_/A _08008_/B vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11715__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A1 _11462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__A3 _12522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _11235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _11636_/S _09955_/X _09958_/X vssd1 vssd1 vccd1 vccd1 dest_val[5] sky130_fd_sc_hd__o21ai_4
XANTENNA__11191__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _12970_/A hold244/X vssd1 vssd1 vccd1 vccd1 _13224_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11921_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06757__B _09479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__B _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _11623_/B _11851_/X hold292/A vssd1 vssd1 vccd1 vccd1 _11852_/Y sky130_fd_sc_hd__a21oi_1
X_10803_ _11124_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__and2_1
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ _09138_/X _11782_/X _06611_/B vssd1 vssd1 vccd1 vccd1 _11783_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__A2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ _11950_/A fanout37/X _08233_/B _12095_/A vssd1 vssd1 vccd1 vccd1 _10735_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _10663_/A _10663_/B _10666_/B vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12404_ _12410_/B _12404_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XFILLER_0_36_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12335_ reg1_val[3] curr_PC[3] _12444_/S vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10596_ _10566_/Y _10567_/X _10595_/X _10565_/Y vssd1 vssd1 vccd1 vccd1 _10596_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09295__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12266_ _12223_/B _12223_/C _12223_/A vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12197_ _06592_/B _06905_/Y _12196_/X _12080_/A vssd1 vssd1 vccd1 vccd1 dest_val[28]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__08178__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _11218_/B _11218_/A vssd1 vssd1 vccd1 vccd1 _11217_/X sky130_fd_sc_hd__and2b_1
X_11148_ _09135_/Y _11135_/X _11247_/B _09064_/Y _11146_/Y vssd1 vssd1 vccd1 vccd1
+ _11148_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11182__A1 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__B2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12131__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ _11297_/A fanout7/X fanout5/X _11169_/A vssd1 vssd1 vccd1 vccd1 _11080_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07310_ fanout36/X _12690_/A _07305_/X fanout92/X vssd1 vssd1 vccd1 vccd1 _07311_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07310__B1 _07305_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ _08698_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06664__A2 _06665_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ _09979_/A _07241_/B vssd1 vssd1 vccd1 vccd1 _07243_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07172_ _10252_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09063__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07613__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__B2 _06940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout304 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__buf_8
X_09813_ _11448_/A _09805_/X _09806_/Y _09812_/X vssd1 vssd1 vccd1 vccd1 _09813_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07019__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06956_ _10529_/A _10156_/A _06961_/B vssd1 vssd1 vccd1 vccd1 _06957_/B sky130_fd_sc_hd__nand3_1
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__or2_1
X_06887_ instruction[29] _06887_/B vssd1 vssd1 vccd1 vccd1 _06887_/X sky130_fd_sc_hd__or2_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _10117_/A _12141_/A fanout45/X _12684_/A vssd1 vssd1 vccd1 vccd1 _09676_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08341__A2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _08626_/A _08626_/B vssd1 vssd1 vccd1 vccd1 _08627_/B sky130_fd_sc_hd__and2_1
XFILLER_0_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08557_ _08472_/Y _08555_/A _08556_/Y _08422_/A vssd1 vssd1 vccd1 vccd1 _08846_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11228__A2 _11164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07730_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07689__A _07689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ _08219_/B _10506_/A _10647_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08489_/B
+ sky130_fd_sc_hd__o22a_1
X_07439_ _07439_/A _07439_/B vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _10450_/A _10450_/B _10450_/C vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__and3_1
XANTENNA__11936__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _09107_/X _09108_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09109_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10739__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10381_ _10490_/B2 fanout14/X fanout52/X fanout80/X vssd1 vssd1 vccd1 vccd1 _10382_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _12061_/A _12058_/Y _12060_/B vssd1 vssd1 vccd1 vccd1 _12124_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ _12051_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09357__B2 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__A1 _09885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11002_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11002_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12953_ hold78/X _12665_/A _12955_/B1 hold138/A _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold79/A sky130_fd_sc_hd__o221a_1
XFILLER_0_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _11905_/A _11905_/B _11905_/C vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__o21ai_4
X_12884_ _13062_/A hold232/X vssd1 vssd1 vccd1 vccd1 _13183_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _12110_/A _12110_/C _09621_/A vssd1 vssd1 vccd1 vccd1 _11836_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _06794_/X _11765_/X _12053_/A vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07843__A1 _12704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06934__C _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10717_ curr_PC[11] _10832_/C vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _11696_/A _11695_/Y _11696_/Y _09156_/B vssd1 vssd1 vccd1 vccd1 _11708_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07843__B2 _12706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08399__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ _10957_/A fanout11/X fanout44/X fanout81/X vssd1 vssd1 vccd1 vccd1 _10649_/B
+ sky130_fd_sc_hd__o22a_1
X_10579_ _09480_/X _09484_/X _11033_/A vssd1 vssd1 vccd1 vccd1 _10580_/A sky130_fd_sc_hd__mux2_1
X_12318_ _12499_/B _12319_/B vssd1 vssd1 vccd1 vccd1 _12326_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ _12250_/B _12250_/C _12250_/A vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06810_ _12175_/A _06809_/X _06819_/A vssd1 vssd1 vccd1 vccd1 _06810_/X sky130_fd_sc_hd__o21a_1
X_07790_ _07875_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__xnor2_1
X_06741_ _06739_/Y _06741_/B vssd1 vssd1 vccd1 vccd1 _06834_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09460_ _09283_/A _09283_/B _09459_/X vssd1 vssd1 vccd1 vccd1 _09460_/Y sky130_fd_sc_hd__a21oi_1
X_06672_ _06963_/A reg1_val[14] vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__and2b_1
X_08411_ _08411_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08412_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11863__C1 _11862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _09217_/A _09216_/Y _09220_/X vssd1 vssd1 vccd1 vccd1 _09396_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__B _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ _10853_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _06938_/A _06938_/B _08765_/A vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10647__B _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07224_ _07225_/A _07225_/B vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07155_ _07156_/A _07156_/B vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__nor2_8
XANTENNA_fanout301_A _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__B _06862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07086_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07087_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout101 _07165_/Y vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__buf_8
Xfanout112 _11887_/A vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout134 _07290_/X vssd1 vssd1 vccd1 vccd1 _12686_/A sky130_fd_sc_hd__buf_8
Xfanout145 _07137_/Y vssd1 vssd1 vccd1 vccd1 _08689_/B1 sky130_fd_sc_hd__buf_8
Xfanout156 _06952_/X vssd1 vssd1 vccd1 vccd1 _10853_/A sky130_fd_sc_hd__clkbuf_16
Xfanout123 _08430_/B vssd1 vssd1 vccd1 vccd1 _10852_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout189 _08698_/A vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__clkbuf_16
Xfanout167 _07056_/Y vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__buf_8
X_07988_ _08755_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__nor2_1
X_06939_ _06939_/A _10761_/A vssd1 vssd1 vccd1 vccd1 _06939_/X sky130_fd_sc_hd__or2_2
X_09727_ _09727_/A fanout3/X vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _12182_/B vssd1 vssd1 vccd1 vccd1 _09658_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A _07156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _08734_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08643_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10838__A _11799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _09590_/A _09590_/B vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__nor2_1
X_11620_ hold210/A _11620_/B _11701_/B vssd1 vssd1 vccd1 vccd1 _11620_/X sky130_fd_sc_hd__and3_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _12089_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _11555_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ fanout7/X fanout93/X _10647_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _10503_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ _12086_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11483_/B sky130_fd_sc_hd__xnor2_1
X_13221_ _13222_/CLK _13221_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10433_ _10433_/A _10433_/B vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__xnor2_1
X_13152_ _13250_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07589__B1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12103_ _12157_/B _12103_/B vssd1 vssd1 vccd1 vccd1 _12104_/C sky130_fd_sc_hd__or2_1
X_13083_ hold271/X _13082_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10161_/A _10160_/B _10158_/X vssd1 vssd1 vccd1 vccd1 _10297_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12034_ _11966_/A _11966_/B _11965_/A vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08002__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ _07301_/B _12962_/B2 hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__o21a_1
XFILLER_0_87_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10112__A2 _10370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ hold218/X _13070_/B2 _13070_/A2 hold184/X vssd1 vssd1 vccd1 vccd1 hold219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ _11819_/A _11819_/B _11819_/C vssd1 vssd1 vccd1 vccd1 _11902_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08069__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12798_ _12989_/B _12990_/A _12777_/X vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__a21o_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__A _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__A _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11749_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__and2_1
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07292__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06961__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06680__B _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _08962_/B sky130_fd_sc_hd__xnor2_1
X_07911_ _10398_/A _07911_/B vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__xnor2_2
X_08891_ fanout15/X _09885_/A _09880_/B2 _07513_/B vssd1 vssd1 vccd1 vccd1 _08892_/B
+ sky130_fd_sc_hd__o22a_1
X_07842_ _07842_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09741__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__B2 _10099_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09512_ _09467_/X _09469_/X _09511_/Y _06847_/X vssd1 vssd1 vccd1 vccd1 _09512_/X
+ sky130_fd_sc_hd__a31o_2
X_07773_ fanout81/X _06977_/A _06985_/A _06947_/X vssd1 vssd1 vccd1 vccd1 _07774_/B
+ sky130_fd_sc_hd__o22a_1
X_06724_ reg1_val[6] _07158_/A vssd1 vssd1 vccd1 vccd1 _06725_/B sky130_fd_sc_hd__nand2_1
X_06655_ instruction[26] _12498_/C vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ _09191_/A _09191_/B _09192_/X vssd1 vssd1 vccd1 vccd1 _09448_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ fanout49/X fanout92/X _12690_/A fanout51/X vssd1 vssd1 vccd1 vccd1 _09375_/B
+ sky130_fd_sc_hd__o22a_1
X_06586_ _06584_/X _06586_/B vssd1 vssd1 vccd1 vccd1 _12221_/A sky130_fd_sc_hd__and2b_1
X_08325_ _08714_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ _08196_/A _08196_/B _08194_/Y vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__A1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__B2 _08740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07207_ fanout82/X _10099_/A1 _12702_/A _06940_/A vssd1 vssd1 vccd1 vccd1 _07208_/B
+ sky130_fd_sc_hd__o22a_1
X_08187_ _08188_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08187_/Y sky130_fd_sc_hd__nand2b_1
X_07138_ _07138_/A _11727_/A vssd1 vssd1 vccd1 vccd1 _07138_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__11367__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11367__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07069_ _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__and2_2
XANTENNA__08798__A _09313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ hold285/A hold294/A _10080_/C vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__or3_1
XANTENNA__07991__B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10982_/A fanout4/X vssd1 vssd1 vccd1 vccd1 _10983_/C sky130_fd_sc_hd__nor2_1
X_12721_ hold31/X _12720_/B _12720_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__o211a_1
XANTENNA__09422__A _09422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12652_ _12646_/B _12648_/B _12646_/A vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_127_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ _11603_/A _11603_/B _11603_/C vssd1 vssd1 vccd1 vccd1 _11834_/B sky130_fd_sc_hd__and3_1
XFILLER_0_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ reg1_val[15] _12576_/B _12579_/A vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11534_ hold283/A _11623_/B _11622_/B _12313_/A1 vssd1 vssd1 vccd1 vccd1 _11534_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11465_ _11474_/A vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13204_ _13217_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 _13204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11358__A1 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__nor2_1
X_11396_ _11304_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__nand2b_1
X_13135_ _13260_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_10347_ hold279/A _12304_/B1 _10345_/X _09810_/A vssd1 vssd1 vccd1 vccd1 _10347_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ hold269/X _13070_/A2 _13065_/X _13070_/B2 vssd1 vssd1 vccd1 vccd1 hold270/A
+ sky130_fd_sc_hd__a22o_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ fanout71/X _11564_/A fanout38/X fanout77/X vssd1 vssd1 vccd1 vccd1 _10279_/B
+ sky130_fd_sc_hd__o22a_1
X_12017_ _11955_/A _07112_/B fanout4/X _11887_/A vssd1 vssd1 vccd1 vccd1 _12017_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ hold97/X _12662_/A _13112_/B hold150/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold158/A sky130_fd_sc_hd__o221a_1
XFILLER_0_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__B1 _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12243__C1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09478__S _09630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ _09088_/X _09089_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08110_ _08110_/A _08110_/B vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__xnor2_2
X_08041_ _08043_/A vssd1 vssd1 vccd1 vccd1 _08041_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08214__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _07157_/X _12029_/B _09870_/Y _09874_/Y vssd1 vssd1 vccd1 vccd1 _09993_/B
+ sky130_fd_sc_hd__a211o_1
X_08943_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08874_ _08045_/Y _08871_/Y _08873_/Y _07973_/X vssd1 vssd1 vccd1 vccd1 _08986_/B
+ sky130_fd_sc_hd__a211o_2
X_07825_ _07825_/A _07825_/B vssd1 vssd1 vccd1 vccd1 _07826_/B sky130_fd_sc_hd__and2_1
XANTENNA__07027__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _07756_/A _07756_/B _07756_/C vssd1 vssd1 vccd1 vccd1 _07883_/A sky130_fd_sc_hd__and3_1
X_06707_ reg2_val[8] _06748_/B vssd1 vssd1 vccd1 vccd1 _06707_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07687_ _09862_/B _07687_/B vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__xnor2_1
X_09426_ _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06638_ _06646_/A _12512_/B vssd1 vssd1 vccd1 vccd1 _06638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06569_ reg2_val[30] _06748_/B _06657_/B1 _06568_/X vssd1 vssd1 vccd1 vccd1 _07255_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _09885_/A _12141_/A fanout45/X _09880_/B2 vssd1 vssd1 vccd1 vccd1 _09358_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _09617_/B _09286_/Y _09287_/Y vssd1 vssd1 vccd1 vccd1 _09288_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07256__A2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _08308_/A _08308_/B vssd1 vssd1 vccd1 vccd1 _08310_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08239_ _08239_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08241_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10260__A1 _11295_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11781_/B _11348_/B hold184/A vssd1 vssd1 vccd1 vccd1 _11250_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09402__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09953__B2 _09293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _09630_/X _09634_/B _10201_/S vssd1 vssd1 vccd1 vccd1 _10201_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08756__A2 _08782_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _11308_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11760__A1 _12110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _10132_/A _10275_/A _10132_/C vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09705__A1 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _09931_/A _09928_/Y _09930_/B vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09705__B2 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _12704_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12704_/Y sky130_fd_sc_hd__nand2_1
X_10965_ _11656_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13017__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ _10896_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ _12635_/A _12640_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
X_12566_ _12566_/A _12574_/A vssd1 vssd1 vccd1 vccd1 _12568_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _11838_/A _09045_/B _09045_/C _09146_/X vssd1 vssd1 vccd1 vccd1 _11517_/X
+ sky130_fd_sc_hd__a31o_1
X_12497_ _12497_/A _12497_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _11448_/A _11448_/B _11448_/C vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__or3_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _11491_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13118_ _13121_/A _13118_/B _13118_/C vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__and3_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13049_/A _13049_/B vssd1 vssd1 vccd1 vccd1 _13050_/B sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07610_ _06963_/Y fanout43/X _07239_/A fanout80/X vssd1 vssd1 vccd1 vccd1 _07611_/B
+ sky130_fd_sc_hd__o22a_1
X_08590_ _08590_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__nand2_1
X_07541_ _07541_/A _07541_/B vssd1 vssd1 vccd1 vccd1 _07543_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11267__B1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07472_ _07538_/A _07538_/B _07437_/Y vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09880__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _09235_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10490__B2 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__A1 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10447__D_N _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ _09151_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__or2_4
XANTENNA__08435__A1 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08435__B2 _10876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ reg1_val[7] reg1_val[24] _09092_/S vssd1 vssd1 vccd1 vccd1 _09073_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout214_A _06890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout3 fanout4/X vssd1 vssd1 vccd1 vccd1 fanout3/X sky130_fd_sc_hd__clkbuf_8
X_08024_ _08257_/A _08257_/B _08023_/A vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09237__A _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A2 _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__nand2b_1
X_08926_ _09422_/A fanout17/X fanout9/X _09222_/B2 vssd1 vssd1 vccd1 vccd1 _08927_/B
+ sky130_fd_sc_hd__o22a_1
X_08857_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__nand2_1
X_07808_ _07808_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _07813_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10702__C1 _12303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08788_ _08814_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__xnor2_1
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10750_ _10638_/X _10644_/A _07277_/X _12029_/B vssd1 vssd1 vccd1 vccd1 _10890_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _11231_/B sky130_fd_sc_hd__nor2_1
X_09409_ fanout82/X fanout74/X fanout68/X _06940_/A vssd1 vssd1 vccd1 vccd1 _09410_/B
+ sky130_fd_sc_hd__o22a_1
X_12420_ _12576_/B _12421_/B vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _12522_/B _12351_/B vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__or2_1
XANTENNA__06988__A1 _06977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _12276_/Y _12277_/X _12281_/X _12274_/X vssd1 vssd1 vccd1 vccd1 _12282_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06988__B2 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _11302_/A _11302_/B vssd1 vssd1 vccd1 vccd1 _11303_/B sky130_fd_sc_hd__nand2_1
X_11233_ _11233_/A _11233_/B vssd1 vssd1 vccd1 vccd1 _11233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__nand2_1
X_10115_ _10115_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__and2_1
X_11095_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__xnor2_4
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11997_ _11994_/Y _11995_/X _11996_/Y vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__B1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948_ _10948_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10950_/C sky130_fd_sc_hd__and2_1
XANTENNA__10472__A1 _07289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _10996_/B _10878_/B _10878_/C vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ reg1_val[24] _12656_/A vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10224__A1 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ _12550_/A _12550_/C _12550_/B vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 curr_PC[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12690__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10491__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ reg1_val[7] _06970_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _06973_/B sky130_fd_sc_hd__o21a_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09760_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__xnor2_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__xnor2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _09587_/A _09587_/B _09583_/X vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08642_ _08755_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__or2_1
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout164_A _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _08734_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08605_/B sky130_fd_sc_hd__xnor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07524_/A _07524_/B vssd1 vssd1 vccd1 vccd1 _07525_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07455_ _12714_/A _09422_/A _09222_/B2 _12716_/A vssd1 vssd1 vccd1 vccd1 _07456_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07386_ _07389_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07391_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08136__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _09123_/X _09124_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09056_ _12178_/A _09056_/B _09056_/C _09055_/Y vssd1 vssd1 vccd1 vccd1 _12223_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08007_ _10876_/A1 _08699_/A2 fanout93/X _08670_/A2 vssd1 vssd1 vccd1 vccd1 _08008_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11715__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _11153_/A _09958_/B _10092_/B vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__or3_1
XANTENNA_fanout77_A _06983_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _09725_/B2 fanout63/X _11950_/A _10009_/A vssd1 vssd1 vccd1 vccd1 _08910_/B
+ sky130_fd_sc_hd__o22a_1
X_09889_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__or2_1
XANTENNA__12691__A2 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _11849_/A _11849_/B _11847_/B vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__o21a_1
XANTENNA__10151__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ hold291/A _11931_/C vssd1 vssd1 vccd1 vccd1 _11851_/X sky130_fd_sc_hd__or2_1
X_11782_ _09501_/B _11625_/B _11782_/S vssd1 vssd1 vccd1 vccd1 _11782_/X sky130_fd_sc_hd__mux2_1
X_10802_ _10692_/A _10690_/X _10706_/S vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__A _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ _10733_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11651__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10664_ _10520_/A _10520_/B _10518_/Y vssd1 vssd1 vccd1 vccd1 _10666_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _12403_/A _12403_/B _12403_/C vssd1 vssd1 vccd1 vccd1 _12404_/B sky130_fd_sc_hd__nand3_1
X_10595_ _12303_/A _10582_/X _10594_/X _10571_/X vssd1 vssd1 vccd1 vccd1 _10595_/X
+ sky130_fd_sc_hd__o211a_1
X_12334_ _12340_/B _12334_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11706__B2 _09330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ _12264_/A _12264_/B _12264_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _12265_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _12170_/Y _12171_/X _12179_/Y _12195_/X vssd1 vssd1 vccd1 vccd1 _12196_/X
+ sky130_fd_sc_hd__a211o_1
X_11216_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11218_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _10809_/A _09128_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11182__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _12089_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__xnor2_1
X_10029_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07310__B2 fanout92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07310__A1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _12694_/A fanout42/X _07239_/A _10490_/B2 vssd1 vssd1 vccd1 vccd1 _07241_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07171_ fanout77/X _06985_/A _12706_/A _06977_/A vssd1 vssd1 vccd1 vccd1 _07172_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09063__A1 _09464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__B2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__A1 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09486__S _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__B2 _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10933__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__A2 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout305 instruction[7] vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__buf_4
X_09812_ _06739_/Y _09138_/X _09501_/B _06834_/A _09811_/X vssd1 vssd1 vccd1 vccd1
+ _09812_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10381__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__B _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _12498_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08326__B1 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ _10529_/A _06961_/B vssd1 vssd1 vccd1 vccd1 _06955_/Y sky130_fd_sc_hd__nand2_1
X_09743_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__nand2_1
X_06886_ instruction[21] _06850_/Y _06885_/X _06637_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__o211a_4
X_09674_ _09567_/A _09567_/B _09565_/Y vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__a21o_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08625_ _08625_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08647_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08556_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08629__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _07507_/A _07507_/B vssd1 vssd1 vccd1 vccd1 _07730_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08629__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08487_ _08490_/A _08490_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__or2_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07438_ _07438_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07439_/B sky130_fd_sc_hd__and2_1
XFILLER_0_52_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _07369_/A _07369_/B vssd1 vssd1 vccd1 vccd1 _07397_/B sky130_fd_sc_hd__and2_1
X_09108_ reg1_val[15] reg1_val[16] _09120_/S vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10739__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ _11458_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09039_ _11426_/B _09039_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__or3_1
X_12050_ _09465_/A _09056_/B _09056_/C _12179_/A vssd1 vssd1 vccd1 vccd1 _12051_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09357__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _11003_/A _11003_/B vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__nand2_1
X_12952_ _07112_/B _12962_/B2 hold107/X vssd1 vssd1 vccd1 vccd1 _13217_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10124__B1 _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _11973_/B _11903_/B vssd1 vssd1 vccd1 vccd1 _11905_/C sky130_fd_sc_hd__and2_1
X_12883_ hold220/X _13070_/B2 _13070_/A2 hold231/X vssd1 vssd1 vccd1 vccd1 hold232/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11834_ _11834_/A _11834_/B _11834_/C _11834_/D vssd1 vssd1 vccd1 vccd1 _12110_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11689_/A _11687_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11696_/A _11696_/B vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07843__A2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716_ _10684_/Y _10685_/X _10688_/X _10715_/X vssd1 vssd1 vccd1 vccd1 _10716_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _10647_/A _11296_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ _12125_/S _10578_/B vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__nand2_1
X_12317_ _12499_/A curr_PC[0] _12444_/S vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12248_ _12728_/A _12248_/B _12248_/C vssd1 vssd1 vccd1 vccd1 _12250_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12179_ _12179_/A _12179_/B vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06678__B _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ reg1_val[4] _07108_/C vssd1 vssd1 vccd1 vccd1 _06741_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06671_ _06763_/B _06613_/A _12576_/B _06670_/X vssd1 vssd1 vccd1 vccd1 _06963_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08410_ _08410_/A _08410_/B vssd1 vssd1 vccd1 vccd1 _08474_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09390_ _09600_/B _09390_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09284__A1 _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ fanout79/X _09237_/A _09428_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08342_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _08272_/A _08272_/B _08272_/C vssd1 vssd1 vccd1 vccd1 _08272_/X sky130_fd_sc_hd__and3_1
XANTENNA__10969__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07223_ _07832_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07225_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09036__A1 _09001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ _07156_/A _07156_/B _11799_/A vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_30_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07085_ reg1_val[14] reg1_val[15] vssd1 vssd1 vccd1 vccd1 _07091_/C sky130_fd_sc_hd__or2_2
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__A2 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 _11887_/A vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__buf_8
Xfanout102 _11470_/A vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout135 _11068_/A vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__buf_12
Xfanout146 _07122_/X vssd1 vssd1 vccd1 vccd1 _08715_/A2 sky130_fd_sc_hd__buf_6
Xfanout124 _06961_/Y vssd1 vssd1 vccd1 vccd1 _08430_/B sky130_fd_sc_hd__buf_8
Xfanout168 _09727_/A vssd1 vssd1 vccd1 vccd1 _08782_/A2 sky130_fd_sc_hd__buf_6
X_07987_ _08022_/A _07987_/B _07987_/C vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__nand3_1
Xfanout179 _08607_/A vssd1 vssd1 vccd1 vccd1 _10607_/A sky130_fd_sc_hd__buf_12
Xfanout157 _08535_/A vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__buf_8
XANTENNA__06588__B _12565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__nand2_4
XANTENNA__10106__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _10126_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__xor2_1
X_06869_ instruction[18] _06887_/B vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__or2_1
X_09657_ _10809_/A _09656_/X _09159_/Y vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09434_/A _09433_/B _09433_/A vssd1 vssd1 vccd1 vccd1 _09590_/B sky130_fd_sc_hd__a21boi_2
X_08608_ _08219_/B _08715_/A2 _08689_/B1 _08815_/B vssd1 vssd1 vccd1 vccd1 _08609_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08539_ _08539_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ fanout64/X fanout11/X fanout44/X _11876_/A vssd1 vssd1 vccd1 vccd1 _11551_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _10400_/A _10399_/B _10399_/A vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__o21ba_1
X_13220_ _13222_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ _11876_/A fanout14/X fanout52/X _11950_/A vssd1 vssd1 vccd1 vccd1 _11482_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07589__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10433_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13151_ _13250_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07589__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10363_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__nand2_1
X_13082_ _13082_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13082_/Y sky130_fd_sc_hd__xnor2_1
X_12102_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12103_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _12104_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__nand2_1
X_10294_ _10146_/A _10146_/C _10146_/B vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_109_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08002__A2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__A1 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ hold39/X _12665_/A _12955_/B1 _13209_/Q _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold40/A sky130_fd_sc_hd__o221a_1
XFILLER_0_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10648__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ _13062_/A hold172/X vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11895_/B _11817_/B vssd1 vssd1 vccd1 vccd1 _11819_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08069__A2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ _12781_/B _12985_/B _12779_/X vssd1 vssd1 vccd1 vccd1 _12990_/A sky130_fd_sc_hd__a21o_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ _11828_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _11757_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__B _06961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07910_ _10876_/A1 _08670_/A2 _08699_/A2 _10957_/A vssd1 vssd1 vccd1 vccd1 _07911_/B
+ sky130_fd_sc_hd__o22a_1
X_08890_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09065__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _06828_/A _12714_/A _08765_/A _12712_/A vssd1 vssd1 vccd1 vccd1 _07842_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09741__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _07782_/B _07854_/A _07782_/A vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__o21a_1
X_06723_ reg1_val[6] _07158_/A vssd1 vssd1 vccd1 vccd1 _06723_/Y sky130_fd_sc_hd__nor2_1
X_09511_ _09136_/B _09506_/X _09510_/X vssd1 vssd1 vccd1 vccd1 _09511_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06654_ instruction[0] instruction[1] _06850_/B instruction[26] pred_val vssd1 vssd1
+ vccd1 vccd1 _12502_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ _09268_/A _09268_/B _09267_/A vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__o21ai_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06585_ reg1_val[29] _06585_/B vssd1 vssd1 vccd1 vccd1 _06586_/B sky130_fd_sc_hd__or2_1
XANTENNA__07313__A _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout244_A _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08324_ _08670_/A2 _08715_/A2 _08689_/B1 _08699_/A2 vssd1 vssd1 vccd1 vccd1 _08325_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06871__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08255_ _08163_/A _08162_/B _08162_/A vssd1 vssd1 vccd1 vccd1 _08261_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__08480__A2 _08715_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _08186_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08188_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ _07137_/A _07137_/B vssd1 vssd1 vccd1 vccd1 _07137_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__11367__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10393__B _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07440__B1 _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _07068_/A _07068_/B vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__nand2_8
XANTENNA__12316__A1 _07184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__B _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07991__B2 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10981_ _06955_/Y fanout4/X _10156_/A vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__o21a_1
X_09709_ fanout83/X fanout65/X fanout58/X _06940_/A vssd1 vssd1 vccd1 vccd1 _09710_/B
+ sky130_fd_sc_hd__o22a_1
X_12720_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09422__B fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07223__A _07832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _11602_/A vssd1 vssd1 vccd1 vccd1 _11834_/A sky130_fd_sc_hd__inv_2
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12582_ _12584_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__nor2_2
X_11533_ _11623_/B _11622_/B hold283/A vssd1 vssd1 vccd1 vccd1 _11533_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12004__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ _11579_/B _11464_/B vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13203_ _13208_/CLK _13203_/D vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11395_ _11395_/A _11395_/B vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _12304_/B1 _10345_/X hold279/A vssd1 vssd1 vccd1 vccd1 _10346_/Y sky130_fd_sc_hd__a21oi_1
X_13134_ _13222_/CLK _13134_/D vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ hold263/X _13064_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__mux2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _11271_/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10281_/A sky130_fd_sc_hd__xnor2_1
X_12016_ _12142_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13169_/CLK sky130_fd_sc_hd__clkbuf_8
X_12918_ _10398_/A _12926_/A2 hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__o21a_1
XANTENNA__06956__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07133__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09239__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ hold213/X _12885_/A2 _12885_/B1 hold241/X vssd1 vssd1 vccd1 vccd1 hold242/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06691__B _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ _08042_/A _08042_/B _08042_/C vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08214__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09991_ _09870_/Y _09874_/Y _07157_/X _12029_/B vssd1 vssd1 vccd1 vccd1 _09991_/X
+ sky130_fd_sc_hd__o211a_1
X_08942_ _08942_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ _09055_/A _08988_/A _08987_/B _08041_/Y _07974_/X vssd1 vssd1 vccd1 vccd1
+ _08873_/Y sky130_fd_sc_hd__o32ai_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _07824_/A _07824_/B vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07755_ _07811_/B _07752_/B _07750_/X vssd1 vssd1 vccd1 vccd1 _07756_/C sky130_fd_sc_hd__o21bai_2
X_06706_ _06704_/Y _06706_/B vssd1 vssd1 vccd1 vccd1 _06830_/C sky130_fd_sc_hd__nand2b_1
X_07686_ _06983_/Y _09727_/A _08798_/B _12710_/A vssd1 vssd1 vccd1 vccd1 _07687_/B
+ sky130_fd_sc_hd__o22a_1
X_06637_ instruction[28] _06637_/B vssd1 vssd1 vccd1 vccd1 _12512_/B sky130_fd_sc_hd__and2_4
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08139__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09425_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06568_ _06613_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _06568_/X sky130_fd_sc_hd__or2_1
XFILLER_0_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ _09356_/A _09356_/B vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09287_ _09617_/B _09286_/Y _09061_/X vssd1 vssd1 vccd1 vccd1 _09287_/Y sky130_fd_sc_hd__a21oi_1
X_08307_ _08307_/A _08307_/B vssd1 vssd1 vccd1 vccd1 _08308_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08238_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__and2_1
XFILLER_0_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10260__A2 _07988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ _10198_/X _10199_/X _11134_/S vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__mux2_1
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08170_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09402__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ _11180_/A _11180_/B _11180_/C vssd1 vssd1 vccd1 vccd1 _11181_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10130_/B _10130_/C _10130_/A vssd1 vssd1 vccd1 vccd1 _10132_/C sky130_fd_sc_hd__a21o_1
X_10062_ _06832_/A _10060_/X _10061_/Y vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__09705__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ hold5/X _12730_/B _12702_/Y _13080_/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__o211a_1
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08049__A _10853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ fanout64/X fanout50/X _07988_/B _11876_/A vssd1 vssd1 vccd1 vccd1 _10965_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13017__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ _11003_/B _10895_/B vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__and2_1
X_12634_ reg1_val[27] _12656_/A vssd1 vssd1 vccd1 vccd1 _12640_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12565_ reg1_val[13] _12565_/B vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _11838_/A _09045_/B _09045_/C vssd1 vssd1 vccd1 vccd1 _11516_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12497_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _10208_/B _11529_/B hold182/A vssd1 vssd1 vccd1 vccd1 _11448_/C sky130_fd_sc_hd__a21oi_1
X_11378_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__or2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10761__B _11385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ hold164/X hold100/X hold161/X vssd1 vssd1 vccd1 vccd1 _13118_/C sky130_fd_sc_hd__a21o_1
X_10329_ _06717_/A _10189_/X _06719_/B vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__o21a_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13085_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _13240_/D sky130_fd_sc_hd__and2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _07540_/A _07540_/B vssd1 vssd1 vccd1 vccd1 _07543_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06686__B _07278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07471_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07538_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09880__A1 _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__B2 _09880_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _09210_/A _09210_/B vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10490__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _09151_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _09141_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ _09068_/X _09071_/X _09630_/S vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08435__A2 _10957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08257_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout4 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__buf_6
XANTENNA_fanout207_A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09237__B _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _09194_/B _08925_/B vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09699__A1 _09564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _07816_/A _07816_/B vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09253__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _06511_/Y _08765_/B _08765_/C _08765_/A _09568_/A vssd1 vssd1 vccd1 vccd1
+ _08788_/B sky130_fd_sc_hd__o32a_2
X_07738_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout22_A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _10680_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__xnor2_4
X_09408_ _09979_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__xnor2_1
X_09339_ _12115_/A _12668_/A _09337_/Y _12265_/C1 vssd1 vssd1 vccd1 vccd1 _09340_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11023__A _11238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _12522_/B _12351_/B vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06988__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12281_ _09330_/A _09293_/B _09324_/Y _09293_/A _12280_/Y vssd1 vssd1 vccd1 vccd1
+ _12281_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _11301_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__or2_1
XFILLER_0_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _11232_/A _12110_/A vssd1 vssd1 vccd1 vccd1 _11233_/B sky130_fd_sc_hd__or2_1
XANTENNA__09428__A _09428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12930__A1 _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _11163_/A _11163_/B _11163_/C _08982_/A vssd1 vssd1 vccd1 vccd1 _11164_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__11194__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _10115_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10941__B1 _10940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11094_ _11094_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__and2_1
XANTENNA__08986__B _08986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
X_11996_ _12302_/A _10088_/Y _12303_/A vssd1 vssd1 vccd1 vccd1 _11996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__B2 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__B2 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ _10867_/A _10867_/B _10864_/A vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10472__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ reg1_val[24] _12656_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _10996_/B _10878_/B _10878_/C vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__and3_1
XFILLER_0_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12029__A _12095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ _12544_/A _12548_/B vssd1 vssd1 vccd1 vccd1 _12550_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12479_ _12465_/B _12473_/B _12484_/A vssd1 vssd1 vccd1 vccd1 _12480_/D sky130_fd_sc_hd__o21ai_1
XANTENNA_2 curr_PC[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__B1 _12313_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ reg1_val[7] _06971_/B vssd1 vssd1 vccd1 vccd1 _06971_/X sky130_fd_sc_hd__xor2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__nand2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09559_/A _09559_/B _09555_/Y vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__o21ai_2
X_08641_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08652_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08572_ _08219_/B _08689_/B1 _09180_/B2 _08815_/B vssd1 vssd1 vccd1 vccd1 _08573_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _07533_/A _07671_/A _07533_/C vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07454_ _07458_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout157_A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07385_ _09862_/B _07385_/B vssd1 vssd1 vccd1 vccd1 _07389_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ reg1_val[7] reg1_val[24] _09124_/S vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10215__A2 _09501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _09055_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08006_ _08010_/A _08010_/B vssd1 vssd1 vccd1 vccd1 _08006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11715__A2 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09957_ curr_PC[4] curr_PC[5] _09957_/C vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__and3_1
X_08908_ _10607_/A _08908_/B vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _09888_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10151__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__A1 _11739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ _09029_/B _09030_/A _08621_/X vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__a21o_1
X_11850_ _10350_/Y _11849_/Y _12271_/S vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ hold191/A _11781_/B _11854_/B vssd1 vssd1 vccd1 vccd1 _11781_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12979__B2 _13110_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ _11232_/A _10800_/C _10800_/B vssd1 vssd1 vccd1 vccd1 _10801_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_95_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11651__A1 _07069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _10733_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08327__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11651__B2 _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ _10663_/A _10663_/B vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__or2_1
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _12403_/A _12403_/B _12403_/C vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__a21o_1
X_10594_ _12073_/B2 _10581_/X _11696_/B _09124_/S _10592_/X vssd1 vssd1 vccd1 vccd1
+ _10594_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12333_ _12333_/A _12333_/B _12333_/C vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12264_ _12264_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12264_/Y sky130_fd_sc_hd__nand2_1
X_12195_ _12195_/A _12195_/B _12195_/C _12195_/D vssd1 vssd1 vccd1 vccd1 _12195_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11215_ _11104_/A _11104_/B _11103_/A vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11138_/Y _11139_/X _11145_/X vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11077_ _11295_/B2 fanout11/X fanout44/X _11462_/A vssd1 vssd1 vccd1 vccd1 _11078_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10028_ _10028_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09621__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10848__B1_N _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__B1 _07041_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _11909_/Y _11910_/X _12112_/A vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07310__A2 _12690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07170_ _07174_/A _07174_/B vssd1 vssd1 vccd1 vccd1 _07170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06980__A _06980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__A2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11945__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07287__S _07875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09811_ _06737_/Y _06905_/Y _09148_/X _06741_/B _09810_/X vssd1 vssd1 vccd1 vccd1
+ _09811_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout306 instruction[7] vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__buf_4
XANTENNA__10381__A1 _10490_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _11654_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08700__A _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__B2 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A1 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06954_ _10529_/A _10156_/A _06961_/B vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__or3_1
X_06885_ instruction[28] _06887_/B vssd1 vssd1 vccd1 vccd1 _06885_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout274_A _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _09605_/A _09605_/B _09606_/Y vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__a21bo_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08651_/A sky130_fd_sc_hd__nor2_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08555_/A vssd1 vssd1 vccd1 vccd1 _08555_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07507_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08629__A2 _08735_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08486_ _08814_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08490_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13234_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12892__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07437_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ _07368_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11936__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ reg1_val[14] reg1_val[17] _09120_/S vssd1 vssd1 vccd1 vccd1 _09107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07299_ _11271_/A _07301_/B vssd1 vssd1 vccd1 vccd1 _07305_/A sky130_fd_sc_hd__and2_1
XFILLER_0_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ _09039_/B _09039_/C vssd1 vssd1 vccd1 vccd1 _11426_/C sky130_fd_sc_hd__or2_1
XFILLER_0_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08014__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _11000_/A _11000_/B vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09706__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ hold106/X _12662_/A _12955_/B1 hold78/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold107/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12882_ _13071_/A hold221/X vssd1 vssd1 vccd1 vccd1 _13182_/D sky130_fd_sc_hd__and2_1
X_11902_ _11902_/A _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__or3_1
X_11833_ _11833_/A _11833_/B vssd1 vssd1 vccd1 vccd1 _12110_/B sky130_fd_sc_hd__xnor2_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ _11838_/A _09052_/B _09052_/C _09146_/X vssd1 vssd1 vccd1 vccd1 _11764_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11695_/A _11695_/B vssd1 vssd1 vccd1 vccd1 _11695_/Y sky130_fd_sc_hd__xnor2_1
X_10715_ _10715_/A _10715_/B _10715_/C vssd1 vssd1 vccd1 vccd1 _10715_/X sky130_fd_sc_hd__and3_1
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10646_ _11296_/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ _10577_/A _10577_/B _10577_/C vssd1 vssd1 vccd1 vccd1 _10578_/B sky130_fd_sc_hd__or3_1
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _07184_/B _06905_/Y _12294_/X _12315_/Y _12080_/A vssd1 vssd1 vccd1 vccd1
+ dest_val[31] sky130_fd_sc_hd__o221a_4
XFILLER_0_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12247_ _12728_/A _12246_/X _12248_/C vssd1 vssd1 vccd1 vccd1 _12250_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12178_ _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__xnor2_1
X_11129_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ reg2_val[14] _06748_/B vssd1 vssd1 vccd1 vccd1 _06670_/X sky130_fd_sc_hd__and2_1
XANTENNA__12696__B _12730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__A _08698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__B2 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _08607_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _11072_/A _08271_/B vssd1 vssd1 vccd1 vccd1 _08272_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ fanout77/X _07000_/A _12706_/A _10481_/A vssd1 vssd1 vccd1 vccd1 _07223_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07153_ _07150_/Y _07152_/X _11726_/A vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09543__A_N _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ _07339_/A _07339_/B _07024_/Y vssd1 vssd1 vccd1 vccd1 _07204_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 _11470_/A vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__buf_6
XANTENNA__06869__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout114 _08642_/B vssd1 vssd1 vccd1 vccd1 _07000_/A sky130_fd_sc_hd__buf_6
Xfanout147 _07122_/X vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__buf_6
Xfanout125 _12694_/A vssd1 vssd1 vccd1 vccd1 _10876_/A1 sky130_fd_sc_hd__buf_8
Xfanout136 _07282_/X vssd1 vssd1 vccd1 vccd1 _11068_/A sky130_fd_sc_hd__buf_12
XANTENNA__08430__A _08755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 _07054_/X vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__buf_8
X_07986_ _07984_/A _07984_/C _07984_/B vssd1 vssd1 vccd1 vccd1 _07987_/C sky130_fd_sc_hd__a21o_1
Xfanout158 _08535_/A vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__buf_4
XFILLER_0_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07046__A _09423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06937_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _06937_/X sky130_fd_sc_hd__and2_1
XANTENNA__10106__A1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10106__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _10009_/A fanout17/X fanout9/A _09725_/B2 vssd1 vssd1 vccd1 vccd1 _09726_/B
+ sky130_fd_sc_hd__o22a_1
X_09656_ _11033_/A _09655_/X _09166_/B vssd1 vssd1 vccd1 vccd1 _09656_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_69_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06868_ instruction[15] _06868_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _08607_/A _08607_/B vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__xnor2_1
X_06799_ _06798_/X _06839_/A vssd1 vssd1 vccd1 vccd1 _06799_/X sky130_fd_sc_hd__and2b_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09587_/A _09587_/B vssd1 vssd1 vccd1 vccd1 _09590_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08539_/B sky130_fd_sc_hd__and2_1
XFILLER_0_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _08427_/X _08510_/A vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08483__B1 _09180_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _10500_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ _11480_/A _11480_/B vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10431_ _10429_/A _10429_/B _10432_/B vssd1 vssd1 vccd1 vccd1 _10431_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _13250_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__A2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _11470_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13081_ _12743_/X _13081_/B vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11790__B1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12157_/B sky130_fd_sc_hd__o21a_1
X_10293_ _10111_/A _10111_/B _10109_/Y vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__a21o_1
X_12032_ _12032_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__or2_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08340__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ _09979_/A _12962_/B2 hold84/X vssd1 vssd1 vccd1 vccd1 _13208_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_88_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12865_ hold171/X _13070_/B2 _13070_/A2 hold218/A vssd1 vssd1 vccd1 vccd1 hold172/A
+ sky130_fd_sc_hd__a22o_1
X_12796_ _12784_/B _12981_/B _12782_/X vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__a21o_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11816_ _11816_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__and2_1
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ _11747_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__or2_1
XANTENNA__12963__C fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11757_/B _11678_/B vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__or2_2
XFILLER_0_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ _11295_/B2 fanout13/X fanout47/X _11462_/A vssd1 vssd1 vccd1 vccd1 _10630_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11876__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ _07929_/A _07838_/X _07835_/X vssd1 vssd1 vccd1 vccd1 _07850_/B sky130_fd_sc_hd__o21a_1
X_07771_ _07771_/A _07771_/B _07771_/C vssd1 vssd1 vccd1 vccd1 _07854_/A sky130_fd_sc_hd__and3_1
X_06722_ _07158_/A reg1_val[6] vssd1 vssd1 vccd1 vccd1 _06772_/A sky130_fd_sc_hd__nand2b_1
X_09510_ _09156_/B _09507_/X _09509_/X _09498_/Y vssd1 vssd1 vccd1 vccd1 _09510_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06653_ _06653_/A _06653_/B vssd1 vssd1 vccd1 vccd1 _11339_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ _09441_/A _09441_/B vssd1 vssd1 vccd1 vccd1 _09454_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06584_ reg1_val[29] _06585_/B vssd1 vssd1 vccd1 vccd1 _06584_/X sky130_fd_sc_hd__and2_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _09372_/A _09372_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10020__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08323_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout237_A _06737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08254_ _08198_/A _08198_/B _08199_/Y vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07205_ _07204_/B _07205_/B vssd1 vssd1 vccd1 vccd1 _07206_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08217__B1 _12702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 _12080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08185_ _08113_/Y _08120_/B _08118_/Y vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__a21oi_4
X_07136_ _07109_/A _06932_/C _07303_/A vssd1 vssd1 vccd1 vccd1 _07137_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09965__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10393__C _10845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__A1 _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _07067_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _07068_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07440__B2 _09237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ _07969_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _08039_/B sky130_fd_sc_hd__xnor2_1
X_09708_ _10398_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout52_A _07513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _11271_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__xnor2_1
X_09639_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ reg1_val[30] _12656_/A vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _11679_/B _11601_/B vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ reg1_val[16] _12615_/B vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__and2_1
X_11532_ hold287/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10076__S _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08208__B1 _08689_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _11462_/A _12245_/B _11462_/C vssd1 vssd1 vccd1 vccd1 _11464_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _13222_/CLK _13202_/D vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10015__B1 _07763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13222_/CLK _13133_/D vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11696__A _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _11394_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11395_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ hold300/A _10469_/C vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__or2_1
X_13064_ _13064_/A _13064_/B vssd1 vssd1 vccd1 vccd1 _13064_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08070__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ fanout65/X fanout42/X _07239_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _10277_/B
+ sky130_fd_sc_hd__o22a_1
X_12015_ _12201_/A fanout11/X _07391_/B fanout9/A vssd1 vssd1 vccd1 vccd1 _12016_/B
+ sky130_fd_sc_hd__o22a_1
X_12917_ _13199_/Q _12662_/A _13112_/B hold97/X _12955_/C1 vssd1 vssd1 vccd1 vccd1
+ hold98/A sky130_fd_sc_hd__o221a_1
XFILLER_0_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__C _06961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12848_ _13071_/A hold214/X vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__and2_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ hold51/X hold294/A vssd1 vssd1 vccd1 vccd1 _12779_/X sky130_fd_sc_hd__and2b_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08447__B1 _08735_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ _09865_/A _09865_/B _09864_/A vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__o21ai_4
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _08863_/B _08991_/B _08861_/X vssd1 vssd1 vccd1 vccd1 _08987_/B sky130_fd_sc_hd__a21o_1
X_07823_ _07823_/A _07823_/B _07823_/C vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__and3_1
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _07754_/A _07754_/B vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06705_ reg1_val[9] _06931_/B vssd1 vssd1 vccd1 vccd1 _06706_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07324__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ _07695_/B _07695_/C _07695_/A vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11690__C1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06636_ _11535_/A _06636_/B vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__and2_1
XFILLER_0_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__xor2_2
X_06567_ instruction[40] _12498_/C vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__and2_4
X_09355_ _09277_/A _09277_/B _09278_/Y vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08438__B1 _10647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ _09464_/A _10320_/A _09465_/A vssd1 vssd1 vccd1 vccd1 _09286_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _08306_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__A2 _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _08246_/B _08246_/A vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08168_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__A2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ _07149_/A _07149_/B vssd1 vssd1 vccd1 vccd1 _07119_/X sky130_fd_sc_hd__and2_1
X_08099_ _08207_/B _08207_/A vssd1 vssd1 vccd1 vccd1 _08099_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08610__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10130_ _10130_/A _10130_/B _10130_/C vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _06832_/A _10060_/X _12265_/C1 vssd1 vssd1 vccd1 vccd1 _10061_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10720__A1 _11636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ _11068_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__xnor2_1
X_12702_ _12702_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _12702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ _10894_/A _10894_/B _10894_/C vssd1 vssd1 vccd1 vccd1 _10895_/B sky130_fd_sc_hd__or3_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _12629_/A _12632_/B _12629_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ reg1_val[13] _12565_/B vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _12223_/A _11514_/C _11514_/B vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ reg1_val[27] curr_PC[27] _12495_/S vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ hold182/A _11620_/B _11529_/B vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__and3_1
XFILLER_0_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ hold161/X _12663_/B _12658_/Y _12664_/A vssd1 vssd1 vccd1 vccd1 _13118_/B
+ sky130_fd_sc_hd__a22o_1
X_10328_ _12263_/S _10328_/B _10328_/C vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__or3_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ hold298/X _13084_/A2 _13046_/X _13084_/B2 vssd1 vssd1 vccd1 vccd1 _13048_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07168__B1 _12712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10259_ _12086_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10711__A1 _07304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07470_ _07468_/A _07468_/B _07469_/Y vssd1 vssd1 vccd1 vccd1 _07538_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09880__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09140_ _09146_/A _09140_/B vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__or2_4
XFILLER_0_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09071_ _09069_/X _09070_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _08022_/A _08160_/A _08022_/C vssd1 vssd1 vccd1 vccd1 _08023_/B sky130_fd_sc_hd__and3_1
XFILLER_0_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout5 fanout6/X vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout102_A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06749__A3 _12512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09973_ _09857_/A _09856_/B _09854_/Y vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__a21o_2
XANTENNA__06750__A_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ _08924_/A _08924_/B vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07159__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A1 _11696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _08855_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08858_/B sky130_fd_sc_hd__nor2_2
XANTENNA__06906__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _07804_/A _07804_/B _07805_/Y vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__o21ai_2
X_08786_ _09423_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _08799_/A sky130_fd_sc_hd__xnor2_1
X_07737_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07668_ _07668_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06619_ _11704_/S _06619_/B vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__nor2_1
X_07599_ _07609_/A vssd1 vssd1 vccd1 vccd1 _07599_/Y sky130_fd_sc_hd__inv_2
X_09407_ _11297_/A fanout42/X _07239_/A _11295_/B2 vssd1 vssd1 vccd1 vccd1 _09408_/B
+ sky130_fd_sc_hd__o22a_1
X_09338_ _11238_/A _12668_/A _09337_/Y vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09084__A0 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09269_ _08964_/A _08963_/B _08961_/Y vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _11301_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__nand2_1
X_12280_ _12280_/A _12280_/B vssd1 vssd1 vccd1 vccd1 _12280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09428__B _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ _10449_/C _11231_/B _11231_/C _11231_/D vssd1 vssd1 vccd1 vccd1 _12110_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07229__A _08916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _10315_/X _11163_/C _11160_/X _11161_/Y vssd1 vssd1 vccd1 vccd1 _11164_/A
+ sky130_fd_sc_hd__o211a_2
XANTENNA__11194__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _11885_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10941__A1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12143__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _11094_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__nor2_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__and2_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold88/X vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ _11994_/A _11994_/B _12302_/A vssd1 vssd1 vccd1 vccd1 _11995_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08114__A2 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__A2 _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10946_ _10896_/A _10896_/B _10897_/Y vssd1 vssd1 vccd1 vccd1 _11010_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10877_ _10997_/B _10877_/B vssd1 vssd1 vccd1 vccd1 _10878_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _12616_/A _12620_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12029__B _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12547_ _12547_/A _12556_/A vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12478_ _12478_/A _12478_/B _12478_/C _12478_/D vssd1 vssd1 vccd1 vccd1 _12480_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA_3 curr_PC[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08523__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ _06652_/Y _11337_/X _06653_/A vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11185__B2 _11271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _07050_/A _06970_/B vssd1 vssd1 vccd1 vccd1 _06971_/B sky130_fd_sc_hd__nand2_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06697__B _07296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ _08640_/A _08657_/A _08640_/C vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__or3_1
XANTENNA__07561__B1 _07157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ _08814_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08605_/A sky130_fd_sc_hd__xnor2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07533_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10448__B1 _10681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07453_ _09420_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07458_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09066__A0 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__A _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07384_ _12712_/A _09727_/A _08798_/B _12714_/A vssd1 vssd1 vccd1 vccd1 _07385_/B
+ sky130_fd_sc_hd__o22a_1
X_09123_ reg1_val[6] reg1_val[25] _09124_/S vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08813__B1 _08813_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10963__A _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10591__A2_N _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _08044_/Y _08988_/B _08043_/A vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08005_ _08741_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11794__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ curr_PC[4] _09957_/C curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__a21oi_1
X_08907_ fanout74/X _10481_/A _07000_/A fanout68/X vssd1 vssd1 vccd1 vccd1 _08908_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09888_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__nand2b_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A1 _10481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__B2 _07000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10687__B1 _12179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _09002_/A _09002_/B _08650_/X vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10151__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _09222_/B2 _09568_/A _09428_/A _09422_/A vssd1 vssd1 vccd1 vccd1 _08770_/B
+ sky130_fd_sc_hd__o22a_1
X_11780_ _11781_/B _11854_/B hold191/A vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12979__A2 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _11232_/A _10800_/B _10800_/C vssd1 vssd1 vccd1 vccd1 _10800_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__07512__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ _11470_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10733_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _12410_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12403_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ _10539_/A _10538_/B _10538_/A vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ _11135_/S _09939_/X _09168_/A vssd1 vssd1 vccd1 vccd1 _11696_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12332_ _12333_/A _12333_/B _12333_/C vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _06821_/X _12262_/X _12263_/S vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _11214_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__xnor2_1
X_12194_ _09152_/Y _12189_/X _12190_/Y _12193_/X vssd1 vssd1 vccd1 vccd1 _12195_/D
+ sky130_fd_sc_hd__a31o_1
X_11145_ _06936_/A _06905_/Y _11142_/X _11144_/Y vssd1 vssd1 vccd1 vccd1 _11145_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09780__A1 _10320_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__A1 _12248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11212_/B _11087_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__and2_1
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10113__A _11885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__and2_1
X_10929_ hold216/A _11620_/B _11040_/B _10928_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1
+ _10929_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07422__A _11183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07846__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07846__B2 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06980__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09810_ _09810_/A _09810_/B _09810_/C vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__or3_1
Xfanout307 instruction[7] vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06953_ reg1_val[14] _06953_/B vssd1 vssd1 vccd1 vccd1 _06961_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10381__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ fanout80/X _11564_/A fanout38/X _10099_/A1 vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08700__B _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A2 fanout93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ instruction[20] _06850_/Y _06883_/X _06637_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _09610_/A _09610_/B _09608_/X vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__a21o_1
X_08623_ _08623_/A _08623_/B vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__and2_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09287__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08554_ _08842_/A _08843_/B _08843_/A vssd1 vssd1 vccd1 vccd1 _08555_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07505_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07505_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08485_ _08274_/A _10876_/A1 _08813_/A1 fanout93/X vssd1 vssd1 vccd1 vccd1 _08486_/B
+ sky130_fd_sc_hd__o22a_1
X_07436_ _07434_/A _07434_/B _07435_/X vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07367_ _07368_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09104_/X _09105_/X _09313_/S vssd1 vssd1 vccd1 vccd1 _09106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09039_/C sky130_fd_sc_hd__xnor2_2
X_07298_ reg1_val[18] _07298_/B vssd1 vssd1 vccd1 vccd1 _07301_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08014__B2 _08565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__A _12571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _06985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _09938_/Y _09471_/A _11134_/S vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__mux2_1
X_12950_ _11955_/A _12962_/B2 hold109/X vssd1 vssd1 vccd1 vccd1 _13216_/D sky130_fd_sc_hd__o21a_1
X_12881_ hold191/X _13070_/B2 _13070_/A2 hold220/X vssd1 vssd1 vccd1 vccd1 hold221/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _11902_/A _11902_/B _11902_/C vssd1 vssd1 vccd1 vccd1 _11973_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09722__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ _11869_/A _11759_/B _11871_/A vssd1 vssd1 vccd1 vccd1 _11833_/B sky130_fd_sc_hd__a21oi_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11763_ _11838_/A _09052_/C _09052_/B vssd1 vssd1 vccd1 vccd1 _11763_/X sky130_fd_sc_hd__a21o_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11617_/A _11617_/B _11615_/B vssd1 vssd1 vccd1 vccd1 _11695_/B sky130_fd_sc_hd__o21a_1
X_10714_ _09330_/A _10700_/X _10713_/Y _09120_/S _10712_/X vssd1 vssd1 vccd1 vccd1
+ _10715_/C sky130_fd_sc_hd__o221a_1
XFILLER_0_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10645_ _10876_/A1 fanout7/X fanout93/X fanout5/X vssd1 vssd1 vccd1 vccd1 _10646_/B
+ sky130_fd_sc_hd__o22a_1
X_12315_ _09498_/A _12297_/Y _12314_/X vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__o21ai_1
X_10576_ _10577_/A _10577_/B _10577_/C vssd1 vssd1 vccd1 vccd1 _10576_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _07268_/A fanout4/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08801__A _08801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _09053_/Y _09055_/Y _09621_/A vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07417__A _09979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12323__A _12502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _06831_/A _11126_/X _11127_/Y vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11059_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11063_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07152__A _07916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _09313_/S fanout43/X _08333_/B _09237_/A vssd1 vssd1 vccd1 vccd1 _08271_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07221_ _08698_/A _07221_/B vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07152_ _07916_/A _07152_/B vssd1 vssd1 vccd1 vccd1 _07152_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07083_ _07415_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07339_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10018__A _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A1 _07157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout104 _07127_/Y vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__buf_8
Xfanout115 _06999_/Y vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__buf_8
Xfanout126 _12694_/A vssd1 vssd1 vccd1 vccd1 _10377_/A1 sky130_fd_sc_hd__buf_4
Xfanout137 _09979_/A vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08430__B _08430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout148 _09698_/A vssd1 vssd1 vccd1 vccd1 _08733_/B1 sky130_fd_sc_hd__buf_6
X_07985_ _07985_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _07987_/B sky130_fd_sc_hd__xnor2_1
Xfanout159 _06915_/Y vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__clkbuf_16
X_06936_ _06936_/A _06963_/B _06936_/C vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__or3_4
XANTENNA__10106__A2 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _09724_/A _09724_/B vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__xor2_1
X_06867_ instruction[14] _06868_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
X_09655_ _09634_/A _09119_/X _09164_/B vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09542__A _10607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06885__B _06887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08606_ _08755_/A _08606_/A2 _08642_/B _08782_/B2 vssd1 vssd1 vccd1 vccd1 _08607_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07062__A _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06798_ _06798_/A _06798_/B vssd1 vssd1 vccd1 vccd1 _06798_/X sky130_fd_sc_hd__and2_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _11654_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11067__B1 _08233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ _08549_/B _08549_/A vssd1 vssd1 vccd1 vccd1 _08537_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08468_ _08465_/A _08466_/Y _08467_/Y _08427_/X vssd1 vssd1 vccd1 vccd1 _08510_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08483__A1 _08782_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08483__B2 _08756_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07419_ _07875_/A _07419_/B vssd1 vssd1 vccd1 vccd1 _07420_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _08699_/A2 _08715_/A2 _08735_/B1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 _08400_/B
+ sky130_fd_sc_hd__o22a_1
X_10430_ _10271_/A _10271_/B _10269_/X vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08235__A1 _11068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ fanout76/X fanout41/X _08135_/B _11663_/A vssd1 vssd1 vccd1 vccd1 _10362_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13080_ _13080_/A hold272/X vssd1 vssd1 vccd1 vccd1 _13247_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _12157_/A _12100_/B vssd1 vssd1 vccd1 vccd1 _12102_/C sky130_fd_sc_hd__nor2_1
XANTENNA__07994__B1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ _10172_/A _10172_/B _10170_/X vssd1 vssd1 vccd1 vccd1 _10300_/A sky130_fd_sc_hd__a21bo_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ _12032_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__nand2_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A1 _10450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10750__C1 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ hold83/X _12665_/A _12955_/B1 hold39/X _12970_/A vssd1 vssd1 vccd1 vccd1
+ hold84/A sky130_fd_sc_hd__o221a_1
XANTENNA__08171__B1 _08333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12864_ _13062_/A hold206/X vssd1 vssd1 vccd1 vccd1 _13173_/D sky130_fd_sc_hd__and2_1
XANTENNA__08068__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ _12976_/B _12977_/A _12785_/X vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__a21o_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11815_ _11816_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__nor2_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11746_ _11747_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__nand2_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12318__A _12499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ _11677_/A _11677_/B _11677_/C vssd1 vssd1 vccd1 vccd1 _11678_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10628_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ _10445_/A _10442_/X _10444_/B vssd1 vssd1 vccd1 vccd1 _10792_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11876__B _12095_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ _12271_/S _09474_/X _12228_/Y _09156_/B vssd1 vssd1 vccd1 vccd1 _12240_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08531__A _08607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07770_ _10850_/A _07770_/B vssd1 vssd1 vccd1 vccd1 _07771_/C sky130_fd_sc_hd__xnor2_1
X_06721_ _06753_/B _06646_/A _12532_/B _06720_/X vssd1 vssd1 vccd1 vccd1 _07158_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09440_ _09438_/Y _09440_/B vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08701__A2 _08730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06652_ _06653_/B vssd1 vssd1 vccd1 vccd1 _06652_/Y sky130_fd_sc_hd__inv_2
X_06583_ reg2_val[29] _06748_/B _06657_/B1 _06581_/X vssd1 vssd1 vccd1 vccd1 _06585_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09662__B1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__S _09309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08203_/A _08203_/B _08201_/X vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__a21oi_2
X_07204_ _07205_/B _07204_/B vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__and2b_1
XANTENNA_fanout132_A _12686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08217__B2 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08184_ _08128_/A _08128_/B _08129_/X vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07135_ _07138_/A _11727_/A _11796_/A vssd1 vssd1 vccd1 vccd1 _07135_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09965__B2 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A1 _10359_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ _07303_/A _07068_/A _06592_/B vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07440__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__A1 _11297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09717__B2 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__A _13085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07057__A _08798_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07976_/A _07976_/B _07958_/Y vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__a21o_1
X_06919_ reg1_val[12] _06919_/B vssd1 vssd1 vccd1 vccd1 _06922_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__06951__A1 _10920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _08700_/C _10845_/A _10845_/B _07044_/Y _10251_/A vssd1 vssd1 vccd1 vccd1
+ _09708_/B sky130_fd_sc_hd__a32o_1
X_07899_ _07899_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ _09493_/A _09490_/Y _09492_/B vssd1 vssd1 vccd1 vccd1 _09638_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout45_A _07391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _09424_/A _09424_/B _09420_/Y vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__a21oi_2
X_11600_ _11600_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__and3_1
X_12580_ reg1_val[16] _12615_/B vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ hold168/A _11620_/B _11619_/B _11530_/Y _11448_/A vssd1 vssd1 vccd1 vccd1
+ _11531_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09653__B1 _12265_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12004__A2 _09141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08208__B2 _08642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08208__A1 _08606_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _11462_/A _12245_/B _11462_/C vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__nor3_1
X_13201_ _13222_/CLK _13201_/D vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11393_ _11393_/A _11393_/B vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__or2_1
XANTENNA__10015__A1 _12141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10015__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _11184_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__xnor2_1
X_13132_ _13251_/CLK _13132_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ _06712_/B _09141_/Y _09137_/Y vssd1 vssd1 vccd1 vccd1 _10344_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13063_ _12749_/X _13063_/B vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11515__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10275_ _10275_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__nand2_1
X_12014_ _11951_/A _11951_/B _11949_/A vssd1 vssd1 vccd1 vccd1 _12026_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12916_ _06975_/B _12686_/B hold120/X vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10121__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ hold222/A _12885_/A2 _12885_/B1 hold213/X vssd1 vssd1 vccd1 vccd1 hold214/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08447__A1 _08670_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12778_ hold285/X hold68/X vssd1 vssd1 vccd1 vccd1 _12989_/B sky130_fd_sc_hd__nand2b_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__A2 _06905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08447__B2 _08699_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__A _08734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11729_ _11730_/A _11730_/B vssd1 vssd1 vccd1 vccd1 _11803_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11887__A _11887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08940_/Y sky130_fd_sc_hd__nand2_1
X_08871_ _09048_/A _09048_/B _09048_/C _08870_/Y vssd1 vssd1 vccd1 vccd1 _08871_/Y
+ sky130_fd_sc_hd__a31oi_2
X_07822_ _07823_/A _07823_/B _07823_/C vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06933__A1 _06960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _07753_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ reg1_val[9] _06931_/B vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07684_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07695_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06635_ reg1_val[19] _06980_/A vssd1 vssd1 vccd1 vccd1 _06636_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _09282_/A _09282_/B _09280_/X vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06566_ _06566_/A _12005_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__and2_1
XFILLER_0_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _08323_/A _08323_/B _08294_/X vssd1 vssd1 vccd1 vccd1 _08312_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08436__A _08814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__B2 _08219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__A1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09285_ _09461_/B _09285_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08236_ _08268_/A _08234_/X _08229_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08246_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__or2_2
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ reg1_val[23] _07284_/B _07118_/C vssd1 vssd1 vccd1 vccd1 _07149_/B sky130_fd_sc_hd__or3_2
XFILLER_0_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08610__B2 _08274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _07029_/B _07047_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07049_/X sky130_fd_sc_hd__a21o_1
X_10060_ instruction[7] _06730_/Y _06770_/Y _10059_/Y vssd1 vssd1 vccd1 vccd1 _10060_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12421__A _12576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A1 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ fanout60/X fanout37/X _08233_/B _12148_/A vssd1 vssd1 vccd1 vccd1 _10963_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07234__B _11184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _06946_/X _12731_/A2 hold67/X _13085_/A vssd1 vssd1 vccd1 vccd1 _13143_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10893_ _10894_/A _10894_/B _10894_/C vssd1 vssd1 vccd1 vccd1 _11003_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08346__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ _12640_/A _12632_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12563_ _12568_/B _12563_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _12491_/B _12493_/B _12491_/A vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _12223_/A _11514_/B _11514_/C vssd1 vssd1 vccd1 vccd1 _11514_/Y sky130_fd_sc_hd__nand3_1
X_11445_ hold179/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _11654_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11378_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ hold164/X hold100/X _13121_/A _13114_/X vssd1 vssd1 vccd1 vccd1 hold165/A
+ sky130_fd_sc_hd__o211a_1
X_10327_ _10327_/A _10327_/B vssd1 vssd1 vccd1 vccd1 _10327_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ hold253/X _13045_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13046_/X sky130_fd_sc_hd__mux2_1
X_10258_ _10377_/A1 fanout14/X fanout52/X _10490_/B2 vssd1 vssd1 vccd1 vccd1 _10259_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07168__B2 _09725_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07168__A1 _12710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _06723_/Y _10059_/B _06725_/B vssd1 vssd1 vccd1 vccd1 _10189_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10711__A2 _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13110__B1 _06858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07160__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ reg1_val[2] reg1_val[29] _09092_/S vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06851__B1 _06847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08021_ _08021_/A _08157_/A vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13101__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout6 fanout6/A vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__buf_8
XFILLER_0_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09972_/A _09972_/B vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08923_ _08924_/A _08924_/B vssd1 vssd1 vccd1 vccd1 _09194_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout297_A fanout298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A1 _07147_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__B2 _07157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ _07965_/A _07965_/C _07965_/B vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__a21oi_1
X_07805_ _07828_/B _07828_/A vssd1 vssd1 vccd1 vccd1 _07805_/Y sky130_fd_sc_hd__nand2b_1
X_08785_ _09422_/A _09237_/A _08813_/B1 _09222_/B2 vssd1 vssd1 vccd1 vccd1 _08786_/B
+ sky130_fd_sc_hd__o22a_1
X_07736_ _07738_/A _07736_/B vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06618_ reg1_val[21] _06987_/A vssd1 vssd1 vccd1 vccd1 _06619_/B sky130_fd_sc_hd__nor2_1
X_07598_ _09423_/A _07598_/B vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09406_ _09406_/A _09406_/B vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__xnor2_2
X_06549_ reg2_val[26] _06754_/B _06539_/X _06548_/X vssd1 vssd1 vccd1 vccd1 _07064_/A
+ sky130_fd_sc_hd__a22o_2
X_09337_ _09495_/C _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07070__A _10845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _09268_/A _09268_/B vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ _10957_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__or2_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09199_ _09200_/B _09200_/A vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ _11230_/A _11230_/B _11230_/C _11230_/D vssd1 vssd1 vccd1 vccd1 _11231_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _10677_/B _10792_/X _10793_/X _11157_/B vssd1 vssd1 vccd1 vccd1 _11161_/Y
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__11194__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ fanout8/X _10370_/A fanout6/X _12684_/A vssd1 vssd1 vccd1 vccd1 _10113_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12143__A1 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12143__B2 _12201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__xnor2_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ _10043_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__xnor2_2
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07245__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ _11994_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _10899_/A _10899_/B _10901_/Y vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876_ _10876_/A1 _11296_/A _10875_/C vssd1 vssd1 vccd1 vccd1 _10877_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12615_ reg1_val[23] _12615_/B vssd1 vssd1 vccd1 vccd1 _12620_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08822__B2 _12499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ reg1_val[10] _12546_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ _12484_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 curr_PC[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11230__A _11230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _11339_/Y _11340_/X _11347_/X _11358_/X vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06978__B _06978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _12761_/X _13029_/B vssd1 vssd1 vccd1 vccd1 _13030_/B sky130_fd_sc_hd__nand2b_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07561__B2 _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08570_ _08813_/A1 _10506_/A _10647_/A _08274_/A vssd1 vssd1 vccd1 vccd1 _08571_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07521_ _07521_/A _07521_/B vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07452_ _06828_/A _12720_/A _12718_/A _08765_/A vssd1 vssd1 vccd1 vccd1 _07453_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _09420_/A _07383_/B vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _09120_/X _09121_/X _09319_/S vssd1 vssd1 vccd1 vccd1 _09122_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07077__B1 _08276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12070__B1 _12309_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__A1 _08813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__B2 _06828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A _08714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _09056_/B _09056_/C vssd1 vssd1 vccd1 vccd1 _09053_/Y sky130_fd_sc_hd__nor2_1
X_08004_ _10957_/A _08740_/A2 _08755_/B fanout81/X vssd1 vssd1 vccd1 vccd1 _08005_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_114_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__B1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _09061_/X _09918_/Y _09919_/X _09922_/X _09954_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/X sky130_fd_sc_hd__o311a_2
XANTENNA__13067__A _13071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _10252_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__xnor2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10136__B1 _07799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _09886_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11884__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ _09003_/A _09003_/B _08679_/X vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__a21o_1
X_08768_ _09420_/A _08768_/B _08768_/C vssd1 vssd1 vccd1 vccd1 _08771_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07719_ _07830_/A _07830_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07722_/B sky130_fd_sc_hd__a21o_1
X_08699_ _08755_/A _08699_/A2 _10398_/A vssd1 vssd1 vccd1 vccd1 _08730_/B sky130_fd_sc_hd__o21a_1
XANTENNA__13006__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ fanout64/X fanout41/X _08135_/B _11876_/A vssd1 vssd1 vccd1 vccd1 _10731_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _10540_/A _10540_/B _10523_/A vssd1 vssd1 vccd1 vccd1 _10671_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _12559_/B _12400_/B vssd1 vssd1 vccd1 vccd1 _12401_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ _10584_/Y _10585_/X _10587_/Y _10591_/X vssd1 vssd1 vccd1 vccd1 _10592_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12331_ _12340_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _12333_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12262_ _06586_/B _12219_/X _06584_/X vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_121_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10083__A2_N _12238_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _11213_/A _11213_/B vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__nor2_1
X_12193_ _09064_/Y _09637_/X _09658_/Y _09135_/Y _12192_/X vssd1 vssd1 vccd1 vccd1
+ _12193_/X sky130_fd_sc_hd__a221o_1
X_11144_ _12309_/B1 _11143_/X _06669_/B vssd1 vssd1 vccd1 vccd1 _11144_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07240__B1 _07239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10127__B1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11075_ _11075_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11087_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12667__A2 _12926_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08740__B1 _08755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _11976_/A _11976_/B _11976_/C vssd1 vssd1 vccd1 vccd1 _11978_/B sky130_fd_sc_hd__a21o_1
X_10928_ _11620_/B _11040_/B hold216/A vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07846__A2 _07040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ _11656_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _12529_/A _12529_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 instruction[2] vssd1 vssd1 vccd1 vccd1 _06850_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__07231__B1 _07050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09365__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__A_N _09464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06952_ reg1_val[15] _06952_/B vssd1 vssd1 vccd1 vccd1 _06952_/X sky130_fd_sc_hd__xor2_1
X_09740_ _11796_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__xnor2_1
.ends

