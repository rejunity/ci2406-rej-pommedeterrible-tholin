VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO icache
  CLASS BLOCK ;
  FOREIGN icache ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 850.000 ;
  PIN cache_entry[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END cache_entry[0]
  PIN cache_entry[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END cache_entry[100]
  PIN cache_entry[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END cache_entry[101]
  PIN cache_entry[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END cache_entry[102]
  PIN cache_entry[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END cache_entry[103]
  PIN cache_entry[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END cache_entry[104]
  PIN cache_entry[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END cache_entry[105]
  PIN cache_entry[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END cache_entry[106]
  PIN cache_entry[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END cache_entry[107]
  PIN cache_entry[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END cache_entry[108]
  PIN cache_entry[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END cache_entry[109]
  PIN cache_entry[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END cache_entry[10]
  PIN cache_entry[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END cache_entry[110]
  PIN cache_entry[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END cache_entry[111]
  PIN cache_entry[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END cache_entry[112]
  PIN cache_entry[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END cache_entry[113]
  PIN cache_entry[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END cache_entry[114]
  PIN cache_entry[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END cache_entry[115]
  PIN cache_entry[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END cache_entry[116]
  PIN cache_entry[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END cache_entry[117]
  PIN cache_entry[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END cache_entry[118]
  PIN cache_entry[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END cache_entry[119]
  PIN cache_entry[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END cache_entry[11]
  PIN cache_entry[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END cache_entry[120]
  PIN cache_entry[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END cache_entry[121]
  PIN cache_entry[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END cache_entry[122]
  PIN cache_entry[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END cache_entry[123]
  PIN cache_entry[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END cache_entry[124]
  PIN cache_entry[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END cache_entry[125]
  PIN cache_entry[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END cache_entry[126]
  PIN cache_entry[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END cache_entry[127]
  PIN cache_entry[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END cache_entry[12]
  PIN cache_entry[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cache_entry[13]
  PIN cache_entry[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END cache_entry[14]
  PIN cache_entry[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END cache_entry[15]
  PIN cache_entry[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cache_entry[16]
  PIN cache_entry[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END cache_entry[17]
  PIN cache_entry[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END cache_entry[18]
  PIN cache_entry[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END cache_entry[19]
  PIN cache_entry[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END cache_entry[1]
  PIN cache_entry[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END cache_entry[20]
  PIN cache_entry[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END cache_entry[21]
  PIN cache_entry[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END cache_entry[22]
  PIN cache_entry[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END cache_entry[23]
  PIN cache_entry[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END cache_entry[24]
  PIN cache_entry[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END cache_entry[25]
  PIN cache_entry[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END cache_entry[26]
  PIN cache_entry[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END cache_entry[27]
  PIN cache_entry[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END cache_entry[28]
  PIN cache_entry[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END cache_entry[29]
  PIN cache_entry[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END cache_entry[2]
  PIN cache_entry[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END cache_entry[30]
  PIN cache_entry[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END cache_entry[31]
  PIN cache_entry[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END cache_entry[32]
  PIN cache_entry[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END cache_entry[33]
  PIN cache_entry[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END cache_entry[34]
  PIN cache_entry[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END cache_entry[35]
  PIN cache_entry[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END cache_entry[36]
  PIN cache_entry[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END cache_entry[37]
  PIN cache_entry[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END cache_entry[38]
  PIN cache_entry[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END cache_entry[39]
  PIN cache_entry[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END cache_entry[3]
  PIN cache_entry[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END cache_entry[40]
  PIN cache_entry[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END cache_entry[41]
  PIN cache_entry[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END cache_entry[42]
  PIN cache_entry[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END cache_entry[43]
  PIN cache_entry[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END cache_entry[44]
  PIN cache_entry[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END cache_entry[45]
  PIN cache_entry[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END cache_entry[46]
  PIN cache_entry[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END cache_entry[47]
  PIN cache_entry[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END cache_entry[48]
  PIN cache_entry[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END cache_entry[49]
  PIN cache_entry[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END cache_entry[4]
  PIN cache_entry[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END cache_entry[50]
  PIN cache_entry[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END cache_entry[51]
  PIN cache_entry[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END cache_entry[52]
  PIN cache_entry[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END cache_entry[53]
  PIN cache_entry[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END cache_entry[54]
  PIN cache_entry[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END cache_entry[55]
  PIN cache_entry[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END cache_entry[56]
  PIN cache_entry[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END cache_entry[57]
  PIN cache_entry[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END cache_entry[58]
  PIN cache_entry[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END cache_entry[59]
  PIN cache_entry[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END cache_entry[5]
  PIN cache_entry[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END cache_entry[60]
  PIN cache_entry[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END cache_entry[61]
  PIN cache_entry[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END cache_entry[62]
  PIN cache_entry[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END cache_entry[63]
  PIN cache_entry[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END cache_entry[64]
  PIN cache_entry[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END cache_entry[65]
  PIN cache_entry[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END cache_entry[66]
  PIN cache_entry[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END cache_entry[67]
  PIN cache_entry[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END cache_entry[68]
  PIN cache_entry[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END cache_entry[69]
  PIN cache_entry[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END cache_entry[6]
  PIN cache_entry[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END cache_entry[70]
  PIN cache_entry[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END cache_entry[71]
  PIN cache_entry[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END cache_entry[72]
  PIN cache_entry[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END cache_entry[73]
  PIN cache_entry[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END cache_entry[74]
  PIN cache_entry[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END cache_entry[75]
  PIN cache_entry[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END cache_entry[76]
  PIN cache_entry[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END cache_entry[77]
  PIN cache_entry[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END cache_entry[78]
  PIN cache_entry[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END cache_entry[79]
  PIN cache_entry[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END cache_entry[7]
  PIN cache_entry[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END cache_entry[80]
  PIN cache_entry[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END cache_entry[81]
  PIN cache_entry[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END cache_entry[82]
  PIN cache_entry[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END cache_entry[83]
  PIN cache_entry[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END cache_entry[84]
  PIN cache_entry[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END cache_entry[85]
  PIN cache_entry[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END cache_entry[86]
  PIN cache_entry[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END cache_entry[87]
  PIN cache_entry[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END cache_entry[88]
  PIN cache_entry[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cache_entry[89]
  PIN cache_entry[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END cache_entry[8]
  PIN cache_entry[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END cache_entry[90]
  PIN cache_entry[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END cache_entry[91]
  PIN cache_entry[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END cache_entry[92]
  PIN cache_entry[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END cache_entry[93]
  PIN cache_entry[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END cache_entry[94]
  PIN cache_entry[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END cache_entry[95]
  PIN cache_entry[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END cache_entry[96]
  PIN cache_entry[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END cache_entry[97]
  PIN cache_entry[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END cache_entry[98]
  PIN cache_entry[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END cache_entry[99]
  PIN cache_entry[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END cache_entry[9]
  PIN cache_hit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 489.530 846.000 489.810 850.000 ;
    END
  END cache_hit
  PIN curr_PC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 20.440 700.000 21.040 ;
    END
  END curr_PC[0]
  PIN curr_PC[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 319.640 700.000 320.240 ;
    END
  END curr_PC[10]
  PIN curr_PC[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.099500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 696.000 349.560 700.000 350.160 ;
    END
  END curr_PC[11]
  PIN curr_PC[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 379.480 700.000 380.080 ;
    END
  END curr_PC[12]
  PIN curr_PC[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 409.400 700.000 410.000 ;
    END
  END curr_PC[13]
  PIN curr_PC[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 439.320 700.000 439.920 ;
    END
  END curr_PC[14]
  PIN curr_PC[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 469.240 700.000 469.840 ;
    END
  END curr_PC[15]
  PIN curr_PC[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 499.160 700.000 499.760 ;
    END
  END curr_PC[16]
  PIN curr_PC[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 529.080 700.000 529.680 ;
    END
  END curr_PC[17]
  PIN curr_PC[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 559.000 700.000 559.600 ;
    END
  END curr_PC[18]
  PIN curr_PC[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.970000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 588.920 700.000 589.520 ;
    END
  END curr_PC[19]
  PIN curr_PC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 696.000 50.360 700.000 50.960 ;
    END
  END curr_PC[1]
  PIN curr_PC[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 618.840 700.000 619.440 ;
    END
  END curr_PC[20]
  PIN curr_PC[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.207500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 648.760 700.000 649.360 ;
    END
  END curr_PC[21]
  PIN curr_PC[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 678.680 700.000 679.280 ;
    END
  END curr_PC[22]
  PIN curr_PC[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.217500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 708.600 700.000 709.200 ;
    END
  END curr_PC[23]
  PIN curr_PC[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.465000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 738.520 700.000 739.120 ;
    END
  END curr_PC[24]
  PIN curr_PC[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.712500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 768.440 700.000 769.040 ;
    END
  END curr_PC[25]
  PIN curr_PC[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 798.360 700.000 798.960 ;
    END
  END curr_PC[26]
  PIN curr_PC[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.320500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 828.280 700.000 828.880 ;
    END
  END curr_PC[27]
  PIN curr_PC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 80.280 700.000 80.880 ;
    END
  END curr_PC[2]
  PIN curr_PC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 110.200 700.000 110.800 ;
    END
  END curr_PC[3]
  PIN curr_PC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 140.120 700.000 140.720 ;
    END
  END curr_PC[4]
  PIN curr_PC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 696.000 170.040 700.000 170.640 ;
    END
  END curr_PC[5]
  PIN curr_PC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 696.000 199.960 700.000 200.560 ;
    END
  END curr_PC[6]
  PIN curr_PC[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 229.880 700.000 230.480 ;
    END
  END curr_PC[7]
  PIN curr_PC[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 259.800 700.000 260.400 ;
    END
  END curr_PC[8]
  PIN curr_PC[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 289.720 700.000 290.320 ;
    END
  END curr_PC[9]
  PIN entry_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    PORT
      LAYER met2 ;
        RECT 629.370 846.000 629.650 850.000 ;
    END
  END entry_valid
  PIN invalidate
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met2 ;
        RECT 349.690 846.000 349.970 850.000 ;
    END
  END invalidate
  PIN new_entry[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END new_entry[0]
  PIN new_entry[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END new_entry[100]
  PIN new_entry[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END new_entry[101]
  PIN new_entry[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END new_entry[102]
  PIN new_entry[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END new_entry[103]
  PIN new_entry[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END new_entry[104]
  PIN new_entry[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END new_entry[105]
  PIN new_entry[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END new_entry[106]
  PIN new_entry[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END new_entry[107]
  PIN new_entry[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END new_entry[108]
  PIN new_entry[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END new_entry[109]
  PIN new_entry[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END new_entry[10]
  PIN new_entry[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END new_entry[110]
  PIN new_entry[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END new_entry[111]
  PIN new_entry[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END new_entry[112]
  PIN new_entry[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END new_entry[113]
  PIN new_entry[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END new_entry[114]
  PIN new_entry[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END new_entry[115]
  PIN new_entry[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END new_entry[116]
  PIN new_entry[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END new_entry[117]
  PIN new_entry[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END new_entry[118]
  PIN new_entry[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END new_entry[119]
  PIN new_entry[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END new_entry[11]
  PIN new_entry[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END new_entry[120]
  PIN new_entry[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END new_entry[121]
  PIN new_entry[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END new_entry[122]
  PIN new_entry[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END new_entry[123]
  PIN new_entry[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END new_entry[124]
  PIN new_entry[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END new_entry[125]
  PIN new_entry[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END new_entry[126]
  PIN new_entry[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END new_entry[127]
  PIN new_entry[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END new_entry[12]
  PIN new_entry[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END new_entry[13]
  PIN new_entry[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END new_entry[14]
  PIN new_entry[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END new_entry[15]
  PIN new_entry[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END new_entry[16]
  PIN new_entry[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END new_entry[17]
  PIN new_entry[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END new_entry[18]
  PIN new_entry[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END new_entry[19]
  PIN new_entry[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END new_entry[1]
  PIN new_entry[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END new_entry[20]
  PIN new_entry[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END new_entry[21]
  PIN new_entry[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END new_entry[22]
  PIN new_entry[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END new_entry[23]
  PIN new_entry[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END new_entry[24]
  PIN new_entry[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END new_entry[25]
  PIN new_entry[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END new_entry[26]
  PIN new_entry[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END new_entry[27]
  PIN new_entry[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END new_entry[28]
  PIN new_entry[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END new_entry[29]
  PIN new_entry[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END new_entry[2]
  PIN new_entry[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END new_entry[30]
  PIN new_entry[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END new_entry[31]
  PIN new_entry[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END new_entry[32]
  PIN new_entry[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END new_entry[33]
  PIN new_entry[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END new_entry[34]
  PIN new_entry[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END new_entry[35]
  PIN new_entry[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END new_entry[36]
  PIN new_entry[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END new_entry[37]
  PIN new_entry[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END new_entry[38]
  PIN new_entry[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END new_entry[39]
  PIN new_entry[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END new_entry[3]
  PIN new_entry[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END new_entry[40]
  PIN new_entry[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END new_entry[41]
  PIN new_entry[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END new_entry[42]
  PIN new_entry[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END new_entry[43]
  PIN new_entry[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END new_entry[44]
  PIN new_entry[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END new_entry[45]
  PIN new_entry[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END new_entry[46]
  PIN new_entry[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END new_entry[47]
  PIN new_entry[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END new_entry[48]
  PIN new_entry[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END new_entry[49]
  PIN new_entry[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END new_entry[4]
  PIN new_entry[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END new_entry[50]
  PIN new_entry[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END new_entry[51]
  PIN new_entry[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END new_entry[52]
  PIN new_entry[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END new_entry[53]
  PIN new_entry[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END new_entry[54]
  PIN new_entry[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END new_entry[55]
  PIN new_entry[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END new_entry[56]
  PIN new_entry[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END new_entry[57]
  PIN new_entry[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END new_entry[58]
  PIN new_entry[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END new_entry[59]
  PIN new_entry[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END new_entry[5]
  PIN new_entry[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END new_entry[60]
  PIN new_entry[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END new_entry[61]
  PIN new_entry[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END new_entry[62]
  PIN new_entry[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END new_entry[63]
  PIN new_entry[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END new_entry[64]
  PIN new_entry[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END new_entry[65]
  PIN new_entry[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END new_entry[66]
  PIN new_entry[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END new_entry[67]
  PIN new_entry[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END new_entry[68]
  PIN new_entry[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END new_entry[69]
  PIN new_entry[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END new_entry[6]
  PIN new_entry[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END new_entry[70]
  PIN new_entry[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END new_entry[71]
  PIN new_entry[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END new_entry[72]
  PIN new_entry[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END new_entry[73]
  PIN new_entry[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END new_entry[74]
  PIN new_entry[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END new_entry[75]
  PIN new_entry[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END new_entry[76]
  PIN new_entry[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END new_entry[77]
  PIN new_entry[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END new_entry[78]
  PIN new_entry[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END new_entry[79]
  PIN new_entry[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END new_entry[7]
  PIN new_entry[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END new_entry[80]
  PIN new_entry[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 6.520500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END new_entry[81]
  PIN new_entry[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END new_entry[82]
  PIN new_entry[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END new_entry[83]
  PIN new_entry[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END new_entry[84]
  PIN new_entry[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END new_entry[85]
  PIN new_entry[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END new_entry[86]
  PIN new_entry[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END new_entry[87]
  PIN new_entry[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END new_entry[88]
  PIN new_entry[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END new_entry[89]
  PIN new_entry[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END new_entry[8]
  PIN new_entry[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END new_entry[90]
  PIN new_entry[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END new_entry[91]
  PIN new_entry[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END new_entry[92]
  PIN new_entry[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END new_entry[93]
  PIN new_entry[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END new_entry[94]
  PIN new_entry[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END new_entry[95]
  PIN new_entry[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END new_entry[96]
  PIN new_entry[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END new_entry[97]
  PIN new_entry[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END new_entry[98]
  PIN new_entry[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END new_entry[99]
  PIN new_entry[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END new_entry[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.853000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 846.000 210.130 850.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 838.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 838.000 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 846.000 70.290 850.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 837.845 ;
      LAYER met1 ;
        RECT 5.520 10.640 694.440 838.000 ;
      LAYER met2 ;
        RECT 7.000 845.720 69.730 846.000 ;
        RECT 70.570 845.720 209.570 846.000 ;
        RECT 210.410 845.720 349.410 846.000 ;
        RECT 350.250 845.720 489.250 846.000 ;
        RECT 490.090 845.720 629.090 846.000 ;
        RECT 629.930 845.720 693.120 846.000 ;
        RECT 7.000 4.280 693.120 845.720 ;
        RECT 7.000 3.670 28.330 4.280 ;
        RECT 29.170 3.670 33.390 4.280 ;
        RECT 34.230 3.670 38.450 4.280 ;
        RECT 39.290 3.670 43.510 4.280 ;
        RECT 44.350 3.670 48.570 4.280 ;
        RECT 49.410 3.670 53.630 4.280 ;
        RECT 54.470 3.670 58.690 4.280 ;
        RECT 59.530 3.670 63.750 4.280 ;
        RECT 64.590 3.670 68.810 4.280 ;
        RECT 69.650 3.670 73.870 4.280 ;
        RECT 74.710 3.670 78.930 4.280 ;
        RECT 79.770 3.670 83.990 4.280 ;
        RECT 84.830 3.670 89.050 4.280 ;
        RECT 89.890 3.670 94.110 4.280 ;
        RECT 94.950 3.670 99.170 4.280 ;
        RECT 100.010 3.670 104.230 4.280 ;
        RECT 105.070 3.670 109.290 4.280 ;
        RECT 110.130 3.670 114.350 4.280 ;
        RECT 115.190 3.670 119.410 4.280 ;
        RECT 120.250 3.670 124.470 4.280 ;
        RECT 125.310 3.670 129.530 4.280 ;
        RECT 130.370 3.670 134.590 4.280 ;
        RECT 135.430 3.670 139.650 4.280 ;
        RECT 140.490 3.670 144.710 4.280 ;
        RECT 145.550 3.670 149.770 4.280 ;
        RECT 150.610 3.670 154.830 4.280 ;
        RECT 155.670 3.670 159.890 4.280 ;
        RECT 160.730 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.010 4.280 ;
        RECT 170.850 3.670 175.070 4.280 ;
        RECT 175.910 3.670 180.130 4.280 ;
        RECT 180.970 3.670 185.190 4.280 ;
        RECT 186.030 3.670 190.250 4.280 ;
        RECT 191.090 3.670 195.310 4.280 ;
        RECT 196.150 3.670 200.370 4.280 ;
        RECT 201.210 3.670 205.430 4.280 ;
        RECT 206.270 3.670 210.490 4.280 ;
        RECT 211.330 3.670 215.550 4.280 ;
        RECT 216.390 3.670 220.610 4.280 ;
        RECT 221.450 3.670 225.670 4.280 ;
        RECT 226.510 3.670 230.730 4.280 ;
        RECT 231.570 3.670 235.790 4.280 ;
        RECT 236.630 3.670 240.850 4.280 ;
        RECT 241.690 3.670 245.910 4.280 ;
        RECT 246.750 3.670 250.970 4.280 ;
        RECT 251.810 3.670 256.030 4.280 ;
        RECT 256.870 3.670 261.090 4.280 ;
        RECT 261.930 3.670 266.150 4.280 ;
        RECT 266.990 3.670 271.210 4.280 ;
        RECT 272.050 3.670 276.270 4.280 ;
        RECT 277.110 3.670 281.330 4.280 ;
        RECT 282.170 3.670 286.390 4.280 ;
        RECT 287.230 3.670 291.450 4.280 ;
        RECT 292.290 3.670 296.510 4.280 ;
        RECT 297.350 3.670 301.570 4.280 ;
        RECT 302.410 3.670 306.630 4.280 ;
        RECT 307.470 3.670 311.690 4.280 ;
        RECT 312.530 3.670 316.750 4.280 ;
        RECT 317.590 3.670 321.810 4.280 ;
        RECT 322.650 3.670 326.870 4.280 ;
        RECT 327.710 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.990 4.280 ;
        RECT 337.830 3.670 342.050 4.280 ;
        RECT 342.890 3.670 347.110 4.280 ;
        RECT 347.950 3.670 352.170 4.280 ;
        RECT 353.010 3.670 357.230 4.280 ;
        RECT 358.070 3.670 362.290 4.280 ;
        RECT 363.130 3.670 367.350 4.280 ;
        RECT 368.190 3.670 372.410 4.280 ;
        RECT 373.250 3.670 377.470 4.280 ;
        RECT 378.310 3.670 382.530 4.280 ;
        RECT 383.370 3.670 387.590 4.280 ;
        RECT 388.430 3.670 392.650 4.280 ;
        RECT 393.490 3.670 397.710 4.280 ;
        RECT 398.550 3.670 402.770 4.280 ;
        RECT 403.610 3.670 407.830 4.280 ;
        RECT 408.670 3.670 412.890 4.280 ;
        RECT 413.730 3.670 417.950 4.280 ;
        RECT 418.790 3.670 423.010 4.280 ;
        RECT 423.850 3.670 428.070 4.280 ;
        RECT 428.910 3.670 433.130 4.280 ;
        RECT 433.970 3.670 438.190 4.280 ;
        RECT 439.030 3.670 443.250 4.280 ;
        RECT 444.090 3.670 448.310 4.280 ;
        RECT 449.150 3.670 453.370 4.280 ;
        RECT 454.210 3.670 458.430 4.280 ;
        RECT 459.270 3.670 463.490 4.280 ;
        RECT 464.330 3.670 468.550 4.280 ;
        RECT 469.390 3.670 473.610 4.280 ;
        RECT 474.450 3.670 478.670 4.280 ;
        RECT 479.510 3.670 483.730 4.280 ;
        RECT 484.570 3.670 488.790 4.280 ;
        RECT 489.630 3.670 493.850 4.280 ;
        RECT 494.690 3.670 498.910 4.280 ;
        RECT 499.750 3.670 503.970 4.280 ;
        RECT 504.810 3.670 509.030 4.280 ;
        RECT 509.870 3.670 514.090 4.280 ;
        RECT 514.930 3.670 519.150 4.280 ;
        RECT 519.990 3.670 524.210 4.280 ;
        RECT 525.050 3.670 529.270 4.280 ;
        RECT 530.110 3.670 534.330 4.280 ;
        RECT 535.170 3.670 539.390 4.280 ;
        RECT 540.230 3.670 544.450 4.280 ;
        RECT 545.290 3.670 549.510 4.280 ;
        RECT 550.350 3.670 554.570 4.280 ;
        RECT 555.410 3.670 559.630 4.280 ;
        RECT 560.470 3.670 564.690 4.280 ;
        RECT 565.530 3.670 569.750 4.280 ;
        RECT 570.590 3.670 574.810 4.280 ;
        RECT 575.650 3.670 579.870 4.280 ;
        RECT 580.710 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.990 4.280 ;
        RECT 590.830 3.670 595.050 4.280 ;
        RECT 595.890 3.670 600.110 4.280 ;
        RECT 600.950 3.670 605.170 4.280 ;
        RECT 606.010 3.670 610.230 4.280 ;
        RECT 611.070 3.670 615.290 4.280 ;
        RECT 616.130 3.670 620.350 4.280 ;
        RECT 621.190 3.670 625.410 4.280 ;
        RECT 626.250 3.670 630.470 4.280 ;
        RECT 631.310 3.670 635.530 4.280 ;
        RECT 636.370 3.670 640.590 4.280 ;
        RECT 641.430 3.670 645.650 4.280 ;
        RECT 646.490 3.670 650.710 4.280 ;
        RECT 651.550 3.670 655.770 4.280 ;
        RECT 656.610 3.670 660.830 4.280 ;
        RECT 661.670 3.670 665.890 4.280 ;
        RECT 666.730 3.670 670.950 4.280 ;
        RECT 671.790 3.670 693.120 4.280 ;
      LAYER met3 ;
        RECT 3.070 829.280 696.000 837.925 ;
        RECT 3.070 827.880 695.600 829.280 ;
        RECT 3.070 799.360 696.000 827.880 ;
        RECT 3.070 797.960 695.600 799.360 ;
        RECT 3.070 770.800 696.000 797.960 ;
        RECT 4.400 769.440 696.000 770.800 ;
        RECT 4.400 769.400 695.600 769.440 ;
        RECT 3.070 768.040 695.600 769.400 ;
        RECT 3.070 765.360 696.000 768.040 ;
        RECT 4.400 763.960 696.000 765.360 ;
        RECT 3.070 759.920 696.000 763.960 ;
        RECT 4.400 758.520 696.000 759.920 ;
        RECT 3.070 754.480 696.000 758.520 ;
        RECT 4.400 753.080 696.000 754.480 ;
        RECT 3.070 749.040 696.000 753.080 ;
        RECT 4.400 747.640 696.000 749.040 ;
        RECT 3.070 743.600 696.000 747.640 ;
        RECT 4.400 742.200 696.000 743.600 ;
        RECT 3.070 739.520 696.000 742.200 ;
        RECT 3.070 738.160 695.600 739.520 ;
        RECT 4.400 738.120 695.600 738.160 ;
        RECT 4.400 736.760 696.000 738.120 ;
        RECT 3.070 732.720 696.000 736.760 ;
        RECT 4.400 731.320 696.000 732.720 ;
        RECT 3.070 727.280 696.000 731.320 ;
        RECT 4.400 725.880 696.000 727.280 ;
        RECT 3.070 721.840 696.000 725.880 ;
        RECT 4.400 720.440 696.000 721.840 ;
        RECT 3.070 716.400 696.000 720.440 ;
        RECT 4.400 715.000 696.000 716.400 ;
        RECT 3.070 710.960 696.000 715.000 ;
        RECT 4.400 709.600 696.000 710.960 ;
        RECT 4.400 709.560 695.600 709.600 ;
        RECT 3.070 708.200 695.600 709.560 ;
        RECT 3.070 705.520 696.000 708.200 ;
        RECT 4.400 704.120 696.000 705.520 ;
        RECT 3.070 700.080 696.000 704.120 ;
        RECT 4.400 698.680 696.000 700.080 ;
        RECT 3.070 694.640 696.000 698.680 ;
        RECT 4.400 693.240 696.000 694.640 ;
        RECT 3.070 689.200 696.000 693.240 ;
        RECT 4.400 687.800 696.000 689.200 ;
        RECT 3.070 683.760 696.000 687.800 ;
        RECT 4.400 682.360 696.000 683.760 ;
        RECT 3.070 679.680 696.000 682.360 ;
        RECT 3.070 678.320 695.600 679.680 ;
        RECT 4.400 678.280 695.600 678.320 ;
        RECT 4.400 676.920 696.000 678.280 ;
        RECT 3.070 672.880 696.000 676.920 ;
        RECT 4.400 671.480 696.000 672.880 ;
        RECT 3.070 667.440 696.000 671.480 ;
        RECT 4.400 666.040 696.000 667.440 ;
        RECT 3.070 662.000 696.000 666.040 ;
        RECT 4.400 660.600 696.000 662.000 ;
        RECT 3.070 656.560 696.000 660.600 ;
        RECT 4.400 655.160 696.000 656.560 ;
        RECT 3.070 651.120 696.000 655.160 ;
        RECT 4.400 649.760 696.000 651.120 ;
        RECT 4.400 649.720 695.600 649.760 ;
        RECT 3.070 648.360 695.600 649.720 ;
        RECT 3.070 645.680 696.000 648.360 ;
        RECT 4.400 644.280 696.000 645.680 ;
        RECT 3.070 640.240 696.000 644.280 ;
        RECT 4.400 638.840 696.000 640.240 ;
        RECT 3.070 634.800 696.000 638.840 ;
        RECT 4.400 633.400 696.000 634.800 ;
        RECT 3.070 629.360 696.000 633.400 ;
        RECT 4.400 627.960 696.000 629.360 ;
        RECT 3.070 623.920 696.000 627.960 ;
        RECT 4.400 622.520 696.000 623.920 ;
        RECT 3.070 619.840 696.000 622.520 ;
        RECT 3.070 618.480 695.600 619.840 ;
        RECT 4.400 618.440 695.600 618.480 ;
        RECT 4.400 617.080 696.000 618.440 ;
        RECT 3.070 613.040 696.000 617.080 ;
        RECT 4.400 611.640 696.000 613.040 ;
        RECT 3.070 607.600 696.000 611.640 ;
        RECT 4.400 606.200 696.000 607.600 ;
        RECT 3.070 602.160 696.000 606.200 ;
        RECT 4.400 600.760 696.000 602.160 ;
        RECT 3.070 596.720 696.000 600.760 ;
        RECT 4.400 595.320 696.000 596.720 ;
        RECT 3.070 591.280 696.000 595.320 ;
        RECT 4.400 589.920 696.000 591.280 ;
        RECT 4.400 589.880 695.600 589.920 ;
        RECT 3.070 588.520 695.600 589.880 ;
        RECT 3.070 585.840 696.000 588.520 ;
        RECT 4.400 584.440 696.000 585.840 ;
        RECT 3.070 580.400 696.000 584.440 ;
        RECT 4.400 579.000 696.000 580.400 ;
        RECT 3.070 574.960 696.000 579.000 ;
        RECT 4.400 573.560 696.000 574.960 ;
        RECT 3.070 569.520 696.000 573.560 ;
        RECT 4.400 568.120 696.000 569.520 ;
        RECT 3.070 564.080 696.000 568.120 ;
        RECT 4.400 562.680 696.000 564.080 ;
        RECT 3.070 560.000 696.000 562.680 ;
        RECT 3.070 558.640 695.600 560.000 ;
        RECT 4.400 558.600 695.600 558.640 ;
        RECT 4.400 557.240 696.000 558.600 ;
        RECT 3.070 553.200 696.000 557.240 ;
        RECT 4.400 551.800 696.000 553.200 ;
        RECT 3.070 547.760 696.000 551.800 ;
        RECT 4.400 546.360 696.000 547.760 ;
        RECT 3.070 542.320 696.000 546.360 ;
        RECT 4.400 540.920 696.000 542.320 ;
        RECT 3.070 536.880 696.000 540.920 ;
        RECT 4.400 535.480 696.000 536.880 ;
        RECT 3.070 531.440 696.000 535.480 ;
        RECT 4.400 530.080 696.000 531.440 ;
        RECT 4.400 530.040 695.600 530.080 ;
        RECT 3.070 528.680 695.600 530.040 ;
        RECT 3.070 526.000 696.000 528.680 ;
        RECT 4.400 524.600 696.000 526.000 ;
        RECT 3.070 520.560 696.000 524.600 ;
        RECT 4.400 519.160 696.000 520.560 ;
        RECT 3.070 515.120 696.000 519.160 ;
        RECT 4.400 513.720 696.000 515.120 ;
        RECT 3.070 509.680 696.000 513.720 ;
        RECT 4.400 508.280 696.000 509.680 ;
        RECT 3.070 504.240 696.000 508.280 ;
        RECT 4.400 502.840 696.000 504.240 ;
        RECT 3.070 500.160 696.000 502.840 ;
        RECT 3.070 498.800 695.600 500.160 ;
        RECT 4.400 498.760 695.600 498.800 ;
        RECT 4.400 497.400 696.000 498.760 ;
        RECT 3.070 493.360 696.000 497.400 ;
        RECT 4.400 491.960 696.000 493.360 ;
        RECT 3.070 487.920 696.000 491.960 ;
        RECT 4.400 486.520 696.000 487.920 ;
        RECT 3.070 482.480 696.000 486.520 ;
        RECT 4.400 481.080 696.000 482.480 ;
        RECT 3.070 477.040 696.000 481.080 ;
        RECT 4.400 475.640 696.000 477.040 ;
        RECT 3.070 471.600 696.000 475.640 ;
        RECT 4.400 470.240 696.000 471.600 ;
        RECT 4.400 470.200 695.600 470.240 ;
        RECT 3.070 468.840 695.600 470.200 ;
        RECT 3.070 466.160 696.000 468.840 ;
        RECT 4.400 464.760 696.000 466.160 ;
        RECT 3.070 460.720 696.000 464.760 ;
        RECT 4.400 459.320 696.000 460.720 ;
        RECT 3.070 455.280 696.000 459.320 ;
        RECT 4.400 453.880 696.000 455.280 ;
        RECT 3.070 449.840 696.000 453.880 ;
        RECT 4.400 448.440 696.000 449.840 ;
        RECT 3.070 444.400 696.000 448.440 ;
        RECT 4.400 443.000 696.000 444.400 ;
        RECT 3.070 440.320 696.000 443.000 ;
        RECT 3.070 438.960 695.600 440.320 ;
        RECT 4.400 438.920 695.600 438.960 ;
        RECT 4.400 437.560 696.000 438.920 ;
        RECT 3.070 433.520 696.000 437.560 ;
        RECT 4.400 432.120 696.000 433.520 ;
        RECT 3.070 428.080 696.000 432.120 ;
        RECT 4.400 426.680 696.000 428.080 ;
        RECT 3.070 422.640 696.000 426.680 ;
        RECT 4.400 421.240 696.000 422.640 ;
        RECT 3.070 417.200 696.000 421.240 ;
        RECT 4.400 415.800 696.000 417.200 ;
        RECT 3.070 411.760 696.000 415.800 ;
        RECT 4.400 410.400 696.000 411.760 ;
        RECT 4.400 410.360 695.600 410.400 ;
        RECT 3.070 409.000 695.600 410.360 ;
        RECT 3.070 406.320 696.000 409.000 ;
        RECT 4.400 404.920 696.000 406.320 ;
        RECT 3.070 400.880 696.000 404.920 ;
        RECT 4.400 399.480 696.000 400.880 ;
        RECT 3.070 395.440 696.000 399.480 ;
        RECT 4.400 394.040 696.000 395.440 ;
        RECT 3.070 390.000 696.000 394.040 ;
        RECT 4.400 388.600 696.000 390.000 ;
        RECT 3.070 384.560 696.000 388.600 ;
        RECT 4.400 383.160 696.000 384.560 ;
        RECT 3.070 380.480 696.000 383.160 ;
        RECT 3.070 379.120 695.600 380.480 ;
        RECT 4.400 379.080 695.600 379.120 ;
        RECT 4.400 377.720 696.000 379.080 ;
        RECT 3.070 373.680 696.000 377.720 ;
        RECT 4.400 372.280 696.000 373.680 ;
        RECT 3.070 368.240 696.000 372.280 ;
        RECT 4.400 366.840 696.000 368.240 ;
        RECT 3.070 362.800 696.000 366.840 ;
        RECT 4.400 361.400 696.000 362.800 ;
        RECT 3.070 357.360 696.000 361.400 ;
        RECT 4.400 355.960 696.000 357.360 ;
        RECT 3.070 351.920 696.000 355.960 ;
        RECT 4.400 350.560 696.000 351.920 ;
        RECT 4.400 350.520 695.600 350.560 ;
        RECT 3.070 349.160 695.600 350.520 ;
        RECT 3.070 346.480 696.000 349.160 ;
        RECT 4.400 345.080 696.000 346.480 ;
        RECT 3.070 341.040 696.000 345.080 ;
        RECT 4.400 339.640 696.000 341.040 ;
        RECT 3.070 335.600 696.000 339.640 ;
        RECT 4.400 334.200 696.000 335.600 ;
        RECT 3.070 330.160 696.000 334.200 ;
        RECT 4.400 328.760 696.000 330.160 ;
        RECT 3.070 324.720 696.000 328.760 ;
        RECT 4.400 323.320 696.000 324.720 ;
        RECT 3.070 320.640 696.000 323.320 ;
        RECT 3.070 319.280 695.600 320.640 ;
        RECT 4.400 319.240 695.600 319.280 ;
        RECT 4.400 317.880 696.000 319.240 ;
        RECT 3.070 313.840 696.000 317.880 ;
        RECT 4.400 312.440 696.000 313.840 ;
        RECT 3.070 308.400 696.000 312.440 ;
        RECT 4.400 307.000 696.000 308.400 ;
        RECT 3.070 302.960 696.000 307.000 ;
        RECT 4.400 301.560 696.000 302.960 ;
        RECT 3.070 297.520 696.000 301.560 ;
        RECT 4.400 296.120 696.000 297.520 ;
        RECT 3.070 292.080 696.000 296.120 ;
        RECT 4.400 290.720 696.000 292.080 ;
        RECT 4.400 290.680 695.600 290.720 ;
        RECT 3.070 289.320 695.600 290.680 ;
        RECT 3.070 286.640 696.000 289.320 ;
        RECT 4.400 285.240 696.000 286.640 ;
        RECT 3.070 281.200 696.000 285.240 ;
        RECT 4.400 279.800 696.000 281.200 ;
        RECT 3.070 275.760 696.000 279.800 ;
        RECT 4.400 274.360 696.000 275.760 ;
        RECT 3.070 270.320 696.000 274.360 ;
        RECT 4.400 268.920 696.000 270.320 ;
        RECT 3.070 264.880 696.000 268.920 ;
        RECT 4.400 263.480 696.000 264.880 ;
        RECT 3.070 260.800 696.000 263.480 ;
        RECT 3.070 259.440 695.600 260.800 ;
        RECT 4.400 259.400 695.600 259.440 ;
        RECT 4.400 258.040 696.000 259.400 ;
        RECT 3.070 254.000 696.000 258.040 ;
        RECT 4.400 252.600 696.000 254.000 ;
        RECT 3.070 248.560 696.000 252.600 ;
        RECT 4.400 247.160 696.000 248.560 ;
        RECT 3.070 243.120 696.000 247.160 ;
        RECT 4.400 241.720 696.000 243.120 ;
        RECT 3.070 237.680 696.000 241.720 ;
        RECT 4.400 236.280 696.000 237.680 ;
        RECT 3.070 232.240 696.000 236.280 ;
        RECT 4.400 230.880 696.000 232.240 ;
        RECT 4.400 230.840 695.600 230.880 ;
        RECT 3.070 229.480 695.600 230.840 ;
        RECT 3.070 226.800 696.000 229.480 ;
        RECT 4.400 225.400 696.000 226.800 ;
        RECT 3.070 221.360 696.000 225.400 ;
        RECT 4.400 219.960 696.000 221.360 ;
        RECT 3.070 215.920 696.000 219.960 ;
        RECT 4.400 214.520 696.000 215.920 ;
        RECT 3.070 210.480 696.000 214.520 ;
        RECT 4.400 209.080 696.000 210.480 ;
        RECT 3.070 205.040 696.000 209.080 ;
        RECT 4.400 203.640 696.000 205.040 ;
        RECT 3.070 200.960 696.000 203.640 ;
        RECT 3.070 199.600 695.600 200.960 ;
        RECT 4.400 199.560 695.600 199.600 ;
        RECT 4.400 198.200 696.000 199.560 ;
        RECT 3.070 194.160 696.000 198.200 ;
        RECT 4.400 192.760 696.000 194.160 ;
        RECT 3.070 188.720 696.000 192.760 ;
        RECT 4.400 187.320 696.000 188.720 ;
        RECT 3.070 183.280 696.000 187.320 ;
        RECT 4.400 181.880 696.000 183.280 ;
        RECT 3.070 177.840 696.000 181.880 ;
        RECT 4.400 176.440 696.000 177.840 ;
        RECT 3.070 172.400 696.000 176.440 ;
        RECT 4.400 171.040 696.000 172.400 ;
        RECT 4.400 171.000 695.600 171.040 ;
        RECT 3.070 169.640 695.600 171.000 ;
        RECT 3.070 166.960 696.000 169.640 ;
        RECT 4.400 165.560 696.000 166.960 ;
        RECT 3.070 161.520 696.000 165.560 ;
        RECT 4.400 160.120 696.000 161.520 ;
        RECT 3.070 156.080 696.000 160.120 ;
        RECT 4.400 154.680 696.000 156.080 ;
        RECT 3.070 150.640 696.000 154.680 ;
        RECT 4.400 149.240 696.000 150.640 ;
        RECT 3.070 145.200 696.000 149.240 ;
        RECT 4.400 143.800 696.000 145.200 ;
        RECT 3.070 141.120 696.000 143.800 ;
        RECT 3.070 139.760 695.600 141.120 ;
        RECT 4.400 139.720 695.600 139.760 ;
        RECT 4.400 138.360 696.000 139.720 ;
        RECT 3.070 134.320 696.000 138.360 ;
        RECT 4.400 132.920 696.000 134.320 ;
        RECT 3.070 128.880 696.000 132.920 ;
        RECT 4.400 127.480 696.000 128.880 ;
        RECT 3.070 123.440 696.000 127.480 ;
        RECT 4.400 122.040 696.000 123.440 ;
        RECT 3.070 118.000 696.000 122.040 ;
        RECT 4.400 116.600 696.000 118.000 ;
        RECT 3.070 112.560 696.000 116.600 ;
        RECT 4.400 111.200 696.000 112.560 ;
        RECT 4.400 111.160 695.600 111.200 ;
        RECT 3.070 109.800 695.600 111.160 ;
        RECT 3.070 107.120 696.000 109.800 ;
        RECT 4.400 105.720 696.000 107.120 ;
        RECT 3.070 101.680 696.000 105.720 ;
        RECT 4.400 100.280 696.000 101.680 ;
        RECT 3.070 96.240 696.000 100.280 ;
        RECT 4.400 94.840 696.000 96.240 ;
        RECT 3.070 90.800 696.000 94.840 ;
        RECT 4.400 89.400 696.000 90.800 ;
        RECT 3.070 85.360 696.000 89.400 ;
        RECT 4.400 83.960 696.000 85.360 ;
        RECT 3.070 81.280 696.000 83.960 ;
        RECT 3.070 79.920 695.600 81.280 ;
        RECT 4.400 79.880 695.600 79.920 ;
        RECT 4.400 78.520 696.000 79.880 ;
        RECT 3.070 51.360 696.000 78.520 ;
        RECT 3.070 49.960 695.600 51.360 ;
        RECT 3.070 21.440 696.000 49.960 ;
        RECT 3.070 20.040 695.600 21.440 ;
        RECT 3.070 9.695 696.000 20.040 ;
      LAYER met4 ;
        RECT 14.095 10.240 20.640 831.465 ;
        RECT 23.040 10.240 97.440 831.465 ;
        RECT 99.840 10.240 174.240 831.465 ;
        RECT 176.640 10.240 251.040 831.465 ;
        RECT 253.440 10.240 327.840 831.465 ;
        RECT 330.240 10.240 404.640 831.465 ;
        RECT 407.040 10.240 481.440 831.465 ;
        RECT 483.840 10.240 558.240 831.465 ;
        RECT 560.640 10.240 635.040 831.465 ;
        RECT 637.440 10.240 689.705 831.465 ;
        RECT 14.095 9.695 689.705 10.240 ;
  END
END icache
END LIBRARY

