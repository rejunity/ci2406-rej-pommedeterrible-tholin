magic
tech sky130B
magscale 1 2
timestamp 1717509706
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 566 2128 48912 48340
<< metal2 >>
rect 754 49200 810 50000
rect 2134 49200 2190 50000
rect 3514 49200 3570 50000
rect 4894 49200 4950 50000
rect 6274 49200 6330 50000
rect 7654 49200 7710 50000
rect 9034 49200 9090 50000
rect 10414 49200 10470 50000
rect 11794 49200 11850 50000
rect 13174 49200 13230 50000
rect 14554 49200 14610 50000
rect 15934 49200 15990 50000
rect 17314 49200 17370 50000
rect 18694 49200 18750 50000
rect 20074 49200 20130 50000
rect 21454 49200 21510 50000
rect 22834 49200 22890 50000
rect 24214 49200 24270 50000
rect 25594 49200 25650 50000
rect 26974 49200 27030 50000
rect 28354 49200 28410 50000
rect 29734 49200 29790 50000
rect 31114 49200 31170 50000
rect 32494 49200 32550 50000
rect 33874 49200 33930 50000
rect 35254 49200 35310 50000
rect 36634 49200 36690 50000
rect 38014 49200 38070 50000
rect 39394 49200 39450 50000
rect 40774 49200 40830 50000
rect 42154 49200 42210 50000
rect 43534 49200 43590 50000
rect 44914 49200 44970 50000
rect 46294 49200 46350 50000
rect 47674 49200 47730 50000
rect 49054 49200 49110 50000
<< obsm2 >>
rect 572 49144 698 49314
rect 866 49144 2078 49314
rect 2246 49144 3458 49314
rect 3626 49144 4838 49314
rect 5006 49144 6218 49314
rect 6386 49144 7598 49314
rect 7766 49144 8978 49314
rect 9146 49144 10358 49314
rect 10526 49144 11738 49314
rect 11906 49144 13118 49314
rect 13286 49144 14498 49314
rect 14666 49144 15878 49314
rect 16046 49144 17258 49314
rect 17426 49144 18638 49314
rect 18806 49144 20018 49314
rect 20186 49144 21398 49314
rect 21566 49144 22778 49314
rect 22946 49144 24158 49314
rect 24326 49144 25538 49314
rect 25706 49144 26918 49314
rect 27086 49144 28298 49314
rect 28466 49144 29678 49314
rect 29846 49144 31058 49314
rect 31226 49144 32438 49314
rect 32606 49144 33818 49314
rect 33986 49144 35198 49314
rect 35366 49144 36578 49314
rect 36746 49144 37958 49314
rect 38126 49144 39338 49314
rect 39506 49144 40718 49314
rect 40886 49144 42098 49314
rect 42266 49144 43478 49314
rect 43646 49144 44858 49314
rect 45026 49144 46238 49314
rect 46406 49144 47618 49314
rect 47786 49144 48648 49314
rect 572 2139 48648 49144
<< metal3 >>
rect 0 46520 800 46640
rect 0 45432 800 45552
rect 0 44344 800 44464
rect 49200 43528 50000 43648
rect 0 43256 800 43376
rect 0 42168 800 42288
rect 0 41080 800 41200
rect 0 39992 800 40112
rect 0 38904 800 39024
rect 0 37816 800 37936
rect 0 36728 800 36848
rect 0 35640 800 35760
rect 0 34552 800 34672
rect 0 33464 800 33584
rect 0 32376 800 32496
rect 0 31288 800 31408
rect 49200 31016 50000 31136
rect 0 30200 800 30320
rect 0 29112 800 29232
rect 0 28024 800 28144
rect 0 26936 800 27056
rect 0 25848 800 25968
rect 0 24760 800 24880
rect 0 23672 800 23792
rect 0 22584 800 22704
rect 0 21496 800 21616
rect 0 20408 800 20528
rect 0 19320 800 19440
rect 49200 18504 50000 18624
rect 0 18232 800 18352
rect 0 17144 800 17264
rect 0 16056 800 16176
rect 0 14968 800 15088
rect 0 13880 800 14000
rect 0 12792 800 12912
rect 0 11704 800 11824
rect 0 10616 800 10736
rect 0 9528 800 9648
rect 0 8440 800 8560
rect 0 7352 800 7472
rect 0 6264 800 6384
rect 49200 5992 50000 6112
rect 0 5176 800 5296
rect 0 4088 800 4208
rect 0 3000 800 3120
<< obsm3 >>
rect 790 46720 49200 47701
rect 880 46440 49200 46720
rect 790 45632 49200 46440
rect 880 45352 49200 45632
rect 790 44544 49200 45352
rect 880 44264 49200 44544
rect 790 43728 49200 44264
rect 790 43456 49120 43728
rect 880 43448 49120 43456
rect 880 43176 49200 43448
rect 790 42368 49200 43176
rect 880 42088 49200 42368
rect 790 41280 49200 42088
rect 880 41000 49200 41280
rect 790 40192 49200 41000
rect 880 39912 49200 40192
rect 790 39104 49200 39912
rect 880 38824 49200 39104
rect 790 38016 49200 38824
rect 880 37736 49200 38016
rect 790 36928 49200 37736
rect 880 36648 49200 36928
rect 790 35840 49200 36648
rect 880 35560 49200 35840
rect 790 34752 49200 35560
rect 880 34472 49200 34752
rect 790 33664 49200 34472
rect 880 33384 49200 33664
rect 790 32576 49200 33384
rect 880 32296 49200 32576
rect 790 31488 49200 32296
rect 880 31216 49200 31488
rect 880 31208 49120 31216
rect 790 30936 49120 31208
rect 790 30400 49200 30936
rect 880 30120 49200 30400
rect 790 29312 49200 30120
rect 880 29032 49200 29312
rect 790 28224 49200 29032
rect 880 27944 49200 28224
rect 790 27136 49200 27944
rect 880 26856 49200 27136
rect 790 26048 49200 26856
rect 880 25768 49200 26048
rect 790 24960 49200 25768
rect 880 24680 49200 24960
rect 790 23872 49200 24680
rect 880 23592 49200 23872
rect 790 22784 49200 23592
rect 880 22504 49200 22784
rect 790 21696 49200 22504
rect 880 21416 49200 21696
rect 790 20608 49200 21416
rect 880 20328 49200 20608
rect 790 19520 49200 20328
rect 880 19240 49200 19520
rect 790 18704 49200 19240
rect 790 18432 49120 18704
rect 880 18424 49120 18432
rect 880 18152 49200 18424
rect 790 17344 49200 18152
rect 880 17064 49200 17344
rect 790 16256 49200 17064
rect 880 15976 49200 16256
rect 790 15168 49200 15976
rect 880 14888 49200 15168
rect 790 14080 49200 14888
rect 880 13800 49200 14080
rect 790 12992 49200 13800
rect 880 12712 49200 12992
rect 790 11904 49200 12712
rect 880 11624 49200 11904
rect 790 10816 49200 11624
rect 880 10536 49200 10816
rect 790 9728 49200 10536
rect 880 9448 49200 9728
rect 790 8640 49200 9448
rect 880 8360 49200 8640
rect 790 7552 49200 8360
rect 880 7272 49200 7552
rect 790 6464 49200 7272
rect 880 6192 49200 6464
rect 880 6184 49120 6192
rect 790 5912 49120 6184
rect 790 5376 49200 5912
rect 880 5096 49200 5376
rect 790 4288 49200 5096
rect 880 4008 49200 4288
rect 790 3200 49200 4008
rect 880 2920 49200 3200
rect 790 2143 49200 2920
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 795 47456 44285 47701
rect 795 5611 4128 47456
rect 4608 5611 19488 47456
rect 19968 5611 34848 47456
rect 35328 5611 44285 47456
<< labels >>
rlabel metal3 s 49200 31016 50000 31136 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 49200 43528 50000 43648 6 custom_settings[1]
port 2 nsew signal input
rlabel metal2 s 754 49200 810 50000 6 io_in[0]
port 3 nsew signal input
rlabel metal2 s 14554 49200 14610 50000 6 io_in[10]
port 4 nsew signal input
rlabel metal2 s 15934 49200 15990 50000 6 io_in[11]
port 5 nsew signal input
rlabel metal2 s 17314 49200 17370 50000 6 io_in[12]
port 6 nsew signal input
rlabel metal2 s 18694 49200 18750 50000 6 io_in[13]
port 7 nsew signal input
rlabel metal2 s 20074 49200 20130 50000 6 io_in[14]
port 8 nsew signal input
rlabel metal2 s 21454 49200 21510 50000 6 io_in[15]
port 9 nsew signal input
rlabel metal2 s 22834 49200 22890 50000 6 io_in[16]
port 10 nsew signal input
rlabel metal2 s 24214 49200 24270 50000 6 io_in[17]
port 11 nsew signal input
rlabel metal2 s 25594 49200 25650 50000 6 io_in[18]
port 12 nsew signal input
rlabel metal2 s 26974 49200 27030 50000 6 io_in[19]
port 13 nsew signal input
rlabel metal2 s 2134 49200 2190 50000 6 io_in[1]
port 14 nsew signal input
rlabel metal2 s 28354 49200 28410 50000 6 io_in[20]
port 15 nsew signal input
rlabel metal2 s 29734 49200 29790 50000 6 io_in[21]
port 16 nsew signal input
rlabel metal2 s 31114 49200 31170 50000 6 io_in[22]
port 17 nsew signal input
rlabel metal2 s 32494 49200 32550 50000 6 io_in[23]
port 18 nsew signal input
rlabel metal2 s 33874 49200 33930 50000 6 io_in[24]
port 19 nsew signal input
rlabel metal2 s 35254 49200 35310 50000 6 io_in[25]
port 20 nsew signal input
rlabel metal2 s 36634 49200 36690 50000 6 io_in[26]
port 21 nsew signal input
rlabel metal2 s 38014 49200 38070 50000 6 io_in[27]
port 22 nsew signal input
rlabel metal2 s 39394 49200 39450 50000 6 io_in[28]
port 23 nsew signal input
rlabel metal2 s 40774 49200 40830 50000 6 io_in[29]
port 24 nsew signal input
rlabel metal2 s 3514 49200 3570 50000 6 io_in[2]
port 25 nsew signal input
rlabel metal2 s 42154 49200 42210 50000 6 io_in[30]
port 26 nsew signal input
rlabel metal2 s 43534 49200 43590 50000 6 io_in[31]
port 27 nsew signal input
rlabel metal2 s 44914 49200 44970 50000 6 io_in[32]
port 28 nsew signal input
rlabel metal2 s 46294 49200 46350 50000 6 io_in[33]
port 29 nsew signal input
rlabel metal2 s 47674 49200 47730 50000 6 io_in[34]
port 30 nsew signal input
rlabel metal2 s 49054 49200 49110 50000 6 io_in[35]
port 31 nsew signal input
rlabel metal2 s 4894 49200 4950 50000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6274 49200 6330 50000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 7654 49200 7710 50000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 9034 49200 9090 50000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 10414 49200 10470 50000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 11794 49200 11850 50000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 13174 49200 13230 50000 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_oeb[1]
port 40 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 io_oeb[2]
port 41 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 io_oeb[3]
port 42 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 io_oeb[4]
port 43 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 io_out[0]
port 44 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_out[10]
port 45 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_out[11]
port 46 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 io_out[12]
port 47 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 io_out[13]
port 48 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 io_out[14]
port 49 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 io_out[15]
port 50 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_out[16]
port 51 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 io_out[17]
port 52 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 io_out[18]
port 53 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 io_out[19]
port 54 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 io_out[1]
port 55 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 io_out[20]
port 56 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 io_out[21]
port 57 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 io_out[22]
port 58 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 io_out[23]
port 59 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 io_out[24]
port 60 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 io_out[25]
port 61 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_out[26]
port 62 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 io_out[27]
port 63 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 io_out[28]
port 64 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 io_out[29]
port 65 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 io_out[2]
port 66 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 io_out[30]
port 67 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 io_out[31]
port 68 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 io_out[32]
port 69 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 io_out[33]
port 70 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 io_out[34]
port 71 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 io_out[35]
port 72 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 io_out[3]
port 73 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_out[4]
port 74 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_out[5]
port 75 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 io_out[6]
port 76 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 io_out[7]
port 77 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 io_out[8]
port 78 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 io_out[9]
port 79 nsew signal output
rlabel metal3 s 49200 18504 50000 18624 6 rst_n
port 80 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 81 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 81 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 82 nsew ground bidirectional
rlabel metal3 s 49200 5992 50000 6112 6 wb_clk_i
port 83 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9415258
string GDS_FILE /home/lucah/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/S8x305/runs/24_06_04_15_47/results/signoff/wrapped_8x305.magic.gds
string GDS_START 1020860
<< end >>

