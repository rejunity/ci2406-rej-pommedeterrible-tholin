* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_mask[0]
+ dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0] dest_val[10]
+ dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16] dest_val[17]
+ dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22] dest_val[23]
+ dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29] dest_val[2]
+ dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6] dest_val[7]
+ dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11] instruction[12]
+ instruction[13] instruction[14] instruction[15] instruction[16] instruction[17]
+ instruction[18] instruction[19] instruction[1] instruction[20] instruction[21] instruction[22]
+ instruction[23] instruction[24] instruction[25] instruction[26] instruction[27]
+ instruction[28] instruction[29] instruction[2] instruction[30] instruction[31] instruction[32]
+ instruction[33] instruction[34] instruction[35] instruction[36] instruction[37]
+ instruction[38] instruction[39] instruction[3] instruction[40] instruction[41] instruction[4]
+ instruction[5] instruction[6] instruction[7] instruction[8] instruction[9] int_return
+ is_load is_store loadstore_address[0] loadstore_address[10] loadstore_address[11]
+ loadstore_address[12] loadstore_address[13] loadstore_address[14] loadstore_address[15]
+ loadstore_address[16] loadstore_address[17] loadstore_address[18] loadstore_address[19]
+ loadstore_address[1] loadstore_address[20] loadstore_address[21] loadstore_address[22]
+ loadstore_address[23] loadstore_address[24] loadstore_address[25] loadstore_address[26]
+ loadstore_address[27] loadstore_address[28] loadstore_address[29] loadstore_address[2]
+ loadstore_address[30] loadstore_address[31] loadstore_address[3] loadstore_address[4]
+ loadstore_address[5] loadstore_address[6] loadstore_address[7] loadstore_address[8]
+ loadstore_address[9] loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3]
+ loadstore_dest[4] loadstore_size[0] loadstore_size[1] new_PC[0] new_PC[10] new_PC[11]
+ new_PC[12] new_PC[13] new_PC[14] new_PC[15] new_PC[16] new_PC[17] new_PC[18] new_PC[19]
+ new_PC[1] new_PC[20] new_PC[21] new_PC[22] new_PC[23] new_PC[24] new_PC[25] new_PC[26]
+ new_PC[27] new_PC[2] new_PC[3] new_PC[4] new_PC[5] new_PC[6] new_PC[7] new_PC[8]
+ new_PC[9] pred_idx[0] pred_idx[1] pred_idx[2] pred_val reg1_idx[0] reg1_idx[1] reg1_idx[2]
+ reg1_idx[3] reg1_idx[4] reg1_val[0] reg1_val[10] reg1_val[11] reg1_val[12] reg1_val[13]
+ reg1_val[14] reg1_val[15] reg1_val[16] reg1_val[17] reg1_val[18] reg1_val[19] reg1_val[1]
+ reg1_val[20] reg1_val[21] reg1_val[22] reg1_val[23] reg1_val[24] reg1_val[25] reg1_val[26]
+ reg1_val[27] reg1_val[28] reg1_val[29] reg1_val[2] reg1_val[30] reg1_val[31] reg1_val[3]
+ reg1_val[4] reg1_val[5] reg1_val[6] reg1_val[7] reg1_val[8] reg1_val[9] reg2_idx[0]
+ reg2_idx[1] reg2_idx[2] reg2_idx[3] reg2_idx[4] reg2_val[0] reg2_val[10] reg2_val[11]
+ reg2_val[12] reg2_val[13] reg2_val[14] reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18]
+ reg2_val[19] reg2_val[1] reg2_val[20] reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24]
+ reg2_val[25] reg2_val[26] reg2_val[27] reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30]
+ reg2_val[31] reg2_val[3] reg2_val[4] reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8]
+ reg2_val[9] rst sign_extend take_branch vccd1 vssd1 wb_clk_i
X_06883_ _09743_/A _06880_/X _06883_/C _06883_/D vssd1 vssd1 vccd1 vccd1 _06884_/D
+ sky130_fd_sc_hd__and4bb_1
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09673_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08622_ _08622_/A _08622_/B _08620_/Y vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08553_ _08649_/B _08553_/A2 _08553_/B1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08554_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout162_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _08633_/B fanout52/X fanout50/X _09300_/A vssd1 vssd1 vccd1 vccd1 _07505_/B
+ sky130_fd_sc_hd__o22a_1
X_08484_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08484_/X sky130_fd_sc_hd__and2_1
XANTENNA__12830__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ _09787_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12043__A0 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07366_ _11168_/A _07366_/B vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__xnor2_1
X_09105_ _09106_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09105_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07297_ _08650_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07310_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ _09371_/A _09371_/C _09034_/Y vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08014__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout75_A _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _06785_/X _09595_/A _09740_/X _06787_/B vssd1 vssd1 vccd1 vccd1 _09870_/B
+ sky130_fd_sc_hd__a31o_1
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13059__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12880_ hold317/A hold21/X vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__nand2b_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11746_/A _11746_/B _11737_/A vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12806__C1 _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13074__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07289__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11764_/C sky130_fd_sc_hd__xnor2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10715_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _11693_/A _11693_/B vssd1 vssd1 vccd1 vccd1 _11693_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _10645_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10646_/A sky130_fd_sc_hd__or2_2
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13363_ _13363_/CLK _13363_/D vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
X_10575_ _07968_/B _07151_/A _07155_/A _07077_/X vssd1 vssd1 vccd1 vccd1 _10576_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12314_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09450__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07461__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _13352_/CLK hold227/X vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10348__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ _06626_/X _12243_/Y _12244_/X vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12176_ hold188/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__or2_1
XANTENNA__06602__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__A1 _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11018_/B _11020_/B _11018_/A vssd1 vssd1 vccd1 vccd1 _11128_/B sky130_fd_sc_hd__a21bo_1
X_11058_ _12143_/A fanout31/X fanout29/X _06978_/X vssd1 vssd1 vccd1 vccd1 _11059_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10009_ _11021_/S _09569_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09808__A3 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07220_ _09795_/A _07220_/B vssd1 vssd1 vccd1 vccd1 _07221_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ _07151_/A vssd1 vssd1 vccd1 vccd1 _07151_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _07082_/A _07082_/B vssd1 vssd1 vccd1 vccd1 _07360_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11551__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout105 _10227_/B1 vssd1 vssd1 vccd1 vccd1 _10463_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout138 _10613_/A vssd1 vssd1 vccd1 vccd1 _10468_/A sky130_fd_sc_hd__buf_12
Xfanout116 _07178_/Y vssd1 vssd1 vccd1 vccd1 _10585_/B2 sky130_fd_sc_hd__buf_8
Xfanout127 _07115_/Y vssd1 vssd1 vccd1 vccd1 _08553_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07755__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout149 _07017_/X vssd1 vssd1 vccd1 vccd1 _09297_/A1 sky130_fd_sc_hd__buf_4
X_07984_ _07873_/A _07873_/B _07873_/C vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__o21ai_1
X_06935_ instruction[7] is_load _06706_/A _06932_/X vssd1 vssd1 vccd1 vccd1 _06936_/B
+ sky130_fd_sc_hd__a22o_2
X_09723_ _09249_/A _09722_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06866_ _12098_/A _06865_/X _06854_/X vssd1 vssd1 vccd1 vccd1 _06866_/X sky130_fd_sc_hd__a21o_1
X_09654_ fanout55/X _10233_/B2 _10233_/A1 fanout67/X vssd1 vssd1 vccd1 vccd1 _09655_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09542__B _09543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08605_/A _08605_/B _08605_/C vssd1 vssd1 vccd1 vccd1 _08607_/C sky130_fd_sc_hd__and3_1
XANTENNA__13056__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06797_ _12621_/A _09722_/S vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__or2_1
X_09585_ _12621_/A _09722_/S _09396_/S _09219_/A vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08536_ _08536_/A _08536_/B vssd1 vssd1 vccd1 vccd1 _08546_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _09941_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08472_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07418_ _07418_/A _07418_/B vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08398_ _08591_/B1 _10227_/B1 _10463_/A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 _08399_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _07348_/A _07348_/B _07573_/A vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__o21bai_1
X_10360_ _10942_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10291_ hold247/A _10427_/A2 _10554_/C _12433_/A1 vssd1 vssd1 vccd1 vccd1 _10291_/X
+ sky130_fd_sc_hd__a31o_1
X_09019_ _08881_/A _08881_/B _08879_/X vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold170 hold172/X vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__A2 _09728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A0 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _12420_/A _08791_/A _08791_/B _12029_/Y vssd1 vssd1 vccd1 vccd1 _12030_/Y
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__12143__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09499__A1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ hold101/X hold316/A vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10502__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11058__A1 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ hold86/X hold275/X vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09879__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__B2 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _07031_/X fanout40/X _07301_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _11815_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _07114_/X _13078_/B2 hold105/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13246_/D
+ sky130_fd_sc_hd__o211a_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__or2_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10805__A1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _11677_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09423__B2 _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08226__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ _13346_/CLK _13346_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
X_10558_ hold283/A hold313/A _10558_/C vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__or3_1
XANTENNA__07434__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10553__S _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ _13297_/CLK _13277_/D vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _10624_/B _10489_/B vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12228_ _12420_/A _08798_/X _12229_/B vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__a21bo_1
X_12159_ _12158_/A _12279_/C _09149_/X vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11297__A1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _11125_/A _07251_/A vssd1 vssd1 vccd1 vccd1 _11137_/S sky130_fd_sc_hd__and2_1
X_06651_ _07026_/B reg1_val[26] vssd1 vssd1 vccd1 vccd1 _12179_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13038__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06582_ instruction[19] _06922_/B vssd1 vssd1 vccd1 vccd1 _06582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09370_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__xnor2_4
X_08321_ _08605_/A _10222_/A2 _07255_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _08322_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07673__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _07944_/B _10326_/A fanout28/X _09450_/B1 vssd1 vssd1 vccd1 vccd1 _07204_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _08183_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__xor2_2
X_07134_ reg1_val[26] _07134_/B vssd1 vssd1 vccd1 vccd1 _07135_/C sky130_fd_sc_hd__xor2_2
XANTENNA__10024__A2 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07065_ reg1_val[8] _07085_/D _07093_/A vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10699__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _07060_/A _07060_/B _06875_/A vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__a21o_1
X_06918_ instruction[27] _06922_/B vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__or2_1
XANTENNA__06896__B _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _09706_/A _09858_/A _09996_/A _10128_/A vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__or4_1
X_07898_ _07010_/Y _07968_/B _07077_/X _07018_/X vssd1 vssd1 vccd1 vccd1 _07899_/B
+ sky130_fd_sc_hd__a22o_1
X_06849_ reg1_val[30] _08858_/A vssd1 vssd1 vccd1 vccd1 _06849_/Y sky130_fd_sc_hd__nand2_1
X_09637_ _09843_/B _09637_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nand2_1
X_09568_ _09190_/X _09194_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout38_A _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__A1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08542_/B sky130_fd_sc_hd__nor2_1
X_11530_ _11529_/B _11620_/B hold255/A vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__a21o_1
X_09499_ _09671_/A _07010_/B wire8/X _09498_/Y vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__a31o_2
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout4_A fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11461_ _12143_/A _07151_/A _07155_/A _06978_/X vssd1 vssd1 vccd1 vccd1 _11462_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__B _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11392_ _11392_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__nor2_1
X_13200_ hold269/X _13209_/A2 _13199_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold270/A
+ sky130_fd_sc_hd__a22o_1
X_10412_ _06757_/Y _10277_/Y _06759_/B vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _13131_/A _13131_/B vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__xnor2_1
X_10343_ _10235_/A _10237_/B _10344_/B vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07967__A1 _07060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07248__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13062_ _11900_/A _13072_/A2 hold124/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__o21a_1
X_10274_ _10175_/X _10570_/A _10273_/Y vssd1 vssd1 vccd1 vccd1 _10274_/Y sky130_fd_sc_hd__a21oi_1
X_12013_ _11852_/A _11935_/A _11934_/A vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__a21o_1
X_12915_ hold80/X hold311/X vssd1 vssd1 vccd1 vccd1 _13150_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ _08857_/Y _13072_/A2 hold69/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold70/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12778_/B vssd1 vssd1 vccd1 vccd1 _12777_/Y sky130_fd_sc_hd__inv_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11728_ _07031_/X fanout42/X fanout40/X _12143_/A vssd1 vssd1 vccd1 vccd1 _11729_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _11658_/B _11659_/B vssd1 vssd1 vccd1 vccd1 _11660_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07407__B1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ _13334_/CLK hold125/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12951__B2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12064__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ reg1_val[30] _08870_/B vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09580__B1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _07821_/A _07821_/B _07821_/C vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__or3_2
XFILLER_0_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07752_ _12785_/A fanout45/X _09324_/A _07814_/B vssd1 vssd1 vccd1 vccd1 _07753_/B
+ sky130_fd_sc_hd__o22a_2
X_06703_ reg1_val[17] _11446_/A vssd1 vssd1 vccd1 vccd1 _06704_/B sky130_fd_sc_hd__nand2b_1
X_07683_ fanout60/X _08649_/B _08641_/A2 fanout52/X vssd1 vssd1 vccd1 vccd1 _07684_/B
+ sky130_fd_sc_hd__o22a_1
X_06634_ reg1_val[25] _06978_/A vssd1 vssd1 vccd1 vccd1 _06635_/B sky130_fd_sc_hd__and2b_1
X_09422_ hold265/A _13338_/Q _10158_/A2 _09240_/X vssd1 vssd1 vccd1 vccd1 _09422_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10966__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _09353_/A _09353_/B vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__and2_1
XANTENNA__07621__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ instruction[3] vssd1 vssd1 vccd1 vccd1 _06927_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _08301_/A _08301_/B _08303_/Y vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__B2 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _09285_/A _09285_/B vssd1 vssd1 vccd1 vccd1 _09284_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08235_ _08300_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13195__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08166_/X sky130_fd_sc_hd__and2b_1
X_07117_ _07116_/B _11823_/A _11900_/A vssd1 vssd1 vccd1 vccd1 _07117_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08097_ _08591_/B1 _08184_/B fanout32/X _08619_/B1 vssd1 vssd1 vccd1 vccd1 _08098_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07068__A _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _10061_/A _07048_/B vssd1 vssd1 vccd1 vccd1 _07048_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__06700__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__B _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__xor2_1
X_10961_ _11188_/A fanout9/X fanout4/X _11083_/A vssd1 vssd1 vccd1 vccd1 _10962_/B
+ sky130_fd_sc_hd__o22a_1
X_12700_ reg1_val[16] _12767_/B vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__xor2_4
X_10892_ _11110_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12631_ reg1_val[3] _12632_/B vssd1 vssd1 vccd1 vccd1 _12631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ _12574_/A _12574_/B _12575_/B vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11988__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _12502_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12495_/C sky130_fd_sc_hd__nand2_1
X_11513_ _11781_/S _11513_/B vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13186__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _11423_/X _11424_/Y _11428_/Y _11612_/A _11443_/X vssd1 vssd1 vccd1 vccd1
+ _11444_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11375_ _11375_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _13236_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13345_/D sky130_fd_sc_hd__and2_1
X_10326_ _10326_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__nand2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10258_/A _10258_/B vssd1 vssd1 vccd1 vccd1 _10257_/X sky130_fd_sc_hd__and2b_1
X_13045_ hold152/X _13071_/A2 _13071_/B1 hold170/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold173/A sky130_fd_sc_hd__o221a_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06610__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _11359_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10189_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__B _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ hold77/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_1
XANTENNA__12059__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10227__A2 _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09093__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11898__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ _08020_/A _08020_/B vssd1 vssd1 vccd1 vccd1 _08065_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12506__B _12506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout7 fanout7/A vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__buf_6
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09821_/A _09821_/B _09819_/Y vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__09815__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ _09038_/A _09038_/B _12383_/A vssd1 vssd1 vccd1 vccd1 _12420_/B sky130_fd_sc_hd__or3_1
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07616__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08853_ _08941_/B _08853_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nand2_1
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07858_/B sky130_fd_sc_hd__xnor2_1
X_08784_ _08060_/A _08060_/B _08165_/Y vssd1 vssd1 vccd1 vccd1 _08784_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07735_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _09401_/X _09404_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09405_/X sky130_fd_sc_hd__mux2_1
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08447__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06617_ _06706_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _06617_/Y sky130_fd_sc_hd__nor2_1
X_07597_ _09668_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10218__A2 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09336_ _09048_/Y _09051_/B _09056_/A vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09084__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _09766_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _09268_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08292__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08218_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _09194_/X _09197_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10217__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ _08147_/A _08147_/B _08148_/Y vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__a21bo_1
X_11160_ _11305_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11091_ _10976_/B _10976_/C _10976_/A vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__a21bo_1
X_10111_ _09978_/A _09977_/B _09975_/Y vssd1 vssd1 vccd1 vccd1 _10121_/A sky130_fd_sc_hd__a21o_1
X_10042_ _09950_/Y _09952_/Y _07263_/Y _11645_/B vssd1 vssd1 vccd1 vccd1 _10042_/X
+ sky130_fd_sc_hd__o211a_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _12073_/A _11993_/B vssd1 vssd1 vccd1 vccd1 _11995_/B sky130_fd_sc_hd__or2_1
XANTENNA__12300__C1 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ _11169_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07322__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ _10753_/A _10753_/B _10751_/Y vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12614_ _12611_/B _12613_/B _12611_/A vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _12549_/B _12545_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08283__B1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11511__A _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12476_ reg1_val[6] curr_PC[6] _12504_/S vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11427_ _11781_/S _06834_/X _11426_/Y vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__o21a_1
XANTENNA_5 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ fanout29/X _07301_/Y _07593_/Y fanout31/X vssd1 vssd1 vccd1 vccd1 _11359_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09916__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _12490_/S _10306_/X _10307_/X _10308_/Y vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a22o_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _11288_/B _11289_/B vssd1 vssd1 vccd1 vccd1 _11290_/B sky130_fd_sc_hd__and2b_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _07053_/B _12797_/B hold177/X vssd1 vssd1 vccd1 vccd1 _13312_/D sky130_fd_sc_hd__a21boi_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _07520_/A _07520_/B vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10448__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09370__B _09370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07451_ _07451_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07480_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07382_ _09795_/A _07382_/B vssd1 vssd1 vccd1 vccd1 _07419_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11948__A2 _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _08996_/A _08996_/B _08994_/X vssd1 vssd1 vccd1 vccd1 _09123_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13112__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09052_ _07101_/Y fanout41/X _07263_/Y _07402_/B vssd1 vssd1 vccd1 vccd1 _09053_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08003_ _08573_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout205_A _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09955_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07346__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ hold261/A _10427_/A2 _10153_/C _09884_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _09885_/X sky130_fd_sc_hd__a311o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _08905_/A _08905_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__xnor2_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _10231_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _08838_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07001__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08767_ _08776_/B _08767_/B _08767_/C vssd1 vssd1 vccd1 vccd1 _08769_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08177__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _07718_/A _07718_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07719_/B sky130_fd_sc_hd__nand3_1
X_08698_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _07647_/A _07647_/B _07650_/B vssd1 vssd1 vccd1 vccd1 _07649_/X sky130_fd_sc_hd__o21ba_1
X_10660_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10660_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout20_A _08985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _09320_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _11645_/A fanout46/X fanout44/X fanout51/X vssd1 vssd1 vccd1 vccd1 _10592_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12061__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12330_/A _12330_/B _12374_/D vssd1 vssd1 vccd1 vccd1 _12330_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ _12262_/A _12315_/A vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__nor2_1
X_11212_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11214_/C sky130_fd_sc_hd__xor2_2
XANTENNA__09765__B1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__A1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__B2 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _11131_/A _09406_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__o21ai_2
X_11074_ _11074_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__and2_1
X_10025_ _09895_/A _09892_/Y _09894_/B vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11627__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _11975_/A _11972_/X _11973_/X _11975_/Y vssd1 vssd1 vccd1 vccd1 dest_val[23]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ curr_PC[12] _10808_/B _12053_/A1 vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10724_/A _10724_/B _10720_/X vssd1 vssd1 vccd1 vccd1 _10860_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08815__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _09874_/Y _10788_/Y _11237_/S vssd1 vssd1 vccd1 vccd1 _10789_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ _12537_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _12530_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13001__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ _12460_/A _12460_/B _12460_/C vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__A _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06951_ _07145_/A _07152_/A _07129_/A _08476_/A vssd1 vssd1 vccd1 vccd1 _07113_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__09508__B1 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _09670_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06882_ _08655_/A _06876_/Y _10414_/A _06793_/Y _09419_/A vssd1 vssd1 vccd1 vccd1
+ _06883_/D sky130_fd_sc_hd__o2111a_1
X_08621_ _08622_/A _08622_/B _08620_/Y vssd1 vssd1 vccd1 vccd1 _08629_/A sky130_fd_sc_hd__nor3b_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13107__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08552_ _08566_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08585_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07298__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07503_ _07503_/A _07503_/B vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__xnor2_1
X_08483_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07434_ _08354_/A2 _10466_/A fanout71/X fanout85/X vssd1 vssd1 vccd1 vccd1 _07435_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ _08354_/A2 fanout77/X fanout73/X _10327_/B2 vssd1 vssd1 vccd1 vccd1 _07366_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11151__A _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _11645_/B _09104_/B vssd1 vssd1 vccd1 vccd1 _09106_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ fanout67/X _09297_/B2 _09297_/A1 fanout64/X vssd1 vssd1 vccd1 vccd1 _07297_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _09035_/A _09544_/A vssd1 vssd1 vccd1 vccd1 _09371_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07076__A _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09648_/A fanout11/X fanout7/X _08590_/B vssd1 vssd1 vccd1 vccd1 _09938_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout68_A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _12420_/A _08713_/A _08713_/B _11946_/A _09867_/Y vssd1 vssd1 vccd1 vccd1
+ _09868_/Y sky130_fd_sc_hd__a311oi_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__nor2_1
X_08819_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__nor2_1
X_11830_ _11830_/A _11830_/B vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10230__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11850_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07289__B2 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07289__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10712_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11863_/A _11692_/B vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08238__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10574_ _12310_/A _10574_/B vssd1 vssd1 vccd1 vccd1 _10578_/A sky130_fd_sc_hd__xnor2_2
X_13362_ _13372_/CLK _13362_/D vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _12313_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09450__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__A1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13293_ _13352_/CLK hold239/X vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07461__B2 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10348__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ _07029_/A _11446_/B _09235_/X _06628_/B _11975_/A vssd1 vssd1 vccd1 vccd1
+ _12244_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12175_ hold329/A _12175_/A2 _12239_/B _12174_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _12183_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06602__B _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11128_/A sky130_fd_sc_hd__nand2_1
X_11057_ _11057_/A _11057_/B vssd1 vssd1 vccd1 vccd1 _11060_/A sky130_fd_sc_hd__and2_1
XANTENNA__09910__B1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _10008_/A _10008_/B vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _11958_/A _10434_/Y _11958_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _11971_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10286__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _07150_/A _07150_/B vssd1 vssd1 vccd1 vccd1 _07150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07081_ _07427_/A _07427_/B vssd1 vssd1 vccd1 vccd1 _07428_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08280__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout106 _07282_/Y vssd1 vssd1 vccd1 vccd1 _10227_/B1 sky130_fd_sc_hd__buf_8
Xfanout128 _07115_/Y vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07755__A2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _09394_/X _09396_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09722_/X sky130_fd_sc_hd__mux2_1
X_07983_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _07993_/A sky130_fd_sc_hd__nand2b_1
X_06934_ _11975_/A _06934_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
X_06865_ _06655_/B _06848_/B _06855_/X vssd1 vssd1 vccd1 vccd1 _06865_/X sky130_fd_sc_hd__a21o_1
X_09653_ _09653_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__nor2_1
X_09584_ hold325/A _10427_/A2 _09582_/X _12433_/A1 vssd1 vssd1 vccd1 vccd1 _09584_/X
+ sky130_fd_sc_hd__a31o_1
X_08604_ _07101_/A _07101_/B _06973_/A vssd1 vssd1 vccd1 vccd1 _08607_/B sky130_fd_sc_hd__a21oi_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06796_ _06799_/A _06801_/B1 _12627_/B _06794_/X vssd1 vssd1 vccd1 vccd1 _06796_/X
+ sky130_fd_sc_hd__a31o_1
X_08535_ _08562_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08466_ _08619_/A2 _08553_/A2 _08551_/B1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 _08467_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07140__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07417_ _07662_/A _07416_/B _07388_/Y vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__a21o_1
X_08397_ _08397_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _08416_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09968__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _07348_/A _07348_/B _07573_/A vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ _10469_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07281_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10290_ _10427_/A2 _10554_/C hold247/A vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ _08824_/A _08824_/B _08827_/A vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__a21o_2
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10502__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12931_ _13184_/A _12930_/B _12861_/X vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__a21o_1
X_12862_ hold302/X hold65/X vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__10502__B2 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11813_ _11813_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11058__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ hold104/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__or2_1
X_11744_ _11743_/B _11744_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__and2b_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08365__A _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__xnor2_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10626_ _10626_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10569__A1 _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ _13346_/CLK _13345_/D vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__dfxtp_1
X_10557_ _06749_/B _09228_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _10557_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07434__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ _10488_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__nand2_1
X_13276_ _13297_/CLK _13276_/D vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _06858_/A _12225_/X _12226_/Y vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__o21a_1
X_12158_ _12158_/A _12279_/C vssd1 vssd1 vccd1 vccd1 _12158_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13346_/CLK sky130_fd_sc_hd__clkbuf_8
X_12089_ _11935_/A _12010_/Y _12012_/B vssd1 vssd1 vccd1 vccd1 _12089_/Y sky130_fd_sc_hd__a21oi_1
X_11109_ _10886_/A _10999_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__11297__A2 _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ reg2_val[26] _06767_/A _06600_/Y _06649_/Y vssd1 vssd1 vccd1 vccd1 _07026_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06581_ instruction[11] _06575_/X _06580_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12246__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08275__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ _08320_/A _08378_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__or3_1
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _08251_/A _08251_/B vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07673__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ _07202_/A _07202_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07673__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09414__A2 _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _08178_/A _08178_/B _08249_/A vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07133_ _07135_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07133_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07064_ _07093_/A _07085_/D vssd1 vssd1 vccd1 vccd1 _07069_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11509__B1 _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07966_ _08007_/A _08007_/B vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__or2_1
X_06917_ instruction[19] _06575_/X _06916_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__or2_1
X_07897_ _07897_/A _07897_/B _07897_/C vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__and3_1
X_06848_ _06656_/X _06848_/B vssd1 vssd1 vccd1 vccd1 _06864_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06779_ reg1_val[4] _07097_/C vssd1 vssd1 vccd1 vccd1 _06780_/B sky130_fd_sc_hd__nand2_1
X_09567_ _09563_/X _09566_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13091__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _07018_/X wire8/X _09671_/A vssd1 vssd1 vccd1 vccd1 _09498_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_38_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08449_ _08566_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08861__B1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _11390_/A _11390_/B _11390_/C vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10411_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ _13130_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13131_/B sky130_fd_sc_hd__nand2_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07967__A2 _07060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07529__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13061_ hold111/X _13071_/A2 _13071_/B1 hold123/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold124/A sky130_fd_sc_hd__o221a_1
XANTENNA__07248__B _07248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _12012_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12154_/A sky130_fd_sc_hd__or2_2
X_10273_ _10175_/X _10570_/A _09148_/Y vssd1 vssd1 vccd1 vccd1 _10273_/Y sky130_fd_sc_hd__o21ai_1
X_12914_ _13145_/A _13146_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12845_ hold68/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12776_ hold154/X hold197/X hold193/X hold149/X vssd1 vssd1 vccd1 vccd1 _12778_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11987__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ _11988_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11658_ _11659_/B _11658_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11589_ _11589_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11592_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _10609_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08604__B1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07407__B2 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07407__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ _13334_/CLK hold113/X vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12951__A2 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _13364_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09580__A1 _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _09668_/A _07820_/B vssd1 vssd1 vccd1 vccd1 _07821_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07174__A _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _07808_/A _07750_/Y _07746_/Y vssd1 vssd1 vccd1 vccd1 _07765_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__10478__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _11446_/A reg1_val[17] vssd1 vssd1 vccd1 vccd1 _06704_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07682_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _07682_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06633_ _06978_/A reg1_val[25] vssd1 vssd1 vccd1 vccd1 _12115_/S sky130_fd_sc_hd__and2b_1
X_09421_ _13338_/Q _10158_/A2 hold265/A vssd1 vssd1 vccd1 vccd1 _09421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06564_ _06564_/A vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__inv_2
XFILLER_0_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _09353_/A _09353_/B vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08303_/Y sky130_fd_sc_hd__nand2b_1
X_09283_ _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09285_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08843__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09829__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ _08298_/A _08298_/B _08230_/Y vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__13195__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ _08167_/B _08167_/A vssd1 vssd1 vccd1 vccd1 _08165_/Y sky130_fd_sc_hd__nand2b_1
X_07116_ _11900_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07116_/Y sky130_fd_sc_hd__nor2_1
X_08096_ _09403_/S _08096_/B vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__nor2_1
X_07047_ _09668_/A _07053_/B vssd1 vssd1 vccd1 vccd1 _07048_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13086__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__B _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08998_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _08999_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07582__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _09795_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07950_/B sky130_fd_sc_hd__xnor2_1
X_10960_ _10959_/A _10959_/B _10959_/C vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout50_A _07059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _10406_/A _10890_/X _10889_/X vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__a21o_1
X_09619_ _09619_/A _09619_/B _09619_/C vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__and3_1
XFILLER_0_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12629_/A _12626_/Y _12628_/B vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12561_ _12574_/B _12575_/B _12574_/A vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10338__B1_N _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12492_ _12657_/B _12492_/B vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09739__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11512_ _11512_/A _11512_/B vssd1 vssd1 vccd1 vccd1 _11512_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__13186__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11443_ _09243_/B _11434_/X _11437_/X _11442_/X vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11374_ _11375_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__and2_1
X_13113_ hold313/X _13222_/A2 _13112_/X _12781_/A vssd1 vssd1 vccd1 vccd1 _13114_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _11296_/B _10325_/B vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10256_ _10256_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10258_/B sky130_fd_sc_hd__xor2_4
X_13044_ _07248_/B _13052_/A2 hold153/X vssd1 vssd1 vccd1 vccd1 _13320_/D sky130_fd_sc_hd__a21boi_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06610__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _11568_/A fanout31/X fanout29/X _07968_/B vssd1 vssd1 vccd1 vccd1 _10188_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12828_ _11749_/A _12842_/A2 hold66/X _13187_/A vssd1 vssd1 vccd1 vccd1 hold67/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12059__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09078__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A _12759_/B _12759_/C vssd1 vssd1 vccd1 vccd1 _12760_/B sky130_fd_sc_hd__and3_2
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07169__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08921_ _09544_/A _10129_/A vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08852_ _08852_/A _08852_/B vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08356__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _07803_/A _07803_/B vssd1 vssd1 vccd1 vccd1 _07858_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11350__A1_N _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ _08780_/A _08780_/B _11945_/A _11863_/B vssd1 vssd1 vccd1 vccd1 _08791_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__07316__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07794_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07632__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__xnor2_2
X_06616_ instruction[40] _06657_/B vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__and2_4
X_09404_ _09402_/X _09403_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__mux2_1
X_07596_ fanout64/X _08633_/B _09300_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _07597_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08816__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ fanout37/X _10326_/A _07218_/Y _07539_/B vssd1 vssd1 vccd1 vccd1 _09267_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08292__A1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13168__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08217_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08292__B2 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _09195_/X _09196_/X _09396_/S vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09241__B1 _09239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08148_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08079_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11103_/A sky130_fd_sc_hd__xor2_1
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__xor2_4
XANTENNA_fanout98_A _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _09301_/A _09941_/B _09942_/Y vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__o21ai_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__S _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _11992_/A _11992_/B vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__and2_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A3 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ fanout74/X fanout12/X fanout6/X _07249_/Y vssd1 vssd1 vccd1 vccd1 _10944_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11064__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10874_ _10874_/A _10874_/B vssd1 vssd1 vccd1 vccd1 _10876_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12613_ _12613_/A _12613_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12544_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12545_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10614__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__A _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08283__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12475_ _12481_/B _12475_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XFILLER_0_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11426_ _11781_/S _11426_/B vssd1 vssd1 vccd1 vccd1 _11426_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_6 reg1_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11357_ _11259_/A _11809_/C _11451_/A _12347_/B vssd1 vssd1 vccd1 vccd1 _11357_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10308_ curr_PC[7] _10438_/C _12490_/S vssd1 vssd1 vccd1 vccd1 _10308_/Y sky130_fd_sc_hd__a21oi_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11288_ _11289_/B _11288_/B vssd1 vssd1 vccd1 vccd1 _11290_/A sky130_fd_sc_hd__and2b_1
X_13027_ hold157/X _13055_/A2 _13053_/B1 hold176/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold177/A sky130_fd_sc_hd__o221a_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _10086_/A _10372_/A _10239_/C vssd1 vssd1 vccd1 vccd1 _10372_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__B1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13095__B2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__A1 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _07548_/B _07548_/A vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__and2b_1
X_07381_ _07197_/Y _08096_/B fanout24/X _08551_/A2 vssd1 vssd1 vccd1 vccd1 _07382_/B
+ sky130_fd_sc_hd__o22a_1
X_09120_ _09120_/A _09120_/B vssd1 vssd1 vccd1 vccd1 _09123_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _09051_/A _09051_/B vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _08594_/A2 _08354_/A2 _10585_/B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08003_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11030__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout100_A _07068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__A _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09953_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09884_ _10427_/A2 _10153_/C hold261/A vssd1 vssd1 vccd1 vccd1 _09884_/Y sky130_fd_sc_hd__a21oi_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08905_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07537__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A2 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ fanout58/X _07048_/Y _09648_/A fanout56/X vssd1 vssd1 vccd1 vccd1 _08836_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07001__A2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _08758_/B _08758_/C _08687_/B _08758_/A vssd1 vssd1 vccd1 vccd1 _08767_/C
+ sky130_fd_sc_hd__a211o_1
X_07717_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07717_/X sky130_fd_sc_hd__or2_1
XANTENNA__11636__A2 _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ _08705_/A _08705_/B _08803_/A _08695_/X vssd1 vssd1 vccd1 vccd1 _08799_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ _07351_/A _07351_/B _07340_/X vssd1 vssd1 vccd1 vccd1 _07650_/B sky130_fd_sc_hd__a21oi_4
X_07579_ _12193_/A _07346_/B _11813_/A vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11612__A _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09318_ _09318_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09320_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09289__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__A2 _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06706__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _10590_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout13_A _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__A _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _09249_/A _09249_/B vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__and2_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _12131_/A _07581_/A wire8/X _12259_/X vssd1 vssd1 vccd1 vccd1 _12315_/A sky130_fd_sc_hd__a31o_1
X_11211_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11318_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_121_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12191_ _12404_/B _12191_/B vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09765__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11142_ _11135_/Y _11136_/X _11140_/Y _11141_/X vssd1 vssd1 vccd1 vccd1 _11142_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10375__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__A _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10780__C1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11074_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11324__A1 _10406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07528__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _06774_/X _09886_/B _10023_/X vssd1 vssd1 vccd1 vccd1 _10024_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10898__A _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__A1 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ _11975_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09150__C1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10926_ curr_PC[11] curr_PC[12] _10926_/C vssd1 vssd1 vccd1 vccd1 _11149_/C sky130_fd_sc_hd__and3_2
X_10857_ _10982_/B _10857_/B vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12618__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10788_/A vssd1 vssd1 vccd1 vccd1 _10788_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _12685_/B _12527_/B vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ _12467_/A _12458_/B vssd1 vssd1 vccd1 vccd1 _12460_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11409_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11411_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11563__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B2 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ hold263/A _12347_/B _12387_/X _11242_/A vssd1 vssd1 vccd1 vccd1 _12390_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09508__A1 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06950_ _07146_/A _10286_/S _09725_/S _12785_/A vssd1 vssd1 vccd1 vccd1 _06950_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__09508__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06881_ _06765_/A _06765_/B _06774_/X _09886_/A vssd1 vssd1 vccd1 vccd1 _06883_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _09301_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08620_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08278__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _06875_/A _08551_/A2 _08551_/B1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08552_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07502_ _07503_/A _07503_/B vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__nand2_1
X_08482_ _08462_/A _08462_/B _08481_/Y vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07910__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ _07436_/A _07436_/B vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _09467_/A fanout9/A fanout5/X _09324_/A vssd1 vssd1 vccd1 vccd1 _09104_/B
+ sky130_fd_sc_hd__o22a_1
X_07364_ _10230_/A _07364_/B vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07295_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07353_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ _07659_/X _08913_/X _08914_/X vssd1 vssd1 vccd1 vccd1 _09034_/Y sky130_fd_sc_hd__a21oi_1
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__xor2_2
X_09867_ _12420_/A _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _09867_/Y sky130_fd_sc_hd__a21oi_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _11169_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08188__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__and2_1
XANTENNA__12806__A1 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _08749_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__and2_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11760_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07289__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _11813_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07820__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11690_/A _11808_/C _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12438__A _12619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13231__B2 _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _10643_/B _10643_/A vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08238__A1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__B2 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ _11083_/A _07347_/B fanout15/X _10966_/A vssd1 vssd1 vccd1 vccd1 _10574_/B
+ sky130_fd_sc_hd__o22a_1
X_13361_ _13363_/CLK _13361_/D vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dfxtp_1
X_13292_ _13352_/CLK _13292_/D vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__dfxtp_1
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__and2_1
XANTENNA__07461__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12243_ _06628_/B _09228_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10348__A2 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _12175_/A2 _12239_/B hold329/A vssd1 vssd1 vccd1 vccd1 _12174_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10405__B _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _11125_/A curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__or2_1
X_11056_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11057_/B sky130_fd_sc_hd__or2_1
XANTENNA__09482__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _12415_/A _06810_/Y _10006_/Y vssd1 vssd1 vccd1 vccd1 _10008_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08174__B1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08098__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11958_ _11958_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11889_ _11889_/A1 _11861_/X _11862_/Y _11888_/X vssd1 vssd1 vccd1 vccd1 _11889_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10908_/A _10908_/B _10908_/C vssd1 vssd1 vccd1 vccd1 _10910_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13222__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12430__C1 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12981__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ _10234_/A _07080_/B vssd1 vssd1 vccd1 vccd1 _07427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 _07264_/X vssd1 vssd1 vccd1 vccd1 _08551_/B1 sky130_fd_sc_hd__buf_6
Xfanout129 _07100_/X vssd1 vssd1 vccd1 vccd1 _08553_/A2 sky130_fd_sc_hd__clkbuf_8
X_07982_ _08043_/A _08043_/B _07961_/X vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__a21o_1
X_06933_ instruction[24] instruction[7] is_load _06767_/B _06932_/X vssd1 vssd1 vccd1
+ vccd1 _06934_/B sky130_fd_sc_hd__a32o_2
X_09721_ _09717_/X _09720_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _09721_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07905__A _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06864_ instruction[6] _06864_/B _06864_/C _06863_/X vssd1 vssd1 vccd1 vccd1 _06864_/X
+ sky130_fd_sc_hd__or4b_1
X_09652_ _09651_/B _09651_/C _09651_/A vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__a21oi_1
X_09583_ _10427_/A2 _09582_/X hold325/A vssd1 vssd1 vccd1 vccd1 _09583_/Y sky130_fd_sc_hd__a21oi_1
X_06795_ _06799_/A _06801_/B1 _12627_/B _06794_/X vssd1 vssd1 vccd1 vccd1 _09725_/S
+ sky130_fd_sc_hd__a31oi_4
X_08603_ _08611_/A _08611_/B vssd1 vssd1 vccd1 vccd1 _08603_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout265_A _06591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ _08556_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08465_ _08556_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07140__B2 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__A1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13213__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07416_ _07388_/Y _07416_/B vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__and2b_1
X_08396_ _08396_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08426_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09968__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__B2 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07347_ _12785_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07278_ _10469_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07282_/A sky130_fd_sc_hd__nand2_1
X_09017_ _08898_/A _08898_/B _08897_/A vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06703__B _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10750__A2 _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09499__A3 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ _12861_/X _12930_/B vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10502__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ hold77/X hold299/X vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _12202_/A fanout22/X fanout14/X _12059_/A vssd1 vssd1 vccd1 vccd1 _11813_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _07146_/Y _13078_/B2 hold49/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13245_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11463__B1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11743_ _11744_/B _11743_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__and2b_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11674_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13204__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10625_ _10625_/A _10625_/B vssd1 vssd1 vccd1 vccd1 _10626_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09477__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13344_ _13344_/CLK _13344_/D vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__dfxtp_1
X_10556_ hold213/A _11863_/A _10672_/B _12433_/A1 vssd1 vssd1 vccd1 vccd1 _10556_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07434__A2 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _10488_/A _10488_/B vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__or2_1
X_13275_ _13297_/CLK _13275_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
X_12226_ _06858_/A _12225_/X _11612_/A vssd1 vssd1 vccd1 vccd1 _12226_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12157_ _12270_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12279_/C sky130_fd_sc_hd__xor2_2
XANTENNA__07198__A1 _07193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__or2_2
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12088_/Y sky130_fd_sc_hd__nor2_1
X_11039_ curr_PC[13] _11149_/C _12490_/S vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09940__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ instruction[18] _06922_/B vssd1 vssd1 vccd1 vccd1 _06580_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09647__B1 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07673__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07201_ _07202_/A _07201_/B vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__xor2_4
X_08181_ _08248_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07132_ reg1_val[24] _07229_/B _07147_/B reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07135_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10326__A _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ reg1_val[6] reg1_val[7] _07063_/C _07063_/D vssd1 vssd1 vccd1 vccd1 _07085_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12182__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12182__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12541__A _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _08556_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _08007_/B sky130_fd_sc_hd__xnor2_1
X_06916_ instruction[26] _06922_/B vssd1 vssd1 vccd1 vccd1 _06916_/X sky130_fd_sc_hd__or2_1
XANTENNA__11157__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__and2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__nand2_1
X_07896_ _09301_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _07897_/C sky130_fd_sc_hd__xnor2_1
X_06847_ _06684_/Y _06840_/Y _06845_/X _11951_/A _06846_/Y vssd1 vssd1 vccd1 vccd1
+ _06848_/B sky130_fd_sc_hd__o221ai_4
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06778_ reg1_val[4] _07097_/C vssd1 vssd1 vccd1 vccd1 _06780_/A sky130_fd_sc_hd__or2_1
X_09566_ _09564_/X _09565_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _09566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09497_ _09669_/A _09497_/B vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08517_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__and2_1
XFILLER_0_108_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08448_ _06875_/A _10067_/A1 _08926_/B1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08449_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08861__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08861__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _11776_/A _08721_/A _08721_/B _12029_/A vssd1 vssd1 vccd1 vccd1 _10411_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ _08410_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__or2_1
X_11390_ _11390_/A _11390_/B _11390_/C vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__and3_1
XFILLER_0_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06714__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__nor2_2
X_13060_ _07108_/Y _13078_/B2 hold112/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__o21a_1
X_10272_ _10650_/B _10272_/B vssd1 vssd1 vccd1 vccd1 _10570_/A sky130_fd_sc_hd__xor2_4
X_12011_ _12011_/A _12011_/B _12011_/C vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__and3_1
X_12913_ hold53/X hold319/A vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11133__C1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12844_ _07593_/Y _13072_/A2 hold130/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold131/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09629__B1 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ hold197/X hold193/X hold149/X vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__nand3_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11436__B1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07280__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11726_ fanout57/X fanout9/X fanout4/X _11837_/A vssd1 vssd1 vccd1 vccd1 _11727_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11987__B2 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11657_ _12068_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13221__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _11589_/B _11589_/A vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__nand2b_1
X_10608_ _10608_/A _10608_/B _10608_/C vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__and3_1
XANTENNA__06624__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07407__A2 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13327_ _13334_/CLK _13327_/D vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10539_ _10442_/X _10537_/Y _10538_/Y vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09935__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ _13363_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13189_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__xnor2_1
X_12209_ _12267_/B _12209_/B vssd1 vssd1 vccd1 vccd1 _12212_/C sky130_fd_sc_hd__nor2_1
X_07750_ _07808_/B vssd1 vssd1 vccd1 vccd1 _07750_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10478__A1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ reg2_val[17] _06712_/B _06707_/B1 _06700_/Y vssd1 vssd1 vccd1 vccd1 _11446_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09670__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10478__B2 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _09668_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07685_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ hold9/A instruction[7] vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__and2_1
X_06632_ reg2_val[25] _06712_/B _06707_/B1 _06631_/Y vssd1 vssd1 vccd1 vccd1 _06978_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06563_ hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _09351_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _09353_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08302_ _08302_/A _08302_/B vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _09077_/A _09076_/Y _09072_/Y vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _08624_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08298_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08843__A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _08164_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ _08605_/B _08605_/C vssd1 vssd1 vccd1 vccd1 _07115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _08094_/A _08142_/A _08100_/A vssd1 vssd1 vccd1 vccd1 _08095_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07046_ _09668_/A _07053_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08359__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08997_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _08997_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07582__A1 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__B2 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _08591_/B1 _08096_/B fanout24/X _08619_/B1 vssd1 vssd1 vccd1 vccd1 _07949_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08531__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07881_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10890_/A _11112_/A vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__and2_1
X_09618_ _09619_/A _09619_/B _09619_/C vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__a21oi_1
X_09549_ _10128_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _10310_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11969__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _12547_/B _12552_/B _12610_/A vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _12657_/B _12492_/B vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__nand2_1
X_11511_ _11863_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11512_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11442_ _12175_/C1 _11439_/Y _11441_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1 _11442_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11373_ _11900_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11375_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12394__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13112_ hold309/X _13111_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__mux2_1
X_10324_ _10589_/A fanout9/A fanout5/X _10490_/A vssd1 vssd1 vccd1 vccd1 _10325_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10255_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__xnor2_4
X_13043_ hold134/X _13071_/A2 _13071_/B1 hold152/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold153/A sky130_fd_sc_hd__o221a_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _10186_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10189_/A sky130_fd_sc_hd__nor2_2
Xfanout290 reg1_val[15] vssd1 vssd1 vccd1 vccd1 _11231_/A sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ hold65/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09078__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ _12759_/B _12759_/C _12759_/A vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08834__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _11879_/A2 _11790_/B hold302/A vssd1 vssd1 vccd1 vccd1 _11709_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12689_ _12694_/B _12689_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
XFILLER_0_21_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__buf_6
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12803__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08920_ _08805_/B _08918_/X _08919_/X _08803_/X _08917_/X vssd1 vssd1 vccd1 vccd1
+ _10129_/A sky130_fd_sc_hd__o221a_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08851_ _08852_/A _08852_/B vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__or2_1
X_07802_ _08702_/A _08702_/B _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _07802_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08782_ _08786_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _11945_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07316__A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _07733_/A _07733_/B vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout178_A _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07664_/X sky130_fd_sc_hd__and2_1
X_06615_ _06613_/X _06615_/B vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09403_ _09185_/X _09211_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__mux2_1
X_07595_ _09669_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09334_ _09334_/A _09334_/B vssd1 vssd1 vccd1 vccd1 _09335_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08816__B2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A1 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _09930_/A _09265_/B vssd1 vssd1 vccd1 vccd1 _09269_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08292__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09196_ _09219_/A reg1_val[31] _09196_/S vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__mux2_1
X_08216_ _08216_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__or2_1
XANTENNA__12376__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ _08147_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08078_ _08078_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07029_ _07029_/A _07299_/B vssd1 vssd1 vccd1 vccd1 _07029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _09987_/A _09987_/B _09988_/Y vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__07004__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ _11992_/A _11992_/B vssd1 vssd1 vccd1 vccd1 _12073_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10942_ _10942_/A _10942_/B vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10873_ _10873_/A _10873_/B vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12605_/B _12607_/B _12605_/A vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10614__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08283__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11080__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _12474_/A _12474_/B _12474_/C vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ _06710_/Y _11331_/B _06711_/A vssd1 vssd1 vccd1 vccd1 _11426_/B sky130_fd_sc_hd__a21o_1
XANTENNA_7 reg1_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _12053_/A1 _11353_/X _11354_/Y _11355_/X vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__09485__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ curr_PC[7] _10438_/C vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__or2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11287_ _12068_/A _11287_/B vssd1 vssd1 vccd1 vccd1 _11288_/B sky130_fd_sc_hd__xor2_1
X_13026_ _09301_/A _13078_/B2 hold158/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__o21a_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _10237_/B _10237_/C _10237_/A vssd1 vssd1 vccd1 vccd1 _10239_/C sky130_fd_sc_hd__a21o_1
X_10169_ _10143_/Y _10144_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__A1 _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13095__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12842__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07380_ _07385_/B _07380_/B vssd1 vssd1 vccd1 vccd1 _07419_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11802__B1 _11777_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__A1 _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _09766_/A _09050_/B vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12358__A1 _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ _08057_/A _08057_/B vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11030__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12025__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _08902_/A _08902_/B _08904_/A vssd1 vssd1 vccd1 vccd1 _08903_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ hold230/A hold325/A hold285/A hold321/A vssd1 vssd1 vccd1 vccd1 _10153_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__B2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _10230_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__xnor2_2
X_08765_ _08260_/Y _08311_/Y _08263_/Y vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__a21o_1
X_07716_ _07734_/A _07714_/Y _07695_/Y vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11636__A3 _11809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ _07861_/X _08696_/B vssd1 vssd1 vccd1 vccd1 _08803_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _07650_/A sky130_fd_sc_hd__or2_2
XFILLER_0_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07578_ _07325_/A _07324_/Y _07320_/Y vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__a21o_1
X_09317_ _11168_/A _09317_/B vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06706__B _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__B _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _10286_/S _09250_/B vssd1 vssd1 vccd1 vccd1 _09249_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__B1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _11125_/A reg1_val[17] _09180_/S vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _11099_/A _11099_/B _11100_/Y vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__o21ai_2
X_12190_ _12309_/A fanout9/X fanout4/X _07302_/X vssd1 vssd1 vccd1 vccd1 _12191_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09765__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11141_ hold311/A _11879_/A2 _11139_/X _12393_/B1 vssd1 vssd1 vccd1 vccd1 _11141_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08973__B1 _06644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11072_ _11070_/X _11071_/Y _11169_/A vssd1 vssd1 vccd1 vccd1 _11074_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07528__A1 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _06774_/A _12395_/A1 _12394_/A1 _06772_/Y _10022_/X vssd1 vssd1 vccd1 vccd1
+ _10023_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07528__B2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A2 _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13077__A2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11974_ curr_PC[23] _12051_/C vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__and2_1
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10925_ _12029_/A _10895_/X _10896_/X _10924_/Y _10894_/Y vssd1 vssd1 vccd1 vccd1
+ _10925_/X sky130_fd_sc_hd__a311o_1
X_10856_ _10856_/A _10856_/B vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12618__B _12619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _09720_/X _09726_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10788_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12685_/B _12527_/B vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12457_ _12632_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07216__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__B _08831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ _12347_/B _12387_/X hold263/A vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08964__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _12171_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09508__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ hold251/X _12781_/A _12780_/B hold253/X vssd1 vssd1 vccd1 vccd1 hold254/A
+ sky130_fd_sc_hd__a22o_1
X_06880_ _10779_/A _10660_/A _06880_/C _06880_/D vssd1 vssd1 vccd1 vccd1 _06880_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__09154__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13068__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11079__B2 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08550_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08550_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07501_ _07689_/A _07689_/B _07497_/X vssd1 vssd1 vccd1 vccd1 _07503_/B sky130_fd_sc_hd__o21ai_1
X_08481_ _08489_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08481_/Y sky130_fd_sc_hd__nand2b_1
X_07432_ _11168_/A _07432_/B vssd1 vssd1 vccd1 vccd1 _07436_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _08980_/A _08980_/B _08978_/X vssd1 vssd1 vccd1 vccd1 _09106_/A sky130_fd_sc_hd__o21ai_2
X_07363_ fanout83/X _10463_/B2 _10228_/A fanout79/X vssd1 vssd1 vccd1 vccd1 _07364_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07294_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__and2_1
XANTENNA__07455__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout210_A _09101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _11155_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _09759_/X _09904_/B _09865_/Y vssd1 vssd1 vccd1 vccd1 _09866_/Y sky130_fd_sc_hd__a21oi_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _10937_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__xor2_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _11837_/A fanout77/X fanout73/X fanout61/X vssd1 vssd1 vccd1 vccd1 _09798_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12806__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08748_ _08748_/A _08748_/B _08748_/C vssd1 vssd1 vccd1 vccd1 _08749_/B sky130_fd_sc_hd__nand3_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08746_/A _08680_/C _08680_/D vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__nand3_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10710_ _07250_/X _07581_/A _07581_/B _07345_/X _07243_/X vssd1 vssd1 vccd1 vccd1
+ _10711_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07143__C1 _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A _11808_/C vssd1 vssd1 vccd1 vccd1 _11690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10643_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09435__B2 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08238__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _13363_/CLK _13360_/D vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ _10520_/A _10520_/B _10521_/Y vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _13352_/CLK _13291_/D vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__dfxtp_1
X_12311_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__nor2_1
X_12242_ _12242_/A _12242_/B vssd1 vssd1 vccd1 vccd1 _12242_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ hold269/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12239_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11124_ _11125_/A curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__nand2_1
X_11055_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11057_/A sky130_fd_sc_hd__nand2_1
X_10006_ _12415_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10006_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08174__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A2 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ _11957_/A _11957_/B vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ _10908_/A _10908_/B _10908_/C vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__and3_1
X_11888_ _11946_/A _11864_/Y _11869_/X _11887_/X vssd1 vssd1 vccd1 vccd1 _11888_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10839_ _07012_/Y fanout31/X fanout29/X _11917_/B vssd1 vssd1 vccd1 vccd1 _10840_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13222__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__A1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09938__A _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ _12509_/A _12509_/B _12509_/C vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_89_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07458__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout119 _10859_/A vssd1 vssd1 vccd1 vccd1 _08354_/A2 sky130_fd_sc_hd__buf_8
X_07981_ _07981_/A _07981_/B vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__xnor2_1
Xfanout108 _09114_/B1 vssd1 vssd1 vccd1 vccd1 _08926_/B1 sky130_fd_sc_hd__buf_6
X_06932_ instruction[40] _06593_/X _06930_/X _06931_/Y vssd1 vssd1 vccd1 vccd1 _06932_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12811__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _09718_/X _09719_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07193__A _07193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ _12772_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _06863_/X sky130_fd_sc_hd__or2_1
X_09651_ _09651_/A _09651_/B _09651_/C vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__and3_1
XANTENNA__06827__A_N _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ hold285/A hold321/A vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2_1
X_06794_ reg2_val[1] _06794_/B vssd1 vssd1 vccd1 vccd1 _06794_/X sky130_fd_sc_hd__and2_1
X_08602_ _08602_/A _08602_/B vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__nand2_1
X_08533_ _09403_/S _08533_/B vssd1 vssd1 vccd1 vccd1 _08534_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09114__B1 _09114_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08464_ _08507_/A2 _08619_/B1 _08591_/B1 _08533_/B vssd1 vssd1 vccd1 vccd1 _08465_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07140__A2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13213__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A1 _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07415_ _07415_/A _07415_/B vssd1 vssd1 vccd1 vccd1 _07416_/B sky130_fd_sc_hd__nand2_1
X_08395_ _08396_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__nor2_1
X_07346_ _12193_/A _07346_/B vssd1 vssd1 vccd1 vccd1 _07346_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07277_ _10469_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07281_/A sky130_fd_sc_hd__and2_1
XANTENNA__07368__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__B _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08928__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11618__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _09781_/A _09781_/B _09782_/X vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout73_A fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09849_/A _09849_/B vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__xnor2_2
X_12860_ hold316/A hold101/X vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__nand2b_1
X_11811_ _11758_/A _11757_/B _11757_/A vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__o21bai_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07831__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__A _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ hold48/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__or2_1
XANTENNA__11463__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ _11900_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__xnor2_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07667__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ _11723_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13204__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__C1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10624_ _10624_/A _10624_/B _10624_/C vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__and3_1
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13343_ _13343_/CLK _13343_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10555_ _11863_/A _10672_/B hold213/A vssd1 vssd1 vccd1 vccd1 _10555_/Y sky130_fd_sc_hd__a21oi_1
X_10486_ _10624_/A _10486_/B vssd1 vssd1 vccd1 vccd1 _10488_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07278__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ _13297_/CLK _13274_/D vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__dfxtp_2
X_12225_ _12415_/A _06867_/X _12224_/X vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__a21o_1
X_12156_ _12014_/A _11860_/B _12085_/A _12271_/B _12155_/X vssd1 vssd1 vccd1 vccd1
+ _12157_/B sky130_fd_sc_hd__o41a_1
XANTENNA__09592__B1 _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ _11107_/A _11107_/B _11107_/C vssd1 vssd1 vccd1 vccd1 _11108_/B sky130_fd_sc_hd__and3_1
XANTENNA__12631__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ _12087_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12087_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09344__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ curr_PC[13] _11149_/C vssd1 vssd1 vccd1 vccd1 _11038_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989_ hold255/A _13143_/B2 _13186_/A2 hold237/X vssd1 vssd1 vccd1 vccd1 hold238/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09647__A1 _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11454__B2 _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07200_ _07264_/A _06952_/C _07097_/C _07113_/A _07299_/B vssd1 vssd1 vccd1 vccd1
+ _07201_/B sky130_fd_sc_hd__o41ai_4
XANTENNA__09668__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08180_ _08573_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08248_/B sky130_fd_sc_hd__xnor2_1
X_07131_ reg1_val[24] _08868_/C _07229_/B reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07135_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10326__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07062_ _10231_/A _07062_/B vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07830__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08925__A3 _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07964_ _08533_/B _10585_/B2 _10067_/A1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _07965_/B
+ sky130_fd_sc_hd__o22a_1
X_06915_ instruction[18] _06575_/X _06914_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__10061__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__or2_1
X_07895_ _08633_/B fanout83/X fanout79/X _09300_/A vssd1 vssd1 vccd1 vccd1 _07896_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06846_ reg1_val[23] _07016_/A vssd1 vssd1 vccd1 vccd1 _06846_/Y sky130_fd_sc_hd__nand2_1
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06777_ _06799_/A _06801_/B1 _12642_/B _06775_/X vssd1 vssd1 vccd1 vccd1 _11237_/S
+ sky130_fd_sc_hd__a31oi_4
X_09565_ _09181_/X _09202_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09670_/A _09497_/B vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__nor2_1
X_08516_ _08545_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__xnor2_1
X_08447_ _08624_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08477_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08861__A2 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08378_ _08378_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10956__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06714__B _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07329_ _07128_/Y fanout41/X _07153_/Y _07402_/B vssd1 vssd1 vccd1 vccd1 _07330_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _10469_/A _10339_/Y _10338_/X vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ _09710_/B _10267_/X _10270_/Y vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08550__A_N _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _12012_/A vssd1 vssd1 vccd1 vccd1 _12010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10708__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11148__A1_N _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12912_ _13140_/A _13141_/A _13140_/B vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07888__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__A _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ hold129/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__or2_1
XANTENNA__09629__A1 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ hold193/X hold149/X vssd1 vssd1 vccd1 vccd1 _12774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11987__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ _12310_/A _11725_/B vssd1 vssd1 vccd1 vccd1 _11733_/A sky130_fd_sc_hd__xnor2_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _12143_/A fanout42/X fanout40/X _06978_/X vssd1 vssd1 vccd1 vccd1 _11657_/B
+ sky130_fd_sc_hd__a22o_1
Xfanout90 _09766_/A vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__buf_4
XFILLER_0_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12626__B _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11683_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__nand2_1
X_10607_ _10608_/A _10608_/B _10608_/C vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06624__B _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ _13334_/CLK hold119/X vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__dfxtp_1
X_10538_ _10442_/X _10537_/Y _11889_/A1 vssd1 vssd1 vccd1 vccd1 _10538_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13257_ _13363_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12208_/A _12208_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12209_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10469_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11372__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ _13188_/A _13188_/B vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__nand2_1
X_12139_ _12208_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11258__A _11258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13113__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ _06706_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _06700_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07343__A2 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ _08633_/B fanout50/X _09659_/B2 _09300_/A vssd1 vssd1 vccd1 vccd1 _07681_/B
+ sky130_fd_sc_hd__o22a_1
X_06631_ _06631_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _06631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06562_ hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _09350_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_75_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _09120_/A _09120_/B _09116_/X vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__a21o_1
X_08232_ _08641_/A2 _08354_/A2 fanout71/X _08649_/B vssd1 vssd1 vccd1 vccd1 _08233_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08843__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10337__A _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08159_/A _08159_/B _08156_/X vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07114_ _08605_/B _08605_/C vssd1 vssd1 vccd1 vccd1 _07114_/X sky130_fd_sc_hd__and2_4
X_08094_ _08094_/A _08142_/A vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__nor2_1
XANTENNA_wire8_A wire8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07045_ reg1_val[6] _07045_/B vssd1 vssd1 vccd1 vccd1 _07053_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08359__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08359__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11168__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__xnor2_2
X_07947_ _07947_/A _07947_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07582__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _09630_/A _07878_/B vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08531__A1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06829_ _07251_/A _11125_/A vssd1 vssd1 vccd1 vccd1 _06829_/X sky130_fd_sc_hd__and2b_1
X_09617_ _09617_/A _09617_/B vssd1 vssd1 vccd1 vccd1 _09619_/C sky130_fd_sc_hd__or2_1
XANTENNA__08531__B2 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09548_ _10129_/A _10129_/B _09546_/X _09547_/X vssd1 vssd1 vccd1 vccd1 _09549_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_93_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout36_A fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07098__A1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _12178_/A2 _11542_/A _11808_/B _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11510_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout2_A fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ reg1_val[8] curr_PC[8] _12490_/S vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ hold216/A _11441_/B vssd1 vssd1 vccd1 vccd1 _11441_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09101__A _09101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ _12202_/B fanout46/X fanout44/X _12202_/A vssd1 vssd1 vccd1 vccd1 _11373_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _13111_/A _13111_/B vssd1 vssd1 vccd1 vccd1 _13111_/Y sky130_fd_sc_hd__xnor2_1
X_10323_ _10259_/A _10259_/B _10257_/X vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__A1 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _10253_/A _10253_/B _10255_/A vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__o21ai_1
X_13042_ _10942_/A _13078_/B2 hold135/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__o21a_1
X_10185_ _10185_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__nor2_1
Xfanout280 _13016_/A vssd1 vssd1 vccd1 vccd1 _13057_/C1 sky130_fd_sc_hd__buf_4
Xfanout291 reg1_val[14] vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12826_ _11734_/A _12842_/A2 hold87/X _13187_/A vssd1 vssd1 vccd1 vccd1 hold88/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09078__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12757_/A _12757_/B _12757_/C vssd1 vssd1 vccd1 vccd1 _12759_/C sky130_fd_sc_hd__or3_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11708_ hold275/A _11708_/B vssd1 vssd1 vccd1 vccd1 _11790_/B sky130_fd_sc_hd__or2_1
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ _12688_/A _12688_/B _12688_/C vssd1 vssd1 vccd1 vccd1 _12689_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11639_ fanout29/X wire8/X _11559_/A vssd1 vssd1 vccd1 vccd1 _11639_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _13324_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _13309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12790__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__B2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11345__B1 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _11168_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__xnor2_1
X_07801_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _07801_/Y sky130_fd_sc_hd__nand2_1
X_08781_ _08168_/X _08772_/B _08691_/X vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07316__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _07732_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__xnor2_2
X_06614_ reg1_val[28] _08971_/B vssd1 vssd1 vccd1 vccd1 _06615_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09402_ _09208_/X _09210_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _08605_/A _07301_/Y _07593_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _07595_/B
+ sky130_fd_sc_hd__a22o_1
X_09333_ _09334_/A _09334_/B vssd1 vssd1 vccd1 vccd1 _09333_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13142__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__A _11451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08277__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _09928_/A _07347_/B fanout15/X _09815_/A vssd1 vssd1 vccd1 vccd1 _09265_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _12621_/A reg1_val[30] _09196_/S vssd1 vssd1 vccd1 vccd1 _09195_/X sky130_fd_sc_hd__mux2_1
X_08215_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08216_/B sky130_fd_sc_hd__and2_1
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _08143_/A _08143_/B _08216_/A vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09241__A2 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _08106_/A _08106_/B vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07028_ _07050_/A _07028_/B _07028_/C vssd1 vssd1 vccd1 vccd1 _08971_/D sky130_fd_sc_hd__or3_4
XFILLER_0_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07004__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _08979_/A _08979_/B vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__xnor2_4
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ _12068_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__xnor2_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10941_ _11172_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10942_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12300__A2 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ _12611_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__nor2_2
X_10872_ _10870_/A _10870_/B _10873_/B vssd1 vssd1 vccd1 vccd1 _10872_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12457__A _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11361__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12542_ _12549_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12544_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10614__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13013__B1 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ _12474_/A _12474_/B _12474_/C vssd1 vssd1 vccd1 vccd1 _12481_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09766__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _11776_/A _08760_/A _08760_/B _12029_/A vssd1 vssd1 vccd1 vccd1 _11424_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12192__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ curr_PC[16] _11448_/C _12053_/A1 vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11286_ _06993_/Y fanout42/X fanout40/X _11749_/A vssd1 vssd1 vccd1 vccd1 _11287_/B
+ sky130_fd_sc_hd__a22o_1
X_10306_ _12029_/A _10275_/Y _10276_/X _10305_/X _10274_/Y vssd1 vssd1 vccd1 vccd1
+ _10306_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07286__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10237_/A _10237_/B _10237_/C vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11327__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ hold181/A _13055_/A2 _13053_/B1 hold157/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold158/A sky130_fd_sc_hd__o221a_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09435__A1_N _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _09155_/S _10146_/X _10152_/X _09882_/X _10167_/X vssd1 vssd1 vccd1 vccd1
+ _10168_/X sky130_fd_sc_hd__a221o_1
X_10099_ _11359_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09299__A2 _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ hold35/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__or2_1
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__B2 _11778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__C1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08000_ _08000_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08057_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10615__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08431__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09951_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__xnor2_4
X_08902_ _08902_/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__nor2_2
X_09882_ _11238_/S _06924_/Y _09222_/Y vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__a21o_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A2 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_A _07043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ fanout52/X _10463_/B2 _10228_/A fanout50/X vssd1 vssd1 vccd1 vccd1 _08834_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13137__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__A _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08759_/A _08759_/B _08763_/A _08763_/B _11511_/B vssd1 vssd1 vccd1 vccd1
+ _11692_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07715_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08695_ _07934_/B _08696_/B _07861_/X vssd1 vssd1 vccd1 vccd1 _08695_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _07160_/Y _07222_/B _07223_/X vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__12046__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__xnor2_4
X_09316_ fanout50/X fanout77/X fanout73/X _09659_/B2 vssd1 vssd1 vccd1 vccd1 _09317_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09725_/S _09250_/B _09246_/X vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__A1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__C _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07473__B2 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09178_ _09176_/X _09177_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08445_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08134_/A sky130_fd_sc_hd__xnor2_2
X_11140_ _11879_/A2 _11139_/X hold311/A vssd1 vssd1 vccd1 vccd1 _11140_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08973__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _11071_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _11071_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07528__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _09240_/X _10020_/X _10021_/Y _11446_/B _06811_/B vssd1 vssd1 vccd1 vccd1
+ _10022_/X sky130_fd_sc_hd__o32a_1
XANTENNA__08649__B _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A3 _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ curr_PC[23] _12051_/C vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__or2_1
XANTENNA__10296__B1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10924_ _09243_/B _10911_/X _10923_/X _10901_/X vssd1 vssd1 vccd1 vccd1 _10924_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07161__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _10856_/A _10856_/B vssd1 vssd1 vccd1 vccd1 _10982_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10048__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11796__B1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ reg1_val[13] curr_PC[13] _12525_/S vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__mux2_1
X_10786_ _10786_/A _11958_/A _10784_/X vssd1 vssd1 vccd1 vccd1 _10786_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12456_ _12632_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09496__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _11309_/A _11309_/B _11310_/Y vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ hold253/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__or2_1
XANTENNA__07216__A1 _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11338_ _11338_/A _11338_/B vssd1 vssd1 vccd1 vccd1 _11338_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08964__B2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13323_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11269_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__xnor2_1
X_13008_ _13134_/A hold252/X vssd1 vssd1 vccd1 vccd1 _13302_/D sky130_fd_sc_hd__and2_1
XFILLER_0_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11079__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07500_ _07500_/A _07500_/B vssd1 vssd1 vccd1 vccd1 _07689_/B sky130_fd_sc_hd__xnor2_2
X_08480_ _08491_/A _08491_/B _08474_/Y vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__12809__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09170__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ _10327_/B2 fanout77/X fanout73/X _10589_/A vssd1 vssd1 vccd1 vccd1 _07432_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06807__B _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _09101_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ _07291_/A _07291_/B _07399_/A vssd1 vssd1 vccd1 vccd1 _07295_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__xor2_2
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12036__S _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__B1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout203_A _06901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _07201_/X fanout9/A fanout5/X _07264_/X vssd1 vssd1 vccd1 vccd1 _09935_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11711__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09759_/X _09904_/B _09148_/Y vssd1 vssd1 vccd1 vccd1 _09865_/Y sky130_fd_sc_hd__o21ai_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _07114_/X _07402_/B fanout41/X _07146_/Y vssd1 vssd1 vccd1 vccd1 _08817_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09800_/A vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__inv_2
XANTENNA__07391__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ _08748_/B _08748_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__a21o_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07143__B1 _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08746_/C sky130_fd_sc_hd__nor2_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ fanout98/X fanout85/X fanout83/X _10466_/A vssd1 vssd1 vccd1 vccd1 _07630_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06717__B _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11778__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _10526_/A _10525_/B _10525_/A vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _13352_/CLK _13290_/D vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__A1_N _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ hold301/A _12349_/A _12296_/B _12393_/B1 vssd1 vssd1 vccd1 vccd1 _12242_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _12171_/A _12170_/Y _12171_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _12183_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12470__A _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _06879_/B _11121_/Y _11122_/Y vssd1 vssd1 vccd1 vccd1 _11123_/X sky130_fd_sc_hd__a21o_1
X_11054_ _11054_/A _11054_/B vssd1 vssd1 vccd1 vccd1 _11056_/B sky130_fd_sc_hd__xnor2_1
X_10005_ _06780_/A _09870_/B _06780_/B vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__08174__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__A3 _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _11872_/B _11874_/B _11872_/A vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10907_ _10785_/B _10785_/C _10785_/A vssd1 vssd1 vccd1 vccd1 _10908_/C sky130_fd_sc_hd__a21bo_1
X_11887_ _11878_/Y _11879_/X _11886_/X _11876_/X vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10838_ _11172_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12430__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _10769_/A _11003_/A vssd1 vssd1 vccd1 vccd1 _10769_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08634__A0 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _12509_/A _12509_/B _12509_/C vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12439_ _12619_/B _12439_/B vssd1 vssd1 vccd1 vccd1 _12440_/B sky130_fd_sc_hd__or2_1
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _09630_/A _07978_/B _08050_/A vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__o21ai_1
X_06931_ instruction[6] is_load vssd1 vssd1 vccd1 vccd1 _06931_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09165__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07474__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _10231_/A _09650_/B _09650_/C vssd1 vssd1 vccd1 vccd1 _09651_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06862_ _06849_/Y _06861_/Y _06943_/B vssd1 vssd1 vccd1 vccd1 _06864_/C sky130_fd_sc_hd__a21oi_1
X_08601_ _08601_/A _08601_/B vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__or2_1
X_09581_ _09223_/Y _09596_/B _09574_/X vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__a21boi_1
X_06793_ _06793_/A _09595_/A vssd1 vssd1 vccd1 vccd1 _06793_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__12249__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _08573_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08562_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09114__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08463_ _08463_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout153_A _06995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__and2_2
XFILLER_0_107_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09417__A2 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ _08394_/A _08394_/B vssd1 vssd1 vccd1 vccd1 _08396_/B sky130_fd_sc_hd__xnor2_2
X_07345_ _12193_/A _07346_/B vssd1 vssd1 vccd1 vccd1 _07345_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08625__B1 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ reg1_val[10] _07276_/B vssd1 vssd1 vccd1 vccd1 _07280_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__A1 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ _09015_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__and2_2
XANTENNA__08928__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07087__C _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B2 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _09917_/A _09917_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__xor2_1
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout66_A fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10014__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _09695_/A _09695_/B _09693_/Y vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__a21boi_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10432__A2_N _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _09631_/A _09631_/B _09627_/X vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__a21oi_1
X_11810_ _12020_/A _12020_/B _12280_/A vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__a21o_1
X_12790_ _07153_/Y _13078_/B2 hold47/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13244_/D
+ sky130_fd_sc_hd__o211a_1
X_11741_ fanout44/X fanout11/X fanout7/A fanout46/X vssd1 vssd1 vccd1 vccd1 _11742_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09104__A _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__A1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A2 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07667__B2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11672_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__and3_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10623_ _10624_/A _10624_/B _10624_/C vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ hold257/A hold247/A _10554_/C vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__or3_1
X_13342_ _13343_/CLK _13342_/D vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _13374_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
X_10485_ _10484_/B _10485_/B vssd1 vssd1 vccd1 vccd1 _10486_/B sky130_fd_sc_hd__nand2b_1
X_12224_ _12162_/A _12160_/X _12378_/S _06652_/Y vssd1 vssd1 vccd1 vccd1 _12224_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _12013_/X _12271_/B _12153_/Y vssd1 vssd1 vccd1 vccd1 _12155_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11809__A _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11107_/A _11107_/B _11107_/C vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12086_ _12086_/A _12215_/A vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09344__A1 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__B2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _12029_/A _11010_/Y _11011_/X _11036_/X _11009_/X vssd1 vssd1 vccd1 vccd1
+ _11037_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12988_ _13144_/A hold256/X vssd1 vssd1 vccd1 vccd1 _13292_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09647__A2 _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _11939_/A _12086_/A vssd1 vssd1 vccd1 vccd1 _11939_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11454__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09949__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _11125_/A _11231_/A _07121_/C _07123_/A _07229_/B vssd1 vssd1 vccd1 vccd1
+ _07147_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07061_ _08590_/B fanout52/X _09648_/A fanout50/X vssd1 vssd1 vccd1 vccd1 _07062_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07830__A1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__B2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07594__B1 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _08573_/A _07963_/B vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__xnor2_1
X_06914_ instruction[25] _06922_/B vssd1 vssd1 vccd1 vccd1 _06914_/X sky130_fd_sc_hd__or2_1
X_09702_ _09702_/A _09702_/B vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__xnor2_4
X_07894_ _08648_/A _07894_/B _07894_/C vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__or3_1
X_06845_ _11947_/A _06843_/X _06844_/Y vssd1 vssd1 vccd1 vccd1 _06845_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__nand2b_1
X_09564_ _09174_/X _09178_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06776_ _06799_/A _06801_/B1 _12642_/B _06775_/X vssd1 vssd1 vccd1 vccd1 _06776_/X
+ sky130_fd_sc_hd__a31o_1
X_08515_ _08515_/A _08515_/B vssd1 vssd1 vccd1 vccd1 _08542_/A sky130_fd_sc_hd__xnor2_1
X_09495_ _09668_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09497_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08446_ _08649_/B _08521_/A2 _08551_/A2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08447_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08377_ _08409_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08410_/A sky130_fd_sc_hd__or2_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07328_ _07328_/A _07328_/B vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10956__A1 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__B2 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ _07259_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__and2_1
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10270_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10708__B2 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__B _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08003__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__A1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ hold56/X hold277/X vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07888__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07888__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _07301_/Y _12842_/A2 hold115/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold116/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09629__A2 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
X_11724_ _12059_/A fanout22/X fanout14/X _11980_/A vssd1 vssd1 vccd1 vccd1 _11725_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__xor2_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout91 _07133_/X vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__buf_8
Xfanout80 _07242_/Y vssd1 vssd1 vccd1 vccd1 _11188_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__06905__B _06907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__or2_1
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _10606_/A _10694_/A vssd1 vssd1 vccd1 vccd1 _10608_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09801__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13325_ _13334_/CLK hold146/X vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10537_ _10767_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13256_ _13363_/CLK hold55/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
X_10468_ _10468_/A _10468_/B _10468_/C vssd1 vssd1 vccd1 vccd1 _10469_/C sky130_fd_sc_hd__nand3_1
XANTENNA__06817__A_N _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _12208_/A _12208_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12642__B _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _13187_/A _13187_/B vssd1 vssd1 vccd1 vccd1 _13360_/D sky130_fd_sc_hd__and2_1
X_10399_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12138_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__and3_1
XANTENNA__11258__B _11258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _12070_/A _12070_/B vssd1 vssd1 vccd1 vccd1 _12138_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13113__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ instruction[35] _06657_/B vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__and2_4
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06561_ hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09280_ _09082_/X _09280_/B vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__and2b_1
X_08300_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__or2_2
XFILLER_0_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12817__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08776_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07113_ _07113_/A _07113_/B vssd1 vssd1 vccd1 vccd1 _08605_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ _08141_/A _08141_/B vssd1 vssd1 vccd1 vccd1 _08142_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07044_ _07063_/C _07063_/D _07093_/A vssd1 vssd1 vccd1 vccd1 _07045_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__A2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__B1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ _07947_/B _07947_/A vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__and2b_1
X_07877_ _07128_/Y _07944_/B fanout28/X _08476_/A vssd1 vssd1 vccd1 vccd1 _07878_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08531__A2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ _11014_/A _06826_/Y _06827_/X vssd1 vssd1 vccd1 vccd1 _06828_/Y sky130_fd_sc_hd__o21bai_1
X_09616_ _09615_/B _09616_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__and2b_1
X_06759_ _06757_/Y _06759_/B vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__nand2b_2
X_09547_ _09547_/A _09547_/B _09858_/A _09996_/A vssd1 vssd1 vccd1 vccd1 _09547_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_19_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06725__B _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13334_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08429_ _08429_/A _08429_/B vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__xnor2_2
X_11440_ hold326/A _11528_/C _11529_/B vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09101__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11371_ _12068_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11051__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13110_ _13110_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13111_/B sky130_fd_sc_hd__nand2_1
X_10322_ _10262_/A _10262_/B _10260_/X vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11359__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ hold195/A _13071_/A2 _13071_/B1 hold134/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold135/A sky130_fd_sc_hd__o221a_1
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10255_/B sky130_fd_sc_hd__nor2_2
X_10184_ _10185_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__and2_1
Xfanout270 _06590_/X vssd1 vssd1 vccd1 vccd1 _06767_/A sky130_fd_sc_hd__clkbuf_8
Xfanout281 _13109_/A vssd1 vssd1 vccd1 vccd1 _13016_/A sky130_fd_sc_hd__clkbuf_4
Xfanout292 _09219_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ hold86/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__or2_1
XANTENNA__11822__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ _12773_/A _12756_/B vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12637__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ hold225/A _11529_/B _11794_/B _11706_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _11715_/C sky130_fd_sc_hd__a311o_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12688_/A _12688_/B _12688_/C vssd1 vssd1 vccd1 vccd1 _12694_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11638_ _11900_/A _11638_/B vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09786__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11569_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13323_/CLK _13308_/D vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__A2 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ hold184/X _12780_/C _13236_/A vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__o21a_1
XANTENNA__11345__B2 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__nand2_1
X_07800_ _07800_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09173__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _08702_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _07731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07662_ _07662_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__xor2_4
X_06613_ reg1_val[28] _08971_/B vssd1 vssd1 vccd1 vccd1 _06613_/X sky130_fd_sc_hd__and2_1
X_07593_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07593_/Y sky130_fd_sc_hd__nand2_4
X_09401_ _09399_/X _09400_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09401_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _09334_/A _09334_/B vssd1 vssd1 vccd1 vccd1 _09332_/X sky130_fd_sc_hd__or2_1
XANTENNA__08277__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09474__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__B _11451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _09280_/B _09088_/B _09099_/B _09100_/B _09100_/A vssd1 vssd1 vccd1 vccd1
+ _09279_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_118_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13022__A1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09194_ _09192_/X _09193_/X _09396_/S vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08214_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08216_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08624_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08106_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ _07050_/A _07028_/B _07028_/C vssd1 vssd1 vccd1 vccd1 _07300_/A sky130_fd_sc_hd__nor3_4
XANTENNA__10083__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _08979_/A _08979_/B vssd1 vssd1 vccd1 vccd1 _08978_/X sky130_fd_sc_hd__or2_1
XANTENNA__07392__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12836__A1 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _07995_/B _07995_/A vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10847__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ fanout33/X _12257_/A fanout13/X fanout35/X vssd1 vssd1 vccd1 vccd1 _10941_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12610_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__nor2_1
X_10871_ _10728_/A _10728_/B _10727_/A vssd1 vssd1 vccd1 vccd1 _10873_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _12696_/B _12541_/B vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__or2_1
XANTENNA__11272__B1 _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ _12481_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _12474_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11423_ _11776_/A _08760_/A _08760_/B vssd1 vssd1 vccd1 vccd1 _11423_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07779__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ curr_PC[16] _11448_/C vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11327__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _09226_/Y _10279_/X _10280_/Y _10304_/X vssd1 vssd1 vccd1 vccd1 _10305_/X
+ sky130_fd_sc_hd__a31o_1
X_10236_ _10235_/A _10235_/B _10235_/C vssd1 vssd1 vccd1 vccd1 _10237_/C sky130_fd_sc_hd__a21o_1
X_13024_ _06990_/B _12797_/B hold182/X vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__a21boi_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10167_ _12171_/A _12107_/B1 _10166_/Y _10161_/X _10155_/Y vssd1 vssd1 vccd1 vccd1
+ _10167_/X sky130_fd_sc_hd__a311o_1
X_10098_ _07968_/B fanout31/X fanout29/X _07077_/X vssd1 vssd1 vccd1 vccd1 _10099_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11552__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _07179_/X _12842_/A2 hold96/X _13134_/A vssd1 vssd1 vccd1 vccd1 hold97/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06646__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11263__B1 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__A3 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12739_ _12740_/A _12740_/B vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _09951_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08901_ _07627_/A _07627_/B _07625_/X vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__a21o_2
XANTENNA__11727__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _09878_/X _09880_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__mux2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ _08832_/A _08832_/B vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12818__A1 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__B _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _08763_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _11604_/C sky130_fd_sc_hd__nor2_1
XANTENNA__10829__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07714_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ _07861_/A _07931_/A _07861_/C vssd1 vssd1 vccd1 vccd1 _08696_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11462__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07645_ _07355_/A _07354_/B _07352_/Y vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07576_ _07576_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ _09315_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _09196_/X _09250_/B _09396_/S vssd1 vssd1 vccd1 vccd1 _09246_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__A2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09177_ reg1_val[13] reg1_val[18] _09180_/S vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _08551_/A2 _10227_/B1 _10463_/A1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 _08129_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _08059_/A _08059_/B vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__xnor2_4
X_11070_ _11070_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout96_A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ hold293/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10021_/Y sky130_fd_sc_hd__nor2_1
X_11972_ _11972_/A _11972_/B _11972_/C _11971_/X vssd1 vssd1 vccd1 vccd1 _11972_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_98_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10923_ _09223_/Y _10904_/Y _10922_/Y _09196_/S _10921_/X vssd1 vssd1 vccd1 vccd1
+ _10923_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07161__A1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ _10854_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10856_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13234__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__A1_N _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10048__B2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10048__A1 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12530_/B _12524_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XANTENNA__12993__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10785_ _10785_/A _10785_/B _10785_/C vssd1 vssd1 vccd1 vccd1 _10786_/A sky130_fd_sc_hd__and3_1
XANTENNA__08110__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ reg1_val[3] curr_PC[3] _12504_/S vssd1 vssd1 vccd1 vccd1 _12457_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__xnor2_2
X_12386_ _09434_/Y _12385_/Y _12421_/B vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09610__B1 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07297__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11337_ _11335_/Y _11337_/B vssd1 vssd1 vccd1 vccd1 _11338_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08964__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11268_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11397_/A sky130_fd_sc_hd__nor2_1
X_11199_ _11083_/A _11155_/A _11084_/A _11085_/Y vssd1 vssd1 vccd1 vccd1 _11200_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11547__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ hold242/X _12781_/A _13209_/A2 hold251/X vssd1 vssd1 vccd1 vccd1 hold252/A
+ sky130_fd_sc_hd__a22o_1
X_10219_ _10933_/A _10219_/B vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07430_ _10230_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07436_/A sky130_fd_sc_hd__xnor2_1
X_07361_ _07361_/A _07361_/B vssd1 vssd1 vccd1 vccd1 _07362_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09100_ _09100_/A _09100_/B vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12825__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__nor2_1
X_07292_ _07398_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07399_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07455__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__13002__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__B1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08404__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09904_/B sky130_fd_sc_hd__or2_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ _09827_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__xnor2_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07391__A1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__B2 _06973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07670__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ _08746_/A _08746_/B _08746_/C _08746_/D vssd1 vssd1 vccd1 vccd1 _08748_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11475__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A1 _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _08736_/A _08736_/B _08484_/X _08678_/B vssd1 vssd1 vccd1 vccd1 _08680_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07221_/A _07221_/B _07207_/A vssd1 vssd1 vccd1 vccd1 _07640_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12975__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07559_ _07328_/A _07328_/B _07326_/Y vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ _10570_/A _10570_/B _10406_/X _10537_/Y vssd1 vssd1 vccd1 vccd1 _11809_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ _09240_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09229_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12240_ _12349_/A _12296_/B hold301/A vssd1 vssd1 vccd1 vccd1 _12242_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _12171_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11950__B2 _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ _06879_/B _11121_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _11122_/Y sky130_fd_sc_hd__o21ai_1
X_11053_ fanout55/X fanout25/X _12257_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11054_/B
+ sky130_fd_sc_hd__o22a_1
X_10004_ _10315_/A _08715_/A _08715_/B _12029_/A vssd1 vssd1 vccd1 vccd1 _10004_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07906__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _11953_/X _11955_/B vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__or2_1
X_11886_ _11881_/Y _11882_/X _11885_/X vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10837_ fanout35/X _10466_/B _10466_/C fanout33/X _12202_/B vssd1 vssd1 vccd1 vccd1
+ _10838_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12430__A2 _06644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _10530_/Y _11003_/A _10766_/Y vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _12516_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _12509_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_89_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09300__A _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10699_ _11052_/A _10699_/B vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__xnor2_1
X_12438_ _12619_/B _12439_/B vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08398__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _12369_/A _12405_/A vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06930_ instruction[17] _09243_/B _09222_/B _06767_/A vssd1 vssd1 vccd1 vccd1 _06930_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10181__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _06850_/X _06860_/Y _12381_/A vssd1 vssd1 vccd1 vccd1 _06861_/Y sky130_fd_sc_hd__o21ai_1
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06581__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09580_ _12421_/B _09579_/Y _09243_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__a21o_1
X_06792_ reg1_val[2] _07152_/A vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__or2_2
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08531_ _08572_/A2 _08619_/B1 _08591_/B1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 _08532_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09114__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__xnor2_1
X_07413_ _07413_/A _07413_/B _07413_/C vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__or3_1
XFILLER_0_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout146_A _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08393_ _08393_/A vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__inv_2
X_07344_ reg1_val[28] _07344_/B vssd1 vssd1 vccd1 vccd1 _07346_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12957__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07275_ reg1_val[8] reg1_val[9] _07085_/D _07093_/A vssd1 vssd1 vccd1 vccd1 _07276_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_103_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10983__A2 _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__or2_1
XFILLER_0_103_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10196__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__A2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold197 hold202/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__buf_1
X_09916_ _10933_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09917_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09889__B1 _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09849_/A sky130_fd_sc_hd__xnor2_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09666_/A _09666_/B _09663_/A vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__o21a_1
XANTENNA_fanout59_A _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08729_ _08673_/B _08673_/C _08673_/A vssd1 vssd1 vccd1 vccd1 _08730_/B sky130_fd_sc_hd__a21o_1
X_11740_ _11740_/A _11740_/B vssd1 vssd1 vccd1 vccd1 _11744_/B sky130_fd_sc_hd__xnor2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__B _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07667__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__a21oi_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11345__A2_N _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ _10696_/B _10622_/B vssd1 vssd1 vccd1 vccd1 _10624_/C sky130_fd_sc_hd__or2_1
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10553_ _10550_/X _10552_/X _11958_/A vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__mux2_1
X_13341_ _13341_/CLK _13341_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _13375_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10485_/B _10484_/B vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ _12279_/D _12221_/X _12222_/Y vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10187__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12154_ _12154_/A _12324_/A vssd1 vssd1 vccd1 vccd1 _12271_/B sky130_fd_sc_hd__or2_1
XANTENNA__11809__B _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A2 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _11105_/A _11105_/B vssd1 vssd1 vccd1 vccd1 _11107_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_102_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12085_ _12085_/A _12154_/A vssd1 vssd1 vccd1 vccd1 _12215_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09344__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _12107_/B1 _11023_/X _11035_/X _11015_/X vssd1 vssd1 vccd1 vccd1 _11036_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12987_ hold216/X _13143_/B2 _13186_/A2 hold255/X vssd1 vssd1 vccd1 vccd1 hold256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07107__A1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11938_ _11770_/Y _12086_/A _11936_/Y vssd1 vssd1 vccd1 vccd1 _11938_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ _11947_/A _11867_/X _11868_/Y vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13061__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07060_ _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09965__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07830__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09176__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07594__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _09701_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09702_/B sky130_fd_sc_hd__xor2_4
X_07962_ _08572_/A2 _08354_/A2 fanout71/X _08594_/A2 vssd1 vssd1 vccd1 vccd1 _07963_/B
+ sky130_fd_sc_hd__o22a_1
X_06913_ instruction[15] _06913_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
X_07893_ _07894_/B _07894_/C _08648_/A vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__o21ai_1
X_06844_ reg1_val[22] _06994_/A vssd1 vssd1 vccd1 vccd1 _06844_/Y sky130_fd_sc_hd__nand2_1
X_09632_ _09473_/A _09472_/B _09470_/X vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09561_/X _09562_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06775_ reg2_val[4] _06794_/B vssd1 vssd1 vccd1 vccd1 _06775_/X sky130_fd_sc_hd__and2_1
X_08514_ _08514_/A _08514_/B _08514_/C vssd1 vssd1 vccd1 vccd1 _08675_/A sky130_fd_sc_hd__and3_1
XFILLER_0_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09494_ _09300_/A fanout13/X fanout11/X _06991_/Y vssd1 vssd1 vccd1 vccd1 _09495_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08451_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06564__A _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08376_ _08556_/A _08376_/B vssd1 vssd1 vccd1 vccd1 _08409_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11602__B1 _11809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07327_ _07373_/A _07327_/B vssd1 vssd1 vccd1 vccd1 _07328_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10956__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09271__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07258_ _07259_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07611_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07189_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__and2_4
XANTENNA__10708__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11645__A _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _13135_/A _13136_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07888__A2 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ hold114/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09115__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12772_ _12772_/A _12772_/B vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08954__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__or2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11654_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11748_/A sky130_fd_sc_hd__and2b_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout92 _12193_/A vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__buf_8
Xfanout81 fanout82/X vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__buf_6
XFILLER_0_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout70 _07572_/Y vssd1 vssd1 vccd1 vccd1 _09930_/A sky130_fd_sc_hd__buf_4
X_10605_ _10735_/A _07282_/B fanout7/X _10604_/X vssd1 vssd1 vccd1 vccd1 _10694_/A
+ sky130_fd_sc_hd__o31a_2
XANTENNA__12397__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11585_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09785__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ _13324_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 _13324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _09998_/X _10534_/Y _10535_/Y _10532_/Y vssd1 vssd1 vccd1 vccd1 _10537_/B
+ sky130_fd_sc_hd__o211a_2
X_13255_ _13352_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
X_10467_ _10468_/B _10468_/C _10468_/A vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__a21o_1
X_12206_ _12206_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12208_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07025__B1 _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13186_ hold316/X _13186_/A2 _13185_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 _13187_/B
+ sky130_fd_sc_hd__a22o_1
X_10398_ _10398_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__xnor2_1
X_12137_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__a21oi_1
X_12068_ _12068_/A _12068_/B vssd1 vssd1 vccd1 vccd1 _12070_/B sky130_fd_sc_hd__xor2_1
X_11019_ reg1_val[12] curr_PC[12] _10908_/X vssd1 vssd1 vccd1 vccd1 _11020_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11274__B _11275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08230_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09253__B2 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07112_ _07299_/B _07113_/A _07097_/C vssd1 vssd1 vccd1 vccd1 _08605_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_43_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08092_ _08092_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08141_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07043_ reg1_val[7] _07043_/B vssd1 vssd1 vccd1 vccd1 _07043_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13010__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06831__B _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07567__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A1 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07945_ _09630_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07943__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07154__S _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _09616_/B _09615_/B vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__and2b_1
X_07876_ _10081_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__xnor2_1
X_06827_ _07255_/A reg1_val[13] vssd1 vssd1 vccd1 vccd1 _06827_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06758_ reg1_val[7] _07202_/A vssd1 vssd1 vccd1 vccd1 _06759_/B sky130_fd_sc_hd__nand2_1
X_09546_ _09370_/A _09370_/B _09545_/X vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__a21o_1
X_09477_ _10231_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__xnor2_1
X_06689_ reg1_val[19] _07058_/A vssd1 vssd1 vccd1 vccd1 _06690_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ _08428_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10929__A2 _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ _08649_/B _10067_/A1 _08926_/B1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08360_/B
+ sky130_fd_sc_hd__o22a_1
X_11370_ _11917_/B fanout42/X fanout40/X _06993_/Y vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11051__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11051__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12235__S _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ _09863_/C _10319_/X _10320_/X _10318_/Y vssd1 vssd1 vccd1 vccd1 _10406_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_33_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06741__B _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ _07235_/B _13052_/A2 hold196/X vssd1 vssd1 vccd1 vccd1 _13318_/D sky130_fd_sc_hd__a21boi_1
X_10252_ _10078_/A _10078_/B _10076_/Y vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__06766__C1 _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _11557_/A _10183_/B vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout260 _06564_/A vssd1 vssd1 vccd1 vccd1 _12781_/A sky130_fd_sc_hd__buf_4
Xfanout282 _13219_/A vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__buf_4
Xfanout271 _06908_/A vssd1 vssd1 vccd1 vccd1 _06799_/A sky130_fd_sc_hd__buf_8
XANTENNA__08507__B1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A0 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _09219_/A sky130_fd_sc_hd__buf_4
X_12824_ _11568_/A _12842_/A2 hold60/X _13144_/A vssd1 vssd1 vccd1 vccd1 hold61/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12067__B1 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11814__B1 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _12764_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__or2_1
XANTENNA__06916__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11706_ _11529_/B _11794_/B hold225/A vssd1 vssd1 vccd1 vccd1 _11706_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12694_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12688_/C sky130_fd_sc_hd__nand2_1
X_11637_ fanout44/X fanout13/X fanout11/X fanout46/X vssd1 vssd1 vccd1 vccd1 _11638_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11568_ _11568_/A _11917_/C vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09786__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10519_ _10394_/A _10394_/B _10392_/X vssd1 vssd1 vccd1 vccd1 _10520_/B sky130_fd_sc_hd__a21oi_2
X_13307_ _13323_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12790__A1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11499_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11501_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__S _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ hold1/X _12778_/B _13237_/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
X_13169_ _13187_/A hold296/X vssd1 vssd1 vccd1 vccd1 _13356_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07763__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _07800_/A _07800_/B _07664_/X vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07661_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _08702_/A sky130_fd_sc_hd__xnor2_4
X_06612_ _06610_/Y _06707_/B1 _06767_/A reg2_val[28] vssd1 vssd1 vccd1 vccd1 _08971_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_07592_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__and2_2
X_09400_ _09204_/X _09207_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09400_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09334_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09474__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ _09137_/A _09137_/B _09138_/Y vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__13022__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ reg1_val[2] reg1_val[29] _09560_/A vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__mux2_1
X_08213_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08213_/X sky130_fd_sc_hd__and2_1
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08649_/B fanout79/X fanout75/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08076_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07026_ _07029_/A _07026_/B _07026_/C vssd1 vssd1 vccd1 vccd1 _07028_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _09668_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08979_/B sky130_fd_sc_hd__xnor2_4
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12836__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07995_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10847__A1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B2 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _07930_/A _07930_/B _07930_/C vssd1 vssd1 vccd1 vccd1 _07931_/A sky130_fd_sc_hd__o21ai_1
X_10870_ _10870_/A _10870_/B vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12049__B1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09279_/A _09279_/B _09278_/A vssd1 vssd1 vccd1 vccd1 _09534_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06736__B _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12540_ _12696_/B _12541_/B vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__A2 _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ _12642_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12472_/B sky130_fd_sc_hd__or2_1
XFILLER_0_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12221__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ _11357_/X _11451_/B _11421_/Y vssd1 vssd1 vccd1 vccd1 _11422_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08976__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07779__A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _11326_/Y _11327_/X _11328_/Y _11329_/X _11352_/X vssd1 vssd1 vccd1 vccd1
+ _11353_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _12065_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__xor2_1
X_10304_ _09152_/Y _10282_/X _10288_/X _09882_/X _10303_/Y vssd1 vssd1 vccd1 vccd1
+ _10304_/X sky130_fd_sc_hd__a221o_1
X_10235_ _10235_/A _10235_/B _10235_/C vssd1 vssd1 vccd1 vccd1 _10237_/B sky130_fd_sc_hd__nand3_1
X_13023_ _13309_/Q _13055_/A2 _13053_/B1 hold181/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold182/A sky130_fd_sc_hd__o221a_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07400__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _10166_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10166_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10097_ _10933_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ hold95/X _12839_/B vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10449__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06659__A2_N _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ _10999_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__or2_2
XANTENNA__06646__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07467__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12738_ _12719_/B _12737_/X _12767_/B _07123_/A vssd1 vssd1 vccd1 vccd1 _12740_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ _12670_/A _12670_/C _12670_/B vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08431__A2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09880_ _09736_/X _10902_/B _10902_/A vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _07577_/A _07576_/B _07576_/A vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__xor2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08761_/B _08761_/C _08761_/A vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07942__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A1 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _07790_/A _07790_/B _07706_/X vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__a21oi_1
X_08693_ _08061_/X _08168_/X _08772_/B _08690_/Y _08692_/X vssd1 vssd1 vccd1 vccd1
+ _08705_/B sky130_fd_sc_hd__o311a_2
XANTENNA_fanout176_A _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07644_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ _07574_/A _07574_/C _07574_/B vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _11237_/S _09250_/B vssd1 vssd1 vccd1 vccd1 _09245_/X sky130_fd_sc_hd__or2_4
XFILLER_0_29_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07668__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09176_ reg1_val[12] reg1_val[19] _09180_/S vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _08109_/X _08204_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08127_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__11962__C1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _08164_/A _08164_/B _08001_/X vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__a21o_1
X_07009_ _07009_/A _07009_/B vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout89_A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ hold293/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__and2_1
X_11971_ _11971_/A _11971_/B _11971_/C vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__and3_1
XANTENNA__11653__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10296__A2 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _11131_/A _09727_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07161__A2 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10853_ _10854_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10048__A2 _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10785_/A _10785_/B _10785_/C vssd1 vssd1 vccd1 vccd1 _10784_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _12523_/A _12523_/B _12523_/C vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__nand3_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12484__A _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ _12460_/B _12454_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08949__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ reg1_val[30] _12421_/C vssd1 vssd1 vccd1 vccd1 _12385_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09610__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11267_ _11369_/A _11267_/B vssd1 vssd1 vccd1 vccd1 _11269_/B sky130_fd_sc_hd__nand2_1
X_13006_ _13134_/A hold243/X vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__and2_1
XANTENNA__10732__A _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ _11078_/A _11078_/B _11076_/X vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11181__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10218_ _07150_/Y _07243_/X _07250_/X _07155_/A vssd1 vssd1 vccd1 vccd1 _10219_/B
+ sky130_fd_sc_hd__a22o_1
X_10149_ _10147_/X _10148_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09677__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__B2 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__S _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13225__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07360_ _07428_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _07361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08872__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09179__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ _07291_/A _07291_/B vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__xnor2_1
X_09030_ _09030_/A _09030_/B vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12841__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__or2_1
XANTENNA__06718__A2 _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _10319_/A _09863_/B _09863_/C vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__and3_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _11456_/A fanout27/X fanout25/X fanout98/X vssd1 vssd1 vccd1 vccd1 _09795_/B
+ sky130_fd_sc_hd__o22a_1
X_08814_ _07814_/B _07197_/Y _07201_/X fanout45/X vssd1 vssd1 vccd1 vccd1 _08815_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07391__A2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ _08421_/Y _08486_/Y _08424_/X vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__11475__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A1 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _08673_/A _08673_/B _08673_/C _08734_/A _08674_/X vssd1 vssd1 vccd1 vccd1
+ _08736_/B sky130_fd_sc_hd__a41o_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07627_ _07627_/A _07627_/B vssd1 vssd1 vccd1 vccd1 _07642_/A sky130_fd_sc_hd__xor2_1
X_07558_ _07488_/A _07488_/B _07489_/Y vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10817__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07489_ _07490_/B _07490_/A vssd1 vssd1 vccd1 vccd1 _07489_/Y sky130_fd_sc_hd__nand2b_1
X_09228_ _09240_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09228_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _09157_/X _09158_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _12170_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12170_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07603__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _11781_/S _06828_/Y _11120_/Y vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__xnor2_1
X_10003_ _10315_/A _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _10003_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07906__A1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__B2 _09114_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11383__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11954_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06908__C _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ _09155_/S _10552_/X _10565_/Y _09222_/Y _11884_/X vssd1 vssd1 vccd1 vccd1
+ _11885_/X sky130_fd_sc_hd__a221o_1
X_10905_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__nand2_1
X_10836_ _10836_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _10767_/A _10888_/A vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10698_ fanout61/X fanout46/X fanout44/X _11645_/A vssd1 vssd1 vccd1 vccd1 _10699_/B
+ sky130_fd_sc_hd__o22a_1
X_12506_ _12666_/B _12506_/B vssd1 vssd1 vccd1 vccd1 _12507_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__B _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07842__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ _09219_/A curr_PC[0] _12525_/S vssd1 vssd1 vccd1 vccd1 _12439_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09727__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08398__A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__B2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12368_ _12368_/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12405_/B sky130_fd_sc_hd__or2_1
XANTENNA__12661__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11319_ _11317_/Y _11319_/B vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__nand2b_2
X_12299_ _06613_/X _12431_/A2 _09225_/X vssd1 vssd1 vccd1 vccd1 _12299_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11154__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _06851_/Y _06859_/X _06656_/A vssd1 vssd1 vccd1 vccd1 _06860_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10799__A2_N _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ reg1_val[2] _07152_/A vssd1 vssd1 vccd1 vccd1 _06793_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08530_ _08536_/B _08536_/A vssd1 vssd1 vccd1 vccd1 _08530_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07125__A2 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08461_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__xnor2_1
X_07412_ _07413_/A _07413_/B _07413_/C vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08392_ _08392_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08393_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07343_ _08868_/C _12756_/B _07229_/B vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07274_ _07647_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07295_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09015_/A sky130_fd_sc_hd__nand2_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10196__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__B2 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A1 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _07155_/A _10222_/A2 _07255_/Y _07151_/A vssd1 vssd1 vccd1 vccd1 _09916_/B
+ sky130_fd_sc_hd__a22o_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07681__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _09671_/A _06990_/B vssd1 vssd1 vccd1 vccd1 _06991_/A sky130_fd_sc_hd__or2_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09840_/A sky130_fd_sc_hd__xor2_4
X_08728_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _10657_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B1 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ _08650_/A _08653_/A _08659_/S vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__mux2_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11672_/C sky130_fd_sc_hd__xor2_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__and2_1
XANTENNA__06744__B _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ _13343_/CLK _13340_/D vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ _10145_/X _10551_/X _11237_/S vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _13375_/CLK hold131/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08017__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10483_ _12068_/A _10483_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__xor2_1
X_12222_ _12279_/D _12221_/X _09149_/X vssd1 vssd1 vccd1 vccd1 _12222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11384__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A1 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__B2 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11378__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _12012_/A _12082_/Y _12084_/B vssd1 vssd1 vccd1 vccd1 _12153_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11104_ _11105_/B _11105_/A vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ _12082_/Y _12084_/B vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__11136__B1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _09222_/Y _11022_/X _11034_/X _09155_/S _11033_/Y vssd1 vssd1 vccd1 vccd1
+ _11035_/X sky130_fd_sc_hd__a221o_1
X_12986_ _13144_/A hold217/X vssd1 vssd1 vccd1 vccd1 _13291_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11937_ _11937_/A _12014_/A vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__nor2_1
X_11868_ _11947_/A _11867_/X _09226_/Y vssd1 vssd1 vccd1 vccd1 _11868_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12656__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11799_ _09196_/S _10669_/X _10682_/Y _09223_/Y _11798_/X vssd1 vssd1 vccd1 vccd1
+ _11799_/X sky130_fd_sc_hd__o221a_1
X_10819_ _07236_/A fanout6/X _10942_/A vssd1 vssd1 vccd1 vccd1 _10819_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07815__B1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__A2 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _07951_/A _08046_/A _07981_/B vssd1 vssd1 vccd1 vccd1 _07961_/X sky130_fd_sc_hd__o21ba_1
X_06912_ instruction[14] _06913_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
X_09700_ _09701_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__and2_1
X_07892_ _07060_/A _07060_/B _08551_/B2 vssd1 vssd1 vccd1 vccd1 _07894_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09192__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06843_ _11782_/A _06842_/Y _06841_/Y vssd1 vssd1 vccd1 vccd1 _06843_/X sky130_fd_sc_hd__o21a_1
X_09631_ _09631_/A _09631_/B vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13008__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__B _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06774_ _06774_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _06774_/X sky130_fd_sc_hd__or2_1
X_09562_ _09166_/X _09171_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__mux2_1
X_08513_ _08515_/A _08515_/B vssd1 vssd1 vccd1 vccd1 _08514_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout256_A _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _09493_/A _09493_/B vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08444_ _08619_/B1 _10227_/B1 _10463_/A1 _09403_/S vssd1 vssd1 vccd1 vccd1 _08445_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _08533_/B _08553_/B1 _09468_/B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08376_/B
+ sky130_fd_sc_hd__o22a_1
X_07326_ _07373_/A _07327_/B vssd1 vssd1 vccd1 vccd1 _07326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07257_ _11168_/A _07257_/B vssd1 vssd1 vccd1 vccd1 _07259_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ reg1_val[19] _07208_/B _07188_/C vssd1 vssd1 vccd1 vccd1 _07192_/B sky130_fd_sc_hd__or3_2
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07034__B2 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11118__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10830__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11645__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _11359_/A _09829_/B vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__xnor2_2
X_12840_ _07031_/X _12842_/A2 hold72/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold73/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06739__B _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12768_/B _12770_/B _12766_/X vssd1 vssd1 vccd1 vccd1 _12772_/B sky130_fd_sc_hd__a21oi_1
X_11722_ _11542_/A _11808_/B _11809_/D _11808_/C _12347_/B vssd1 vssd1 vccd1 vccd1
+ _11774_/A sky130_fd_sc_hd__o41a_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _12065_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__xnor2_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout82 _07239_/X vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_8
X_10604_ _07284_/X wire8/X _10736_/A vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__a21o_1
Xfanout60 _06999_/X vssd1 vssd1 vccd1 vccd1 fanout60/X sky130_fd_sc_hd__buf_6
Xfanout71 _10966_/A vssd1 vssd1 vccd1 vccd1 fanout71/X sky130_fd_sc_hd__buf_8
XFILLER_0_37_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__xnor2_1
Xfanout93 _10937_/A vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__buf_8
XFILLER_0_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13323_ _13323_/CLK _13323_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08970__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12492__A _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10535_ _09374_/A _09374_/B _09996_/Y _10534_/A _10769_/A vssd1 vssd1 vccd1 vccd1
+ _10535_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_0_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _13350_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_10466_ _10466_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _10468_/C sky130_fd_sc_hd__or3_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13185_ hold299/X _13184_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07025__A1 _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12255_/B _12205_/B _12206_/B vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__and3_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ _12204_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12138_/C sky130_fd_sc_hd__nor2_1
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12306__C1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ fanout40/X _08857_/Y wire8/X fanout42/X vssd1 vssd1 vccd1 vccd1 _12068_/B
+ sky130_fd_sc_hd__a22o_1
X_11018_ _11018_/A _11018_/B vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06649__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12969_ hold257/A _13095_/B2 _13158_/A2 hold213/X vssd1 vssd1 vccd1 vccd1 hold214/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08289__B1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10096__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08160_/Y sky130_fd_sc_hd__nor2_1
X_07111_ _07116_/B _11823_/A vssd1 vssd1 vccd1 vccd1 _07111_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09253__A2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08091_ _10468_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08141_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07042_ reg1_val[6] _07063_/C _07063_/D _07093_/A vssd1 vssd1 vccd1 vccd1 _07043_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__07496__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07567__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _11813_/A _08993_/B vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09372__A1_N _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _08476_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06790__A3 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _09928_/A _08184_/B fanout32/X _09815_/A vssd1 vssd1 vccd1 vccd1 _07876_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ _06733_/Y _06824_/Y _06825_/X vssd1 vssd1 vccd1 vccd1 _06826_/Y sky130_fd_sc_hd__a21oi_1
X_09614_ _10937_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13172__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ reg1_val[7] _07202_/A vssd1 vssd1 vccd1 vccd1 _06757_/Y sky130_fd_sc_hd__nor2_1
X_09545_ _09145_/A _09145_/B _09370_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09545_/X
+ sky130_fd_sc_hd__o22a_1
X_06688_ _07058_/A reg1_val[19] vssd1 vssd1 vccd1 vccd1 _11626_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ fanout55/X _09648_/A _12257_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _09477_/B
+ sky130_fd_sc_hd__o22a_1
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10097__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08358_ _08361_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _08358_/X sky130_fd_sc_hd__or2_1
XANTENNA__11051__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _08594_/A2 _08521_/A2 _08551_/A2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08290_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07309_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07586_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _09042_/A _09042_/B _09858_/X _10319_/X vssd1 vssd1 vccd1 vccd1 _10320_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _10107_/A _10107_/B _10108_/Y vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__a21bo_2
X_10182_ fanout61/X fanout27/X fanout25/X _11645_/A vssd1 vssd1 vccd1 vccd1 _10183_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout250 _12421_/B vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__clkbuf_8
Xfanout283 _13219_/A vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__buf_4
Xfanout261 hold132/X vssd1 vssd1 vccd1 vccd1 _06564_/A sky130_fd_sc_hd__clkbuf_4
Xfanout272 _06589_/X vssd1 vssd1 vccd1 vccd1 _06908_/A sky130_fd_sc_hd__buf_4
XANTENNA__08507__B2 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__A1 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout294 instruction[7] vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__08965__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ hold59/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__or2_1
XANTENNA__12067__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12754_ reg1_val[28] _12773_/A vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__nor2_1
X_11705_ hold237/A _11705_/B vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__or2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ reg1_val[13] _12685_/B vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__or2_1
XFILLER_0_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11636_ _11542_/A _11808_/B _11809_/D _12347_/B vssd1 vssd1 vccd1 vccd1 _11690_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11567_/A _11567_/B vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10735__A _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _10518_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__xnor2_1
X_13306_ _13323_/CLK _13306_/D vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12790__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11498_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__nand2b_1
X_13237_ hold1/X _12780_/B hold198/A _12781_/A vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10449_ _11557_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10002__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ hold295/X _13186_/A2 _13167_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold296/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11566__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12118_/X _12119_/B _12119_/C vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__and3b_1
XANTENNA__12161__S _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ hold317/X _13222_/A2 _13098_/X _13108_/B2 vssd1 vssd1 vccd1 vccd1 hold318/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10305__A1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07660_ _07660_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _09035_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08875__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ reg2_val[28] _06794_/B _06707_/B1 _06610_/Y vssd1 vssd1 vccd1 vccd1 _06851_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_07591_ _07074_/B _07300_/A _07300_/B _08971_/A vssd1 vssd1 vccd1 vccd1 _07593_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09330_ _09330_/A _09330_/B vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09474__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _09142_/A _09142_/B _09140_/X vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_117_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13007__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08212_ _08212_/A _08212_/B vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ reg1_val[3] reg1_val[28] _09560_/A vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07237__A1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout121_A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _08143_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06842__B _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__A1 _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ _08566_/A _08074_/B vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07025_ _07026_/B _06967_/A _06967_/B _07026_/C _07029_/A vssd1 vssd1 vccd1 vccd1
+ _07025_/X sky130_fd_sc_hd__a41o_1
XANTENNA__10792__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09934__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ fanout67/X _09300_/A fanout55/X _08633_/B vssd1 vssd1 vccd1 vccd1 _08977_/B
+ sky130_fd_sc_hd__o22a_2
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07925_/A _07925_/B _07926_/X vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__a21o_2
XANTENNA__10847__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07173__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _07858_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07930_/C sky130_fd_sc_hd__xor2_1
X_06809_ reg1_val[4] _11237_/S vssd1 vssd1 vccd1 vccd1 _06809_/X sky130_fd_sc_hd__and2_1
X_07789_ _07789_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07791_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _09361_/A _09361_/B _09359_/Y vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout34_A _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _09459_/A _09459_/B vssd1 vssd1 vccd1 vccd1 _09526_/A sky130_fd_sc_hd__and2_2
XANTENNA__11272__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _12642_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__nand2_1
X_11421_ _11357_/X _11451_/B _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _11612_/A _11333_/Y _11340_/X _11351_/X vssd1 vssd1 vccd1 vccd1 _11352_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10232__B1 _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__B2 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _11238_/S _09243_/B _10302_/Y _10297_/X vssd1 vssd1 vccd1 vccd1 _10303_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_15_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11283_ _07012_/Y _07151_/A _07155_/A _11917_/B vssd1 vssd1 vccd1 vccd1 _11284_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11327__A3 _11451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _10234_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10235_/C sky130_fd_sc_hd__xor2_2
X_13022_ _09671_/A _12797_/B hold19/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11386__A _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _10163_/Y _10165_/B vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07400__B2 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _07151_/A _07250_/X _07255_/Y _07155_/A vssd1 vssd1 vccd1 vccd1 _10097_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12806_ _07212_/X _12842_/A2 hold33/X _13134_/A vssd1 vssd1 vccd1 vccd1 hold34/A
+ sky130_fd_sc_hd__o211a_1
X_10998_ _10998_/A _10998_/B _10998_/C vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__and3_1
XFILLER_0_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__B2 _06973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__A1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ _12737_/A _12737_/B _12737_/C _12737_/D vssd1 vssd1 vccd1 vccd1 _12737_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__06943__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _12664_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12670_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _11238_/S _10922_/Y _11618_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _11630_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07219__B2 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A1 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ _12585_/B _12593_/B _12616_/A vssd1 vssd1 vccd1 vccd1 _12600_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11296__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08830_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08830_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06745__A3 _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B _08761_/C vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__and3_1
XANTENNA__10829__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _07712_/A _07712_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__xor2_1
X_08692_ _08161_/Y _08165_/Y _08166_/X _08786_/A _08790_/A vssd1 vssd1 vccd1 vccd1
+ _08692_/X sky130_fd_sc_hd__a2111o_1
XANTENNA__12839__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07643_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__nor2_2
XANTENNA__13016__A _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__or2_1
X_07574_ _07574_/A _07574_/B _07574_/C vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__and3_1
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _11237_/S _09250_/B vssd1 vssd1 vccd1 vccd1 _09252_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07949__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _09171_/X _09174_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09175_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08126_ _08124_/A _08124_/B _08203_/A vssd1 vssd1 vccd1 vccd1 _08138_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08958__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09080__B1 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__B2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ _08057_/A _08057_/B vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07008_ _07009_/A _07009_/B vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07684__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08959_ _09787_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__xnor2_1
X_11970_ _11964_/Y _11965_/X _11969_/X vssd1 vssd1 vccd1 vccd1 _11971_/C sky130_fd_sc_hd__o21a_1
X_10921_ _10921_/A _10921_/B _10921_/C vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__and3_1
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__A3 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10852_ _10852_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10048__A3 _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10666_/B _10666_/C _10666_/A vssd1 vssd1 vccd1 vccd1 _10785_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12523_/A _12523_/B _12523_/C vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__a21o_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08110__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _12453_/A _12453_/B _12453_/C vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08949__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ _12383_/A _12383_/B _12029_/A vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09610__A2 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08949__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11335_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11335_/Y sky130_fd_sc_hd__nor2_1
X_11266_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11267_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13005_ _13300_/Q _12781_/A _13209_/A2 hold242/X vssd1 vssd1 vccd1 vccd1 hold243/A
+ sky130_fd_sc_hd__a22o_1
X_10217_ _11813_/A _10217_/B vssd1 vssd1 vccd1 vccd1 _10221_/A sky130_fd_sc_hd__xnor2_1
X_11197_ _11197_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11181__A1 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__B2 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10148_ _09565_/X _09570_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__mux2_1
X_10079_ _09917_/A _09917_/B _09914_/A vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12130__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09429__A2 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12433__A1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07290_ _09787_/A _07290_/B vssd1 vssd1 vccd1 vccd1 _07398_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10195__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__buf_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09195__S _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09862_ _09863_/B _09863_/C _10319_/A vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07376__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06718__A3 _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09814_/A sky130_fd_sc_hd__xor2_1
X_08813_ _07584_/A _07584_/B _07587_/A vssd1 vssd1 vccd1 vccd1 _08824_/A sky130_fd_sc_hd__a21o_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _08739_/X _08740_/Y _08743_/B _08743_/A _08737_/Y vssd1 vssd1 vccd1 vccd1
+ _08750_/A sky130_fd_sc_hd__a221o_2
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11475__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08675_/A _08675_/B vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__nor2_2
XANTENNA__08876__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07627_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ _07661_/A _07661_/B _07491_/X vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__12975__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07679__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07488_ _07488_/A _07488_/B vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ _09233_/A _09227_/B vssd1 vssd1 vccd1 vccd1 _09227_/X sky130_fd_sc_hd__or2_1
XANTENNA__12188__B1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ reg1_val[3] reg1_val[28] _09180_/S vssd1 vssd1 vccd1 vccd1 _09158_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ _09297_/A1 fanout13/X fanout11/X _09297_/B2 vssd1 vssd1 vccd1 vccd1 _09090_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07603__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08109_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _11781_/S _11120_/B vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ _11980_/A fanout46/X fanout45/X fanout57/X vssd1 vssd1 vccd1 vccd1 _11052_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07367__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _12339_/A1 _10038_/A _10313_/A _11889_/A1 vssd1 vssd1 vccd1 vccd1 _10002_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__07906__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11953_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11953_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11884_ reg1_val[22] _06993_/A _09595_/B _11883_/X vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10674__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ _11131_/A _09737_/X _10903_/X vssd1 vssd1 vccd1 vccd1 _10904_/Y sky130_fd_sc_hd__a21oi_2
X_10835_ _10933_/A _10835_/B vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08619__B1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ _10527_/X _10646_/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10697_ _10870_/B _10697_/B vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__nand2_1
X_12505_ _12666_/B _12506_/B vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09300__C _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07842__B2 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07842__A1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ _12414_/X _12418_/X _12434_/X _12435_/Y vssd1 vssd1 vccd1 vccd1 dest_val[31]
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08398__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12367_ _12366_/A _12366_/B _12366_/C vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06940__B _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11318_ _11318_/A _11318_/B _11318_/C vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12298_ hold307/A _12349_/A _12348_/B _12393_/B1 vssd1 vssd1 vccd1 vccd1 _12298_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11154__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13143__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11249_ _11249_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__and3_1
XANTENNA__11154__B2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ _06799_/A _06801_/B1 _12632_/B _06788_/X vssd1 vssd1 vccd1 vccd1 _06790_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__xnor2_1
X_07411_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07413_/C sky130_fd_sc_hd__xnor2_1
X_08391_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07342_ reg1_val[26] reg1_val[27] _07342_/C vssd1 vssd1 vccd1 vccd1 _12756_/B sky130_fd_sc_hd__or3_4
XANTENNA__07499__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12957__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _07273_/A _07273_/B _07359_/A vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09012_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11749__A _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09219__A _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08123__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11145__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09914_ _09914_/A _09914_/B vssd1 vssd1 vccd1 vccd1 _09917_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09889__A2 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _09843_/A _09843_/B _09846_/B vssd1 vssd1 vccd1 vccd1 _09845_/Y sky130_fd_sc_hd__a21oi_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ reg1_val[4] _06988_/B vssd1 vssd1 vccd1 vccd1 _06990_/B sky130_fd_sc_hd__xor2_2
X_09776_ _09776_/A _09776_/B vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__nor2_2
X_08727_ _08726_/A _08726_/C _08726_/B vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08849__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08710_/A sky130_fd_sc_hd__xnor2_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13341_/CLK sky130_fd_sc_hd__clkbuf_8
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _07611_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10828__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08588_/A _08588_/C _08588_/B vssd1 vssd1 vccd1 vccd1 _08595_/B sky130_fd_sc_hd__a21o_1
X_10620_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10696_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13070__A1 _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11081__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _09391_/X _09405_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07202__A _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13270_ _13375_/CLK hold116/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__dfxtp_1
X_10482_ fanout42/X _07243_/X _07250_/X fanout40/X vssd1 vssd1 vccd1 vccd1 _10483_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12374_/D _12279_/B _12279_/C _12280_/A vssd1 vssd1 vccd1 vccd1 _12221_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__B2 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__A_N _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _12324_/B _12324_/C vssd1 vssd1 vccd1 vccd1 _12270_/A sky130_fd_sc_hd__nor2_2
XANTENNA__08033__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__xnor2_1
X_12083_ _12083_/A _12083_/B _12083_/C vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11809__D _11809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _11131_/A _09573_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ hold326/X _13143_/B2 _13186_/A2 hold216/X vssd1 vssd1 vccd1 vccd1 hold217/A
+ sky130_fd_sc_hd__a22o_1
X_11936_ _11766_/A _11852_/A _11851_/A vssd1 vssd1 vccd1 vccd1 _11936_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11867_ _11865_/X _11947_/B instruction[7] vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10818_ _10822_/A vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__inv_2
X_11798_ _12395_/A1 _11797_/X _06682_/B vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10749_ _10602_/A _10602_/B _10600_/Y vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xload_slew1 _07066_/Y vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06951__A _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12672__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06670__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12420_/A _12420_/B _12420_/C vssd1 vssd1 vccd1 vccd1 _12419_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _07959_/B _07959_/C _07959_/A vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__o21ba_1
X_06911_ instruction[13] _06913_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
XANTENNA__07782__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ _12619_/A _07891_/B _07891_/C vssd1 vssd1 vccd1 vccd1 _07894_/B sky130_fd_sc_hd__and3_1
X_06842_ reg1_val[20] _06996_/A vssd1 vssd1 vccd1 vccd1 _06842_/Y sky130_fd_sc_hd__nand2_1
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06773_ _06774_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _10008_/A sky130_fd_sc_hd__nor2_1
X_09561_ _09159_/X _09163_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__mux2_1
X_08512_ _08510_/A _08510_/B _08511_/Y vssd1 vssd1 vccd1 vccd1 _08515_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12847__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ _11168_/A _09492_/B vssd1 vssd1 vccd1 vccd1 _09493_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09256__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08374_ _08573_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _08409_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11063__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07325_ _07325_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07327_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07256_ fanout77/X fanout75/X fanout73/X fanout71/X vssd1 vssd1 vccd1 vccd1 _07257_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06580__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _07208_/B _07188_/C reg1_val[19] vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07034__A2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ fanout31/X _07237_/Y _07243_/X fanout28/X vssd1 vssd1 vccd1 vccd1 _09829_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _10315_/A _09904_/A vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__or2_1
XANTENNA__07742__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12770_/A _12770_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12053_/A1 _11717_/X _11720_/X vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11652_ _12202_/B _07155_/Y _12257_/A _07151_/Y vssd1 vssd1 vccd1 vccd1 _11653_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _10504_/A _10504_/B _10501_/A vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout61 _06999_/X vssd1 vssd1 vccd1 vccd1 fanout61/X sky130_fd_sc_hd__buf_4
Xfanout83 _11296_/A vssd1 vssd1 vccd1 vccd1 fanout83/X sky130_fd_sc_hd__buf_8
Xfanout72 _07254_/X vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__buf_6
Xfanout50 _07059_/X vssd1 vssd1 vccd1 vccd1 fanout50/X sky130_fd_sc_hd__buf_6
X_11583_ _11584_/B _11584_/A vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__nand2b_1
Xfanout94 _07126_/Y vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__buf_8
X_13322_ _13323_/CLK _13322_/D vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12492__B _12492_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ _10534_/A _10769_/A vssd1 vssd1 vccd1 vccd1 _10534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _13372_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_10465_ _07593_/A _07593_/B fanout85/X vssd1 vssd1 vccd1 vccd1 _10468_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13184_/Y sky130_fd_sc_hd__xnor2_1
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12206_/B sky130_fd_sc_hd__xor2_1
X_10396_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10396_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07078__S _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ _12134_/B _12135_/B vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_19_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _12138_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12070_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13109__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11018_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10096__A1 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ _12978_/A hold258/X vssd1 vssd1 vccd1 vccd1 _13282_/D sky130_fd_sc_hd__and2_1
XANTENNA__06946__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _11998_/A _11919_/B vssd1 vssd1 vccd1 vccd1 _11921_/B sky130_fd_sc_hd__nor2_1
X_12899_ hold29/X hold309/X vssd1 vssd1 vccd1 vccd1 _13110_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10096__B2 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13034__A1 _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07110_ _07109_/A _07109_/B _07109_/C _07109_/D vssd1 vssd1 vccd1 vccd1 _11823_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _08553_/A2 fanout82/X _08551_/B1 _08400_/B vssd1 vssd1 vccd1 vccd1 _08091_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07041_ reg1_val[4] reg1_val[5] vssd1 vssd1 vccd1 vccd1 _07063_/D sky130_fd_sc_hd__or2_1
XFILLER_0_42_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10931__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _09675_/A _07347_/B fanout15/X _09467_/A vssd1 vssd1 vccd1 vccd1 _08993_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12848__A1 wire8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07943_ _10081_/A _07943_/B vssd1 vssd1 vccd1 vccd1 _07947_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06688__A_N _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A _13227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__S _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _07873_/B _07873_/C _07873_/A vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__o21ba_1
X_06825_ _07175_/A reg1_val[12] vssd1 vssd1 vccd1 vccd1 _06825_/X sky130_fd_sc_hd__and2b_1
X_09613_ fanout41/X _10326_/A _07218_/Y _07402_/B vssd1 vssd1 vccd1 vccd1 _09614_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06756_ _06799_/A _06801_/B1 _12657_/B _06755_/X vssd1 vssd1 vccd1 vccd1 _07202_/A
+ sky130_fd_sc_hd__a31o_4
X_09544_ _09544_/A _09706_/A _09858_/A _09996_/A vssd1 vssd1 vccd1 vccd1 _10129_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ reg2_val[19] _06712_/B _06707_/B1 _06686_/Y vssd1 vssd1 vccd1 vccd1 _07058_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _10230_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__xnor2_1
X_08426_ _08426_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _08459_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09886__B _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _09941_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08288_ _08445_/A _08288_/B vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07308_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07310_/B sky130_fd_sc_hd__xnor2_2
X_07239_ _07236_/A _07236_/B _09787_/A vssd1 vssd1 vccd1 vccd1 _07239_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10250_ _10117_/A _10117_/B _10115_/X vssd1 vssd1 vccd1 vccd1 _10258_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _11052_/A _10181_/B vssd1 vssd1 vccd1 vccd1 _10185_/A sky130_fd_sc_hd__xnor2_1
Xfanout273 _06573_/X vssd1 vssd1 vccd1 vccd1 _06699_/B sky130_fd_sc_hd__clkbuf_8
Xfanout262 _06944_/X vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__clkbuf_8
Xfanout251 _06766_/X vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__buf_4
XANTENNA__10811__A_N _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08507__A2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 instruction[7] vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__buf_4
Xfanout284 _12025_/S vssd1 vssd1 vccd1 vccd1 _11781_/S sky130_fd_sc_hd__clkbuf_8
X_12822_ _07067_/Y _12782_/Y hold140/X _13226_/A vssd1 vssd1 vccd1 vccd1 _13260_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12067__A2 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ reg1_val[28] _12773_/A vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__and2_1
X_11704_ _11238_/S _10801_/Y _11703_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _11715_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ reg1_val[13] _12685_/B vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__nand2_1
X_11635_ _12053_/A1 _11632_/X _11634_/Y vssd1 vssd1 vccd1 vccd1 dest_val[19] sky130_fd_sc_hd__o21ai_4
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11567_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07597__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13305_ _13372_/CLK hold164/X vssd1 vssd1 vccd1 vccd1 hold162/A sky130_fd_sc_hd__dfxtp_1
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__nand2_1
X_13236_ _13236_/A _13236_/B hold155/X vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__and3_1
XFILLER_0_122_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10448_ fanout56/X fanout27/X fanout25/X fanout62/X vssd1 vssd1 vccd1 vccd1 _10449_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ hold281/X _13166_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__mux2_1
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _09222_/Y _10146_/X _10152_/X _09155_/S _12117_/Y vssd1 vssd1 vccd1 vccd1
+ _12118_/X sky130_fd_sc_hd__a221o_1
X_13098_ hold271/X _13097_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09317__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ _12023_/X _12027_/X _12048_/X _11975_/A vssd1 vssd1 vccd1 vccd1 _12049_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07182__A1 _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _06706_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _06610_/Y sky130_fd_sc_hd__nor2_1
X_07590_ _06851_/B _07300_/A _07074_/B _08971_/A vssd1 vssd1 vccd1 vccd1 _07593_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10069__A1 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__B2 _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _10310_/A _10310_/B _12420_/A vssd1 vssd1 vccd1 vccd1 _09260_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08211_ _08259_/A _08259_/B _08172_/X vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09191_ _09187_/X _09190_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09191_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _08142_/A _08142_/B vssd1 vssd1 vccd1 vccd1 _08143_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ _06875_/A fanout98/X fanout83/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08074_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ _08650_/A _07024_/B vssd1 vssd1 vccd1 vccd1 _07039_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09934__A1 _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B2 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _09670_/A _08975_/B vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08131__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _07937_/B _07937_/A vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__and2b_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07970__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _07864_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__and2b_1
X_06808_ _09743_/A _09739_/B _06807_/Y vssd1 vssd1 vccd1 vccd1 _06808_/Y sky130_fd_sc_hd__o21ai_1
X_07788_ _07788_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__xnor2_1
X_06739_ reg2_val[10] _06767_/A vssd1 vssd1 vccd1 vccd1 _06739_/X sky130_fd_sc_hd__and2_1
X_09527_ _09351_/A _09351_/B _09354_/A vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__a21o_2
XANTENNA__08122__B1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout27_A _07211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _09458_/A _09458_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09459_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10480__B2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__A1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _09180_/X _09200_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08409_ _08409_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__nand2_1
X_11420_ _11595_/A _11420_/B vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _09196_/S _11237_/X _11346_/X _11350_/X vssd1 vssd1 vccd1 vccd1 _11351_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08976__A2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _10302_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10302_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ _11285_/A vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08189__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _10233_/A1 fanout11/X fanout7/X _10233_/B2 vssd1 vssd1 vccd1 vccd1 _10234_/B
+ sky130_fd_sc_hd__o22a_1
X_13021_ hold18/X _13055_/A2 _13053_/B1 _13309_/Q _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold19/A sky130_fd_sc_hd__o221a_1
XANTENNA__11386__B _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07400__A2 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ _09831_/A _09831_/B _09954_/B _09955_/B _09955_/A vssd1 vssd1 vccd1 vccd1
+ _10109_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__09571__S _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__A _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13237__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ hold32/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__or2_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10997_ _10998_/A _10998_/B _10998_/C vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11799__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11799__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ _12741_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12740_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_29_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12437__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12676_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11618_ _11958_/A _11618_/B vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09613__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ _12598_/A _12598_/B _12598_/C _12598_/D vssd1 vssd1 vccd1 vccd1 _12600_/C
+ sky130_fd_sc_hd__or4_1
X_11549_ _11548_/B _11549_/B vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _13219_/A hold288/X vssd1 vssd1 vccd1 vccd1 _13367_/D sky130_fd_sc_hd__and2_1
XANTENNA__10481__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11296__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13324_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _08760_/A _08760_/B _11512_/A vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__and3_1
XANTENNA__08886__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__and2_1
X_08691_ _08161_/Y _08165_/Y _08166_/X vssd1 vssd1 vccd1 vccd1 _08691_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07642_ _07642_/A _07642_/B vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12987__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ _11361_/A _09312_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__xnor2_1
X_07573_ _07573_/A _11813_/A vssd1 vssd1 vccd1 vccd1 _07574_/C sky130_fd_sc_hd__or2_1
XFILLER_0_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout231_A _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _12772_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__nor2_2
XANTENNA__10656__A _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06853__B _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _09172_/X _09173_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10214__A1 _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08125_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__or2_1
XANTENNA__08958__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09080__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A1 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07965__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08056_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__nand2_1
X_07007_ _07009_/A _07009_/B vssd1 vssd1 vccd1 vccd1 _07011_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08591__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ fanout50/X fanout85/X _10466_/A _09659_/B2 vssd1 vssd1 vccd1 vccd1 _08959_/B
+ sky130_fd_sc_hd__o22a_1
X_07909_ _10233_/B2 _08354_/A2 _10585_/B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _07910_/B
+ sky130_fd_sc_hd__o22a_1
X_08889_ _08944_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _08891_/C sky130_fd_sc_hd__or2_1
XFILLER_0_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10920_ _07175_/A _06940_/B _10919_/Y vssd1 vssd1 vccd1 vccd1 _10921_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _10852_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _10972_/C sky130_fd_sc_hd__or2_1
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10785_/B sky130_fd_sc_hd__or2_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11650__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _12530_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12523_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12452_ _12453_/A _12453_/B _12453_/C vssd1 vssd1 vccd1 vccd1 _12460_/B sky130_fd_sc_hd__a21o_1
X_11403_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12781__A _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _12383_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12383_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11334_ _11232_/B _11234_/B _11230_/X vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11265_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand2_1
X_13004_ _13134_/A hold189/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__and2_1
X_10216_ _07212_/X _07581_/A _07581_/B _07345_/X _10712_/A vssd1 vssd1 vccd1 vccd1
+ _10217_/B sky130_fd_sc_hd__a32o_1
XANTENNA__07909__B1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _11097_/A _11097_/B _11095_/Y vssd1 vssd1 vccd1 vccd1 _11205_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11181__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ _09562_/X _09564_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _10147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12130__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__A1 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12418__C1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12969__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _12737_/A _12719_/B _12719_/C vssd1 vssd1 vccd1 vccd1 _12720_/B sky130_fd_sc_hd__and3_2
XFILLER_0_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold315 hold315/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09930_ _09930_/A _09930_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09861_ _10128_/A _09546_/X _10267_/A _09860_/X vssd1 vssd1 vccd1 vccd1 _09863_/C
+ sky130_fd_sc_hd__o31a_2
XANTENNA__07376__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07376__B2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__nand2_1
X_08812_ _07612_/A _07612_/B _07610_/Y vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__o21ai_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _08743_/B vssd1 vssd1 vccd1 vccd1 _08743_/X sky130_fd_sc_hd__and2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout279_A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout181_A _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08876__B2 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__A1 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _08543_/A _08675_/B _08675_/A vssd1 vssd1 vccd1 vccd1 _08674_/X sky130_fd_sc_hd__o21ba_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__B2 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10683__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07625_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07625_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07556_ _07556_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__B2 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _09233_/A _09227_/B vssd1 vssd1 vccd1 vccd1 _09226_/Y sky130_fd_sc_hd__nor2_8
X_07487_ _07487_/A _07487_/B vssd1 vssd1 vccd1 vccd1 _07488_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ reg1_val[2] reg1_val[29] _09180_/S vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07603__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _10081_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__xnor2_1
X_09088_ _09280_/B _09088_/B vssd1 vssd1 vccd1 vccd1 _09099_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _08069_/A _08069_/B _08034_/Y vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07367__B2 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _12420_/A _10038_/A _10313_/A vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06758__B _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _11951_/A _11951_/B _11951_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _11972_/C
+ sky130_fd_sc_hd__o211a_1
X_11883_ _09228_/Y _11966_/B _11883_/S vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__mux2_1
X_10903_ _11235_/S _09877_/X _10902_/X _11237_/S vssd1 vssd1 vccd1 vccd1 _10903_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ _11734_/A _07151_/A _07155_/A _11568_/A vssd1 vssd1 vccd1 vccd1 _10835_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08619__B2 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__A1 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10765_ _10765_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__or2_2
X_12504_ reg1_val[10] curr_PC[10] _12504_/S vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09292__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10696_ _10696_/A _10696_/B _10696_/C vssd1 vssd1 vccd1 vccd1 _10697_/B sky130_fd_sc_hd__or3_1
XANTENNA__07842__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _07127_/B _11446_/B _12504_/S vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ _12366_/A _12366_/B _12366_/C vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__and3_1
X_11317_ _11318_/A _11318_/B _11318_/C vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12297_ _12349_/A _12348_/B hold307/A vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11248_ _07243_/A _06940_/B _11247_/Y vssd1 vssd1 vccd1 vccd1 _11249_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11154__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _11179_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06949__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__B _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _07410_/A _07423_/A vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__nor2_2
X_08390_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09807__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07351_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07272_ _07273_/B _07359_/A _07273_/A vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _09012_/B _09012_/A vssd1 vssd1 vccd1 vccd1 _09011_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__B _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10653__B _10653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _09913_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__nor2_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09844_ _09684_/A _09684_/B _09682_/Y vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__a21oi_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10353__B1 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06578__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ reg1_val[3] _06987_/B vssd1 vssd1 vccd1 vccd1 _06987_/Y sky130_fd_sc_hd__xnor2_1
X_09775_ _09775_/A _09775_/B _09775_/C vssd1 vssd1 vccd1 vccd1 _09776_/B sky130_fd_sc_hd__and3_1
X_08726_ _08726_/A _08726_/B _08726_/C vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08849__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09510__A2 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__xor2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13055__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07608_ _07609_/B _07609_/A vssd1 vssd1 vccd1 vccd1 _07608_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08588_ _08588_/A _08588_/B _08588_/C vssd1 vssd1 vccd1 vccd1 _08595_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13070__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ _08476_/A _07539_/B _07690_/B vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__and3_1
XANTENNA__11081__B2 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11081__A1 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10550_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07285__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ _11296_/B _10481_/B vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09207_/X _09208_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09209_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12220_ _12270_/B _12220_/B vssd1 vssd1 vccd1 vccd1 _12279_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__B2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _12151_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12324_/C sky130_fd_sc_hd__and3_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _11103_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__nand2_1
X_12082_ _12083_/A _12083_/B _12083_/C vssd1 vssd1 vccd1 vccd1 _12082_/Y sky130_fd_sc_hd__a21oi_2
X_11033_ _11033_/A _11033_/B _11033_/C vssd1 vssd1 vccd1 vccd1 _11033_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__10895__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ _13144_/A hold246/X vssd1 vssd1 vccd1 vccd1 _13290_/D sky130_fd_sc_hd__and2_1
X_11935_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_87_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11866_ _11782_/A _11779_/X _06841_/Y vssd1 vssd1 vccd1 vccd1 _11947_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ _11169_/A _10817_/B vssd1 vssd1 vccd1 vccd1 _10822_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11797_ _09886_/B _12394_/A1 _11797_/S vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10748_ _10626_/A _10625_/B _10625_/A vssd1 vssd1 vccd1 vccd1 _10753_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10679_ hold308/A _11029_/A2 _10796_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _10679_/X
+ sky130_fd_sc_hd__a31o_1
X_12418_ _12417_/A _12417_/B _12417_/Y _11612_/A vssd1 vssd1 vccd1 vccd1 _12418_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__06951__B _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__A1 _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08224__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ _12349_/A _12391_/B vssd1 vssd1 vccd1 vccd1 _12349_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06910_ instruction[12] _06913_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
XANTENNA__06679__A _06964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07200__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _07953_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _07954_/A sky130_fd_sc_hd__nor2_1
X_06841_ reg1_val[21] _06964_/B vssd1 vssd1 vccd1 vccd1 _06841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _09560_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__nor2_1
X_06772_ reg1_val[5] _06952_/C vssd1 vssd1 vccd1 vccd1 _06772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09491_ fanout52/X fanout77/X fanout73/X fanout50/X vssd1 vssd1 vccd1 vccd1 _09492_/B
+ sky130_fd_sc_hd__o22a_1
X_08511_ _08545_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08455_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13037__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08373_ _08572_/A2 _08553_/A2 _08551_/B1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 _08374_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout144_A _07054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11063__A1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__B2 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07324_ _07325_/B vssd1 vssd1 vccd1 vccd1 _07324_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07255_ _07255_/A _07255_/B vssd1 vssd1 vccd1 vccd1 _07255_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07019__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07186_ reg1_val[18] reg1_val[31] _12335_/A vssd1 vssd1 vccd1 vccd1 _07188_/C sky130_fd_sc_hd__and3_1
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__xnor2_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07742__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _09758_/A _10310_/C _09710_/Y vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__nor3b_1
XANTENNA__07742__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout57_A _07015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08709_ _08624_/A _08658_/A _08652_/X _08707_/A vssd1 vssd1 vccd1 vccd1 _08710_/B
+ sky130_fd_sc_hd__o31ai_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11434__S _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _12525_/S _11892_/C _11720_/C vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__or3_2
X_09689_ _09526_/A _09526_/B _09525_/A vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ _12310_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__xnor2_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 fanout41/X vssd1 vssd1 vccd1 vccd1 fanout40/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07213__A _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09247__A1 _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10602_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__xor2_2
Xfanout62 _06994_/Y vssd1 vssd1 vccd1 vccd1 fanout62/X sky130_fd_sc_hd__buf_8
XFILLER_0_92_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 fanout74/X vssd1 vssd1 vccd1 vccd1 fanout73/X sky130_fd_sc_hd__buf_6
Xfanout51 _07059_/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__buf_4
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout95 _07096_/X vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__buf_8
X_13321_ _13323_/CLK _13321_/D vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__dfxtp_1
X_10533_ _10270_/A _10769_/A _10530_/Y vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__a21o_1
Xfanout84 _07238_/X vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__buf_6
XANTENNA__10574__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _13350_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
X_10464_ _10735_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ _13187_/A hold300/X vssd1 vssd1 vccd1 vccd1 _13359_/D sky130_fd_sc_hd__and2_1
X_12203_ _12404_/B _12203_/B _12202_/X vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__or3b_1
X_10395_ _10256_/A _10256_/B _10254_/Y vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12134_ _12135_/B _12134_/B vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07883__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12065_ _12065_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__nand2_1
X_11016_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11018_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ hold247/X _13095_/B2 _13158_/A2 hold257/X vssd1 vssd1 vccd1 vccd1 hold258/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09486__A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B2 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A1 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ fanout57/X _11988_/A _11916_/Y vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10096__A2 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ _13105_/A _13106_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__13019__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _11850_/A _11850_/B _11850_/C vssd1 vssd1 vccd1 vccd1 _11852_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07123__A _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12964__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ _07082_/A _07082_/B vssd1 vssd1 vccd1 vccd1 _07084_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10556__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _08865_/A _08865_/B _08863_/X vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12848__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _08553_/B1 _08184_/B fanout32/X _09468_/B2 vssd1 vssd1 vccd1 vccd1 _07943_/B
+ sky130_fd_sc_hd__o22a_1
X_07873_ _07873_/A _07873_/B _07873_/C vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__or3_1
X_06824_ _10779_/A _06822_/X _06823_/X vssd1 vssd1 vccd1 vccd1 _06824_/Y sky130_fd_sc_hd__o21bai_1
X_09612_ _09612_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09616_/B sky130_fd_sc_hd__xor2_1
X_09543_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06755_ reg2_val[7] _06794_/B vssd1 vssd1 vccd1 vccd1 _06755_/X sky130_fd_sc_hd__and2_1
X_06686_ _06706_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _06686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ fanout58/X _10463_/B2 _10228_/A fanout56/X vssd1 vssd1 vccd1 vccd1 _09475_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08129__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07033__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ _08425_/A _08425_/B vssd1 vssd1 vccd1 vccd1 _08746_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11036__A1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ _08619_/B2 _08521_/A2 _08551_/A2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08357_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12784__A1 _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ _08553_/B1 _10227_/B1 _10463_/A1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 _08288_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07238_ _07074_/A _07073_/X _07074_/Y _06959_/Y vssd1 vssd1 vccd1 vccd1 _07238_/X
+ sky130_fd_sc_hd__a22o_1
X_07169_ _11168_/A _07180_/C vssd1 vssd1 vccd1 vccd1 _07169_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ _11386_/A fanout46/X fanout44/X _11296_/A vssd1 vssd1 vccd1 vccd1 _10181_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout230 _09420_/X vssd1 vssd1 vccd1 vccd1 _10158_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout241 _06939_/X vssd1 vssd1 vccd1 vccd1 _11446_/B sky130_fd_sc_hd__clkbuf_8
Xfanout274 _06573_/X vssd1 vssd1 vccd1 vccd1 _06657_/B sky130_fd_sc_hd__buf_2
Xfanout252 _06631_/A vssd1 vssd1 vccd1 vccd1 _06801_/B1 sky130_fd_sc_hd__buf_8
Xfanout263 _06944_/X vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__buf_4
Xfanout285 _12378_/S vssd1 vssd1 vccd1 vccd1 _12025_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__06923__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ hold139/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09468__A1 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12752_ _12752_/A _12757_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
X_11703_ _11958_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11703_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12688_/B _12683_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XANTENNA__07138__A_N _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12224__B1 _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ curr_PC[19] _11718_/C _11633_/Y vssd1 vssd1 vccd1 vccd1 _11634_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__09569__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11496_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__xnor2_2
X_13304_ _13372_/CLK _13304_/D vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
X_10516_ _10515_/A _10515_/B _10517_/A vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10447_ _11169_/A _10447_/B vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__xnor2_1
X_13235_ hold202/A hold193/A hold149/X hold154/X vssd1 vssd1 vccd1 vccd1 hold155/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10538__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13166_ _13166_/A _13166_/B vssd1 vssd1 vccd1 vccd1 _13166_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__nor2_1
X_12117_ _06978_/A _06939_/X _12116_/X vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__o21ai_1
X_13097_ _13097_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13097_/Y sky130_fd_sc_hd__xnor2_1
X_12048_ _12107_/B1 _12036_/X _12047_/Y _12030_/Y vssd1 vssd1 vccd1 vccd1 _12048_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11863__A _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__B _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13007__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08217_/A _08217_/B _08199_/X vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06692__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _09188_/X _09189_/X _09396_/S vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _08141_/A _08141_/B vssd1 vssd1 vccd1 vccd1 _08142_/B sky130_fd_sc_hd__and2_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08072_ _08072_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08103_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07023_ fanout64/X _09297_/B2 fanout58/X _09297_/A1 vssd1 vssd1 vccd1 vccd1 _07024_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__A _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_A _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11741__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08974_ _06973_/Y fanout11/X fanout7/X _06973_/A vssd1 vssd1 vccd1 vccd1 _08975_/B
+ sky130_fd_sc_hd__o22a_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _07925_/A _07925_/B vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__xnor2_2
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07864_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09243__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ reg1_val[3] _10902_/A vssd1 vssd1 vccd1 vccd1 _06807_/Y sky130_fd_sc_hd__nand2_1
X_07787_ _07806_/A _07806_/B _07767_/X vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__a21bo_1
X_06738_ _10794_/S _06738_/B vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__nor2_1
X_09526_ _09526_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__xor2_4
X_09457_ _09458_/A _09458_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08122__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06669_ _11883_/S _06669_/B vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__nor2_2
X_08408_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08412_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10480__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _09177_/X _09179_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10768__B1 _10766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _08392_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08339_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11350_ _09222_/Y _11339_/B _11348_/Y _11349_/X vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10299_/Y _10301_/B vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _12310_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__xnor2_1
X_13020_ _07009_/B _12797_/B hold161/X vssd1 vssd1 vccd1 vccd1 _13308_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__08189__B2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13182__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _10231_/B _10231_/C _10231_/A vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09418__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10940__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10094_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12498__B _12499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09153__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _07218_/Y _12782_/Y hold39/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__o211a_1
XANTENNA__11248__A1 _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10998_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ reg1_val[24] _12773_/A vssd1 vssd1 vccd1 vccd1 _12736_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ reg1_val[10] _12666_/B vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__or2_1
XFILLER_0_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ _12616_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__xnor2_4
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09613__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07401__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ _11549_/B _11548_/B vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07120__B _12717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09613__B2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ _11480_/B _11479_/B vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ hold287/X _13222_/A2 _13217_/X _12781_/A vssd1 vssd1 vccd1 vccd1 hold288/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13173__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13149_ _13187_/A hold312/X vssd1 vssd1 vccd1 vccd1 _13352_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11593__A _11593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _09630_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08690_ _07997_/A _07997_/B _08689_/X vssd1 vssd1 vccd1 vccd1 _08690_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13228__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07641_ _07642_/A _07642_/B vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__and2_1
X_07572_ reg1_val[29] _07572_/B vssd1 vssd1 vccd1 vccd1 _07572_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _11386_/A _08184_/B fanout32/X _11296_/A vssd1 vssd1 vccd1 vccd1 _09312_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10937__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09242_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08407__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09173_ reg1_val[11] reg1_val[20] _09180_/S vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10214__A2 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _08124_/A _08124_/B vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07615__B1 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08055_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07006_ _07009_/A _07009_/B vssd1 vssd1 vccd1 vccd1 _07010_/A sky130_fd_sc_hd__and2_1
XANTENNA__08591__A1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__B2 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13194__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _09064_/B _08957_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__nor2_1
X_07908_ _07908_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__xor2_1
X_08888_ _08888_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__nor2_1
X_07839_ _07845_/B _07845_/A vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__and2b_1
X_10850_ _11296_/B _10850_/B vssd1 vssd1 vccd1 vccd1 _10852_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12427__B1 _09239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__nand2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09795_/A _09509_/B vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__xnor2_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11650__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11650__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12520_ _12679_/B _12520_/B vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__or2_1
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08317__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12451_ _12460_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12453_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07606__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12382_ _08809_/A _08808_/Y _12420_/A vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11333_ _11333_/A _11333_/B vssd1 vssd1 vccd1 vccd1 _11333_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _11559_/A _11264_/B vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11166__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ hold188/X _13143_/B2 _13209_/A2 _13300_/Q vssd1 vssd1 vccd1 vccd1 hold189/A
+ sky130_fd_sc_hd__a22o_1
X_10215_ _10384_/B _10215_/B vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__or2_1
XANTENNA__07909__A1 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _11090_/A _11089_/B _11087_/Y vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07891__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _11131_/A _10145_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__o21a_1
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12130__A2 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ _10864_/A _10864_/B _10867_/A vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12448__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ _12719_/B _12719_/C _12737_/A vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__08227__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12972__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ _12649_/A _12649_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xor2_4
XANTENNA__06970__A _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12691__B _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09860_ _09541_/X _09703_/X _09704_/X vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07376__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10380__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _09791_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__nand2_1
X_08811_ _07653_/A _07653_/B _07654_/Y vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__o21ai_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08680_/C _08680_/D _08746_/A vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__a21o_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _08673_/A _08673_/B _08673_/C vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07306__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07624_ _08891_/B _07624_/B vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__and2_1
XANTENNA__08876__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07555_ _07553_/A _07553_/B _07554_/Y vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__11632__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07486_ _07486_/A _07486_/B vssd1 vssd1 vccd1 vccd1 _07487_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _09238_/B _09229_/B vssd1 vssd1 vccd1 vccd1 _09225_/X sky130_fd_sc_hd__or2_2
XFILLER_0_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09154_/X _09155_/X _12785_/A vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09087_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08107_ _08619_/B1 _08184_/B fanout32/X _09403_/S vssd1 vssd1 vccd1 vccd1 _08108_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout87_A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _10319_/B _10000_/B vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07367__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08316__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08316__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11882_ hold199/A _11529_/B _11960_/B _11242_/A vssd1 vssd1 vccd1 vccd1 _11882_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10674__A2 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _10902_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__or2_1
X_10833_ _10833_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13073__B1 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A1 _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__A2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10764_ _10764_/A _10764_/B _10764_/C vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__and3_1
XANTENNA__07827__A0 _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ _12509_/B _12503_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ _10696_/A _10696_/B _10696_/C vssd1 vssd1 vccd1 vccd1 _10870_/B sky130_fd_sc_hd__o21ai_1
X_12434_ _11946_/A _12419_/Y _12420_/X _12433_/X vssd1 vssd1 vccd1 vccd1 _12434_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12365_ _12365_/A _12365_/B vssd1 vssd1 vccd1 vccd1 _12366_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11316_ _11316_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11318_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ hold301/A _12296_/B vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__or2_1
X_11247_ _12395_/A1 _11246_/X _06716_/B vssd1 vssd1 vccd1 vccd1 _11247_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08004__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11179_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__and2_1
XANTENNA__06949__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _10129_/A _10129_/B _10129_/C vssd1 vssd1 vccd1 vccd1 _10129_/X sky130_fd_sc_hd__or3_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06965__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07340_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07271_ _07358_/A _07358_/B vssd1 vssd1 vccd1 vccd1 _07359_/A sky130_fd_sc_hd__and2_1
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09012_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10050__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _09913_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__and2_1
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10353__A1 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__nand2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10353__B2 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _12619_/A _12621_/A reg1_val[2] _07093_/A vssd1 vssd1 vccd1 vccd1 _06987_/B
+ sky130_fd_sc_hd__o31a_1
X_09774_ _09775_/A _09775_/B _09775_/C vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__a21oi_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08725_ _08720_/A _08720_/B _08581_/X _08599_/X vssd1 vssd1 vccd1 vccd1 _08726_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08849__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06875__A _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _09670_/A _08656_/B _09553_/B vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__or3_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ _08576_/A _08575_/C _08575_/B vssd1 vssd1 vccd1 vccd1 _08588_/C sky130_fd_sc_hd__a21o_1
X_07607_ _10234_/A _07607_/B vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06594__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ _09827_/A _07538_/B vssd1 vssd1 vccd1 vccd1 _07690_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11081__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07814_/B _09675_/A _09467_/A fanout45/X vssd1 vssd1 vccd1 vccd1 _07470_/B
+ sky130_fd_sc_hd__o22a_1
X_10480_ _10585_/B2 fanout9/A fanout5/X _10589_/A vssd1 vssd1 vccd1 vccd1 _10481_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09397__S _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ reg1_val[10] reg1_val[21] _09560_/A vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12150_ _12151_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12324_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07588__A2 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _11101_/A _11101_/B vssd1 vssd1 vccd1 vccd1 _11103_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ _12151_/B _12081_/B vssd1 vssd1 vccd1 vccd1 _12083_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ _07255_/A _06940_/B _11031_/Y vssd1 vssd1 vccd1 vccd1 _11033_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09734__B1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B1 _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__B _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ hold210/X _13143_/B2 _13186_/A2 hold245/X vssd1 vssd1 vccd1 vccd1 hold246/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11934_ _11934_/A vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__inv_2
XFILLER_0_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ _11782_/A _11780_/X _11797_/S vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816_ fanout74/X fanout13/X fanout12/X _08274_/B vssd1 vssd1 vccd1 vccd1 _10817_/B
+ sky130_fd_sc_hd__o22a_1
X_11796_ hold249/A _11529_/B _11880_/B _11242_/A vssd1 vssd1 vccd1 vccd1 _11796_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _10610_/A _10610_/B _10627_/X vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10678_ _11029_/A2 _10796_/B hold308/A vssd1 vssd1 vccd1 vccd1 _10678_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12417_ _12417_/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12417_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06951__C _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ hold307/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ _12374_/D _12279_/B _12279_/C _12279_/D vssd1 vssd1 vccd1 vccd1 _12280_/C
+ sky130_fd_sc_hd__and4_1
X_06840_ _11611_/A _11607_/B _06839_/X vssd1 vssd1 vccd1 vccd1 _06840_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_65_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06771_ reg1_val[5] _06952_/C vssd1 vssd1 vccd1 vccd1 _06774_/B sky130_fd_sc_hd__and2_1
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09490_ _09490_/A _09490_/B vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__nand2_1
X_08510_ _08510_/A _08510_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09071__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08441_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08372_ _08385_/B _08385_/A vssd1 vssd1 vccd1 vccd1 _08372_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11063__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07323_ _10234_/A _07323_/B vssd1 vssd1 vccd1 vccd1 _07325_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08464__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout137_A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07254_ _07255_/A _07255_/B vssd1 vssd1 vccd1 vccd1 _07254_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07019__A1 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07019__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07185_ reg1_val[14] reg1_val[15] _07121_/C _07089_/C _07093_/A vssd1 vssd1 vccd1
+ vccd1 _07208_/B sky130_fd_sc_hd__o41a_2
XANTENNA__10023__B1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09964__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__B1 _11770_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _07814_/B _11083_/A _10966_/A fanout45/X vssd1 vssd1 vccd1 vccd1 _09827_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06969_ _06967_/A _06967_/B _07026_/C _07074_/B vssd1 vssd1 vccd1 vccd1 _06971_/B
+ sky130_fd_sc_hd__a31o_2
X_09757_ _12490_/S _09753_/X _09754_/X _09756_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__07742__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ _09553_/B _08708_/B vssd1 vssd1 vccd1 vccd1 _09714_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _09701_/A sky130_fd_sc_hd__xor2_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08639_ _12619_/A _07146_/Y _07153_/Y _08605_/A vssd1 vssd1 vccd1 vccd1 _08640_/B
+ sky130_fd_sc_hd__a22o_1
X_11650_ _11980_/A fanout22/X fanout14/X fanout57/X vssd1 vssd1 vccd1 vccd1 _11651_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 fanout31/X vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__or2_1
Xfanout63 _06994_/Y vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__buf_4
X_10601_ _10601_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__xnor2_2
Xfanout74 _07252_/X vssd1 vssd1 vccd1 vccd1 fanout74/X sky130_fd_sc_hd__buf_8
XANTENNA__12251__A1 _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout41 _07139_/X vssd1 vssd1 vccd1 vccd1 fanout41/X sky130_fd_sc_hd__buf_6
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout52 _07052_/Y vssd1 vssd1 vccd1 vccd1 fanout52/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout85 _08400_/B vssd1 vssd1 vccd1 vccd1 fanout85/X sky130_fd_sc_hd__buf_6
Xfanout96 _09827_/A vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__clkbuf_8
X_13320_ _13323_/CLK _13320_/D vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
X_10532_ _10270_/A _10769_/A _10530_/Y vssd1 vssd1 vccd1 vccd1 _10532_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08325__A _08328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13251_ _13350_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
X_10463_ _10463_/A1 fanout11/X fanout7/X _10463_/B2 vssd1 vssd1 vccd1 vccd1 _10464_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13182_ hold299/X _13209_/A2 _13181_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold300/A
+ sky130_fd_sc_hd__a22o_1
X_12202_ _12202_/A _12202_/B _12404_/B _12202_/D vssd1 vssd1 vccd1 vccd1 _12202_/X
+ sky130_fd_sc_hd__or4_1
X_10394_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11357__A3 _11451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06769__B1 _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ _07138_/X wire8/X _12132_/Y _12193_/A vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__a22o_1
X_12064_ _12065_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12138_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11015_ _11014_/A _11014_/B _11014_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _11015_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap102_A _07067_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__B1 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _12978_/A hold248/X vssd1 vssd1 vccd1 vccd1 _13281_/D sky130_fd_sc_hd__and2_1
XANTENNA__09486__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ _11916_/Y _11917_/B _11917_/C vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__and3b_1
X_12897_ hold41/X hold293/X vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11850_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07123__B _07342_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08446__B1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _06683_/C _06840_/Y _06842_/Y vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09946__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _11155_/A _08990_/B vssd1 vssd1 vccd1 vccd1 _08996_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07941_ _07941_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07185__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07873_/C sky130_fd_sc_hd__or2_1
X_06823_ _07179_/A reg1_val[11] vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__and2b_1
X_09611_ _09766_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__xor2_1
X_06754_ _06752_/Y _06754_/B vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__nand2b_1
X_09542_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__and2_1
XANTENNA__07314__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ instruction[29] _06699_/B vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__and2_4
X_09473_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09505_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _08424_/A _08424_/B _08425_/B vssd1 vssd1 vccd1 vccd1 _08424_/X sky130_fd_sc_hd__or3_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07968__B _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08355_ _08566_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08361_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12784__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _09668_/A _07306_/B vssd1 vssd1 vccd1 vccd1 _07308_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10795__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08286_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08286_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07237_ _07074_/A _07073_/X _07074_/Y _06959_/Y vssd1 vssd1 vccd1 vccd1 _07237_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09937__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ reg1_val[16] _07168_/B vssd1 vssd1 vccd1 vccd1 _07180_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07099_ _07299_/B _07113_/A _07113_/B _06811_/B vssd1 vssd1 vccd1 vccd1 _07101_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout231 _12393_/B1 vssd1 vssd1 vccd1 vccd1 _12175_/C1 sky130_fd_sc_hd__buf_4
Xfanout220 _07097_/C vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__clkbuf_8
Xfanout264 _12616_/A vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__buf_8
Xfanout253 _06631_/A vssd1 vssd1 vccd1 vccd1 _06706_/A sky130_fd_sc_hd__buf_4
Xfanout242 _12396_/A vssd1 vssd1 vccd1 vccd1 _06940_/B sky130_fd_sc_hd__buf_4
XANTENNA__07176__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _12978_/A vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__clkbuf_4
Xfanout286 _06569_/Y vssd1 vssd1 vccd1 vccd1 _12378_/S sky130_fd_sc_hd__clkbuf_8
X_09809_ _09810_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09704__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _07077_/X _12782_/Y hold51/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__o211a_1
XANTENNA__11251__A1_N _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09468__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ reg1_val[27] _12773_/A vssd1 vssd1 vccd1 vccd1 _12757_/C sky130_fd_sc_hd__xnor2_2
X_11702_ _11702_/A _11702_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__xnor2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A _12682_/B _12682_/C vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ curr_PC[19] _11718_/C _12525_/S vssd1 vssd1 vccd1 vccd1 _11633_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ _11645_/B _11564_/B vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13303_ _13372_/CLK _13303_/D vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dfxtp_1
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10517_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13234_ hold154/X _12780_/B _12777_/Y _12781_/A vssd1 vssd1 vccd1 vccd1 _13236_/B
+ sky130_fd_sc_hd__a22o_1
X_10446_ _12202_/B _08274_/B fanout74/X _12202_/A vssd1 vssd1 vccd1 vccd1 _10447_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _12865_/X _13165_/B vssd1 vssd1 vccd1 vccd1 _13166_/B sky130_fd_sc_hd__nand2b_1
X_10377_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__and2_1
X_12116_ _09225_/X _12115_/X _06635_/B vssd1 vssd1 vccd1 vccd1 _12116_/X sky130_fd_sc_hd__a21o_1
X_13096_ _13109_/A hold272/X vssd1 vssd1 vccd1 vccd1 _13341_/D sky130_fd_sc_hd__and2_1
X_12047_ _12041_/Y _12042_/X _12046_/Y _12039_/X vssd1 vssd1 vccd1 vccd1 _12047_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_46_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09614__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__A1 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__B2 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__B _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ hold62/X _12948_/B hold279/X vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06973__A _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06692__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _08140_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ _08071_/A _08170_/A vssd1 vssd1 vccd1 vccd1 _08104_/A sky130_fd_sc_hd__or2_1
XFILLER_0_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ _07389_/A _07389_/B _07003_/X vssd1 vssd1 vccd1 vccd1 _07082_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_113_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11726__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08973_ _12335_/A _08971_/X _06644_/X vssd1 vssd1 vccd1 vccd1 fanout7/A sky130_fd_sc_hd__a21o_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07924_ _07922_/A _07922_/B _07999_/A vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__a21bo_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07855_ _07852_/A _07852_/B _07936_/A vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09243__B _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ _06793_/Y _06804_/X _06805_/X vssd1 vssd1 vccd1 vccd1 _09739_/B sky130_fd_sc_hd__a21oi_1
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__xnor2_4
X_06737_ reg1_val[11] _07179_/A vssd1 vssd1 vccd1 vccd1 _06738_/B sky130_fd_sc_hd__nor2_1
X_09525_ _09525_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__nor2_2
X_06668_ reg1_val[22] _06993_/A vssd1 vssd1 vccd1 vccd1 _06669_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10465__B1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09458_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08122__A2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__A2 _11041_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ _08624_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06599_ instruction[24] _06591_/X _06908_/B instruction[41] _06595_/X vssd1 vssd1
+ vccd1 vccd1 _06600_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09387_ _09385_/X _09386_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08338_ _08338_/A _08338_/B vssd1 vssd1 vccd1 vccd1 _08392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08308_/B sky130_fd_sc_hd__xnor2_1
X_11280_ _11645_/A fanout22/X fanout14/X fanout51/X vssd1 vssd1 vccd1 vccd1 _11281_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nand2_1
X_10231_ _10231_/A _10231_/B _10231_/C vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08189__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13182__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__B _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _10029_/A _10026_/Y _10028_/B vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_30_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10940__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10094_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ hold38/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__or2_1
XANTENNA__11248__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _11107_/B sky130_fd_sc_hd__or2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ reg1_val[24] _12773_/A vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ reg1_val[10] _12666_/B vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12596_ reg1_val[24] curr_PC[24] _12615_/S vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__mux2_2
X_11616_ _11520_/B _11522_/B _11520_/A vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09613__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12748__A2 _07342_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09074__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _12065_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11548_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_92_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _12068_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13217_ hold307/A _13216_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13173__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ hold313/A _10558_/C vssd1 vssd1 vccd1 vccd1 _10429_/X sky130_fd_sc_hd__or2_1
X_13148_ hold311/X _13186_/A2 _13147_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold312/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__A _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ hold273/X hold3/X fanout3/X vssd1 vssd1 vccd1 vccd1 _13079_/Y sky130_fd_sc_hd__nand3_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ _07640_/A _07640_/B vssd1 vssd1 vccd1 vccd1 _07642_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07571_ reg1_val[29] _07572_/B vssd1 vssd1 vccd1 vccd1 _11813_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07560__B1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ _09787_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09241_ hold321/A _09237_/Y _09239_/Y _13338_/Q _09236_/X vssd1 vssd1 vccd1 vccd1
+ _09242_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09172_ reg1_val[10] reg1_val[21] _09180_/S vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08123_ _08573_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _08202_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07615__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07615__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ _08054_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07005_ reg1_val[2] _07005_/B vssd1 vssd1 vccd1 vccd1 _07009_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08591__A2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _08955_/B _08956_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__and2b_1
X_07907_ _08445_/A _07907_/B vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__xnor2_1
X_08887_ _08888_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__and2_1
X_07838_ _07834_/A _07834_/B _07872_/A vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _08096_/B _11296_/A _11188_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _09509_/B
+ sky130_fd_sc_hd__o22a_1
X_07769_ _10067_/A1 _08400_/B fanout82/X _08926_/B1 vssd1 vssd1 vccd1 vccd1 _07770_/B
+ sky130_fd_sc_hd__o22a_1
X_10780_ _10779_/A _10779_/B _10779_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _10780_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07303__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout32_A _07181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09439_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12627_/B _12450_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07606__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12381_/A _12381_/B vssd1 vssd1 vccd1 vccd1 _12381_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07606__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ _11781_/S _06832_/Y _11331_/Y vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _07031_/X fanout29/X _07301_/Y fanout31/X vssd1 vssd1 vccd1 vccd1 _11264_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11166__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11166__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ _13134_/A hold229/X vssd1 vssd1 vccd1 vccd1 _13299_/D sky130_fd_sc_hd__and2_1
X_10214_ _10213_/A _11645_/B _10213_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07909__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10913__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _11021_/S _09398_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _10145_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10076_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12969__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08508__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12717_ _12767_/B _12717_/B vssd1 vssd1 vccd1 vccd1 _12719_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12648_ _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12649_/B sky130_fd_sc_hd__or2_2
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ reg1_val[21] curr_PC[21] _12615_/S vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08810_ _07658_/A _07658_/B _07656_/X vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__a21oi_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10380__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _09791_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__or2_1
XANTENNA__07781__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08739_/X _08740_/Y _08737_/Y vssd1 vssd1 vccd1 vccd1 _08741_/X sky130_fd_sc_hd__a21o_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _08672_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09802__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07623_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__or2_1
XFILLER_0_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout167_A _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09286__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _07663_/B _07663_/A vssd1 vssd1 vccd1 vccd1 _07554_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11632__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07485_ _07486_/A _07486_/B vssd1 vssd1 vccd1 vccd1 _07485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ _09238_/B _09229_/B vssd1 vssd1 vccd1 vccd1 _09595_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09155_ _09219_/A reg1_val[31] _09155_/S vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08106_ _08106_/A _08106_/B vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__xor2_1
X_09086_ _09087_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__or2_1
XANTENNA__13275__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08037_ _09795_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09988_ _09989_/B _09989_/A vssd1 vssd1 vccd1 vccd1 _09988_/Y sky130_fd_sc_hd__nand2b_1
X_08939_ _08938_/B _08939_/B vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ _11947_/X _11948_/Y _11949_/X _12378_/S vssd1 vssd1 vccd1 vccd1 _11951_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08316__A2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ _06879_/D _10899_/Y _10900_/Y vssd1 vssd1 vccd1 vccd1 _10901_/X sky130_fd_sc_hd__a21o_1
X_11881_ _11529_/B _11960_/B hold199/A vssd1 vssd1 vccd1 vccd1 _11881_/Y sky130_fd_sc_hd__a21oi_1
X_10832_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08328__A _08328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__A1 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ _10764_/A _10764_/B _10764_/C vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12503_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _10694_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10696_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12284__S _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _12433_/A1 _12425_/Y _12432_/X _12423_/Y vssd1 vssd1 vccd1 vccd1 _12433_/X
+ sky130_fd_sc_hd__o211a_1
X_12364_ _12364_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__or2_1
X_11315_ _11316_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11411_/B sky130_fd_sc_hd__or2_1
XANTENNA__13128__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ hold251/A _12347_/B _12345_/B _12433_/A1 vssd1 vssd1 vccd1 vccd1 _12295_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09201__A0 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ _09886_/B _12394_/A1 _11246_/S vssd1 vssd1 vccd1 vccd1 _11246_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _11359_/A _11177_/B vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09752__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _10128_/A _10267_/A _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10129_/C
+ sky130_fd_sc_hd__or4_2
X_10059_ _10233_/A1 fanout13/X fanout11/X _10233_/B2 vssd1 vssd1 vccd1 vccd1 _10060_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06965__B _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13144__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09807__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ _09795_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07358_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06981__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09069__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _11052_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__xnor2_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_09842_ _09621_/A _09621_/B _09620_/A vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__a21o_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10353__A2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09775_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07317__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout284_A _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ _09668_/A vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__inv_4
X_08724_ _08723_/A _08723_/B _08721_/B _08721_/A vssd1 vssd1 vccd1 vccd1 _10656_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06875__B _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _08655_/A _09430_/A vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__or2_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ fanout60/X _10233_/B2 _10233_/A1 fanout52/X vssd1 vssd1 vccd1 vccd1 _07607_/B
+ sky130_fd_sc_hd__o22a_1
X_08586_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08588_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_49_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ fanout45/X _09324_/A _08591_/B1 _07814_/B vssd1 vssd1 vccd1 vccd1 _07538_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12802__A1 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07468_ _08648_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07285__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ reg1_val[11] reg1_val[20] _09560_/A vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__mux2_1
X_07399_ _07399_/A _07399_/B vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07198__S _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _09139_/B _09139_/A vssd1 vssd1 vccd1 vccd1 _09138_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10041__A1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11100_ _11101_/B _11101_/A vssd1 vssd1 vccd1 vccd1 _11100_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _10231_/A _09069_/B vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12080_ _12080_/A _12080_/B _12080_/C vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11031_ _12395_/A1 _11030_/X _06727_/B vssd1 vssd1 vccd1 vccd1 _11031_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07227__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12982_ _13144_/A hold211/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__and2_1
XANTENNA__12787__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__B1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _11933_/A _11933_/B _11933_/C vssd1 vssd1 vccd1 vccd1 _11934_/A sky130_fd_sc_hd__and3_1
XANTENNA__10588__A _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__A1 _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ _11864_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11864_/Y sky130_fd_sc_hd__xnor2_2
X_10815_ _10702_/A _10702_/B _10707_/A vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__a21o_1
X_11795_ _11529_/B _11880_/B hold249/A vssd1 vssd1 vccd1 vccd1 _11795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10746_ _10746_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__and2_1
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10677_ hold303/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10796_/B sky130_fd_sc_hd__or2_1
XANTENNA__12308__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ _12335_/A _06871_/X _12381_/X _12415_/Y vssd1 vssd1 vccd1 vccd1 _12417_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06951__D _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09422__B1 _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B2 _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__A1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12347_ hold253/A _12347_/B _12387_/B vssd1 vssd1 vccd1 vccd1 _12347_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _12278_/A _12278_/B _12279_/C _12279_/D vssd1 vssd1 vccd1 vccd1 _12330_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13139__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _11228_/A _11228_/B _11228_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _11253_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12978__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ reg1_val[5] _06952_/C vssd1 vssd1 vccd1 vccd1 _06774_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10498__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06695__B _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08440_ _08440_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08441_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08397_/A _08369_/Y _08366_/Y vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ fanout52/X _10233_/B2 _10233_/A1 fanout50/X vssd1 vssd1 vccd1 vccd1 _07323_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08464__A1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08464__B2 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07253_ _07175_/A _07299_/B _07175_/B vssd1 vssd1 vccd1 vccd1 _07255_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07019__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ _11361_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09964__A1 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09964__B2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07047__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _09609_/Y _09612_/B _09617_/A vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__a21o_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06968_ _06978_/A _06975_/A vssd1 vssd1 vccd1 vccd1 _07026_/C sky130_fd_sc_hd__and2_1
X_09756_ _12490_/S _10035_/C vssd1 vssd1 vccd1 vccd1 _09756_/Y sky130_fd_sc_hd__nor2_1
X_09687_ _09685_/Y _09687_/B vssd1 vssd1 vccd1 vccd1 _09688_/B sky130_fd_sc_hd__and2b_1
X_08707_ _08707_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__and2_1
X_06899_ _06767_/A _06593_/X _09240_/B instruction[4] _06897_/Y vssd1 vssd1 vccd1
+ vccd1 _12782_/B sky130_fd_sc_hd__a221oi_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08638_ _08638_/A _08638_/B _08638_/C vssd1 vssd1 vccd1 vccd1 _08663_/B sky130_fd_sc_hd__and3_1
XFILLER_0_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout31 _07193_/Y vssd1 vssd1 vccd1 vccd1 fanout31/X sky130_fd_sc_hd__clkbuf_8
Xfanout20 _08985_/Y vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__buf_8
X_08569_ _08619_/B2 _09468_/B2 _08591_/B1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08570_/B
+ sky130_fd_sc_hd__o22a_1
X_11580_ _11490_/A _11490_/B _11488_/X vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__a21boi_1
Xfanout53 _07052_/Y vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__buf_4
X_10600_ _10601_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10600_/Y sky130_fd_sc_hd__nand2_1
Xfanout42 _07402_/B vssd1 vssd1 vccd1 vccd1 fanout42/X sky130_fd_sc_hd__clkbuf_8
Xfanout64 _06977_/Y vssd1 vssd1 vccd1 vccd1 fanout64/X sky130_fd_sc_hd__buf_8
XFILLER_0_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout9_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout86 _07236_/Y vssd1 vssd1 vccd1 vccd1 _08400_/B sky130_fd_sc_hd__buf_8
Xfanout97 _07096_/X vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__buf_12
X_10531_ _10650_/B _10650_/C vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__nor2_2
XANTENNA__09201__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout75 _11083_/A vssd1 vssd1 vccd1 vccd1 fanout75/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07510__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ _13346_/CLK hold17/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12539__A0 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10462_ _10382_/A _10382_/B _10379_/A vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__a21oi_2
X_12201_ _12202_/A _12202_/D _12202_/B vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13181_ hold302/A _13180_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__mux2_1
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _12132_/A wire8/X vssd1 vssd1 vccd1 vccd1 _12132_/Y sky130_fd_sc_hd__nand2_1
X_12063_ _12310_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__xnor2_1
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12965_ hold232/X _13095_/B2 _13158_/A2 hold247/X vssd1 vssd1 vccd1 vccd1 hold248/A
+ sky130_fd_sc_hd__a22o_1
X_11916_ _12310_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__xnor2_1
X_12896_ _12881_/B _13101_/B _12879_/X vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__a21o_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11777_/A _11777_/B _11946_/A vssd1 vssd1 vccd1 vccd1 _11778_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08446__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08446__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10729_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10745_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ instruction[14] vssd1 vssd1 vccd1 vccd1 loadstore_dest[3] sky130_fd_sc_hd__buf_12
XANTENNA__09946__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13375_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10556__A2 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07709__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _07837_/B _07871_/B vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__and2b_1
X_06822_ _10660_/A _06820_/Y _06821_/X vssd1 vssd1 vccd1 vccd1 _06822_/X sky130_fd_sc_hd__o21ba_1
X_09610_ _07539_/B _10712_/A _07212_/X fanout37/X vssd1 vssd1 vccd1 vccd1 _09611_/B
+ sky130_fd_sc_hd__a22o_1
X_06753_ reg1_val[8] _07195_/A vssd1 vssd1 vccd1 vccd1 _06754_/B sky130_fd_sc_hd__nand2_1
X_09541_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06684_ _06884_/B vssd1 vssd1 vccd1 vccd1 _06684_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09882__B1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _09470_/X _09472_/B vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08423_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout247_A _06893_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ _06875_/A _08354_/A2 _10585_/B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08355_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08988__A2 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07330__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07305_ _08633_/B fanout58/X fanout56/X _09300_/A vssd1 vssd1 vccd1 vccd1 _07306_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08285_ _08335_/A _08335_/B _08281_/X vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _07236_/A _07236_/B vssd1 vssd1 vccd1 vccd1 _07236_/Y sky130_fd_sc_hd__nand2_1
X_07167_ _11231_/A _07167_/B vssd1 vssd1 vccd1 vccd1 _07167_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__09937__B2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__A1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07948__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _11237_/S _06950_/X _06949_/Y _06952_/C vssd1 vssd1 vccd1 vccd1 _07101_/A
+ sky130_fd_sc_hd__a211o_1
Xfanout232 _09240_/X vssd1 vssd1 vccd1 vccd1 _12393_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout221 _07097_/C vssd1 vssd1 vccd1 vccd1 _10288_/S sky130_fd_sc_hd__clkbuf_4
Xfanout210 _09101_/A vssd1 vssd1 vccd1 vccd1 _12785_/A sky130_fd_sc_hd__buf_6
Xfanout265 _06591_/X vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__buf_4
Xfanout254 _13071_/A2 vssd1 vssd1 vccd1 vccd1 _13055_/A2 sky130_fd_sc_hd__buf_4
Xfanout243 _12525_/S vssd1 vssd1 vccd1 vccd1 _12490_/S sky130_fd_sc_hd__buf_6
Xfanout276 _13219_/A vssd1 vssd1 vccd1 vccd1 _13187_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10180__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _09301_/A _06991_/A fanout7/X _09807_/Y vssd1 vssd1 vccd1 vccd1 _09810_/B
+ sky130_fd_sc_hd__o31ai_2
Xfanout287 _06566_/Y vssd1 vssd1 vccd1 vccd1 _06875_/A sky130_fd_sc_hd__buf_6
XANTENNA__08373__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout62_A _06994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ _12415_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09739_/X sky130_fd_sc_hd__and2_1
XANTENNA__07505__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12750_ _12746_/B _12749_/B _12744_/X vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__a21o_1
X_11701_ _11615_/B _11617_/B _11615_/A vssd1 vssd1 vccd1 vccd1 _11702_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12682_/A _12682_/B _12682_/C vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__a21o_1
X_11632_ _07058_/A _11446_/B _06941_/X _11631_/X vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ fanout61/X fanout9/X fanout4/X _11645_/A vssd1 vssd1 vccd1 vccd1 _11564_/B
+ sky130_fd_sc_hd__o22a_1
X_13302_ _13372_/CLK _13302_/D vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11494_/A _11494_/B vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10514_ _10458_/B _10333_/B _10357_/B _10356_/B _10356_/A vssd1 vssd1 vccd1 vccd1
+ _10517_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _13236_/A _13233_/B hold203/X vssd1 vssd1 vccd1 vccd1 _13372_/D sky130_fd_sc_hd__and3_1
X_10445_ _10345_/A _10345_/B _10343_/Y vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13164_ _13187_/A hold282/X vssd1 vssd1 vccd1 vccd1 _13355_/D sky130_fd_sc_hd__and2_1
XFILLER_0_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10376_ _11359_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10378_/B sky130_fd_sc_hd__xnor2_1
X_12115_ _12431_/A2 _09235_/X _12115_/S vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__mux2_1
X_13095_ hold271/X _13222_/A2 _13094_/X _13095_/B2 vssd1 vssd1 vccd1 vccd1 hold272/A
+ sky130_fd_sc_hd__a22o_1
X_12046_ _09155_/S _10288_/X _12045_/X vssd1 vssd1 vccd1 vccd1 _12046_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08364__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__C _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ hold62/X _12948_/B vssd1 vssd1 vccd1 vccd1 _12950_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12879_ hold21/X hold317/A vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09630__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06973__B _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _08071_/A _08070_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07021_ _07021_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07389_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11726__B2 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _12335_/A _08971_/X _06644_/X vssd1 vssd1 vccd1 vccd1 wire8/A sky130_fd_sc_hd__a21oi_2
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _07998_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07854_ _07935_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__nor2_1
X_06805_ reg1_val[2] _10286_/S vssd1 vssd1 vccd1 vccd1 _06805_/X sky130_fd_sc_hd__and2_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08107__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _07853_/A _07853_/B _07778_/X vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__a21o_2
X_06736_ reg1_val[11] _07179_/A vssd1 vssd1 vccd1 vccd1 _10794_/S sky130_fd_sc_hd__and2_1
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__nor2_1
X_06667_ reg1_val[22] _06993_/A vssd1 vssd1 vccd1 vccd1 _11883_/S sky130_fd_sc_hd__and2_1
XANTENNA__10465__A1 _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ _09283_/A _09283_/B _09284_/X vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08406_ _08641_/A2 _08521_/A2 _08926_/B1 _08649_/B vssd1 vssd1 vccd1 vccd1 _08407_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06598_ instruction[41] _06908_/B _06595_/X vssd1 vssd1 vccd1 vccd1 _06631_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__07060__A _07060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ _09173_/X _09176_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08337_ _08337_/A _08337_/B vssd1 vssd1 vccd1 vccd1 _08392_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ _08268_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _08096_/B _10589_/A fanout24/X _08926_/B1 vssd1 vssd1 vccd1 vccd1 _07220_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__11717__A1 _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _10230_/A _10230_/B _10230_/C vssd1 vssd1 vccd1 vccd1 _10231_/C sky130_fd_sc_hd__nand3_1
X_08199_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08594__B1 _07043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _10143_/A _09228_/Y _11966_/B _06765_/B _10160_/X vssd1 vssd1 vccd1 vccd1
+ _10161_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10940__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__and2_1
XANTENNA__12142__A1 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__B2 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _10876_/A _10876_/B _10877_/Y vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__o21a_1
X_12802_ _10326_/A _13072_/A2 hold16/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold17/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12795__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12733_/A _12737_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12664_/A _12664_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
X_12595_ _12598_/D _12595_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
X_11615_ _11615_/A _11615_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09074__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09074__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ _07031_/X _07151_/A _07155_/A _12143_/A vssd1 vssd1 vccd1 vccd1 _11547_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08821__B2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13216_ _13216_/A _13216_/B vssd1 vssd1 vccd1 vccd1 _13216_/Y sky130_fd_sc_hd__xnor2_1
X_11477_ _07012_/Y fanout42/X fanout40/X _11917_/B vssd1 vssd1 vccd1 vccd1 _11478_/B
+ sky130_fd_sc_hd__a22o_1
X_10428_ _06754_/B _09228_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _10428_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ hold319/A _13146_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
X_10359_ _08400_/B _10466_/B _10466_/C fanout82/X _12202_/B vssd1 vssd1 vccd1 vccd1
+ _10360_/B sky130_fd_sc_hd__o32a_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ hold273/X _13227_/B _11645_/B _13078_/B2 hold7/X vssd1 vssd1 vccd1 vccd1
+ hold8/A sky130_fd_sc_hd__o221a_1
XFILLER_0_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12133__B2 _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12029_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _12029_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10144__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__A _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ reg1_val[28] _08868_/C _12756_/B _07229_/B vssd1 vssd1 vccd1 vccd1 _07572_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__07560__B2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _09240_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09240_/X sky130_fd_sc_hd__or2_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _09169_/X _09170_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _08594_/A2 _10585_/B2 _10067_/A1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08123_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07615__A2 _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08053_ _08052_/A _08063_/A vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ _12619_/A reg1_val[1] _07093_/A vssd1 vssd1 vccd1 vccd1 _07005_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ _08956_/B _08955_/B vssd1 vssd1 vccd1 vccd1 _09064_/B sky130_fd_sc_hd__and2b_1
X_07906_ _10067_/A1 _10227_/B1 _10463_/A1 _09114_/B1 vssd1 vssd1 vccd1 vccd1 _07907_/B
+ sky130_fd_sc_hd__o22a_1
X_08886_ _09630_/A _08886_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__xnor2_1
X_07837_ _07871_/B _07837_/B vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__and2b_1
X_07768_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06719_ _11125_/A _07251_/A vssd1 vssd1 vccd1 vccd1 _06721_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09828__B1 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _09507_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_94_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08500__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07303__B2 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07303__A1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _10081_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07701_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout25_A _07215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__nand3_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ _09370_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11307_/A _11307_/B _11306_/A vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11938__A1 _11770_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _12381_/A _12379_/B _11612_/A vssd1 vssd1 vccd1 vccd1 _12380_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07606__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11781_/S _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _11900_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__xnor2_1
X_11193_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11166__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ hold228/X _13143_/B2 _13209_/A2 hold188/X vssd1 vssd1 vccd1 vccd1 hold229/A
+ sky130_fd_sc_hd__a22o_1
X_10213_ _10213_/A _11645_/B _10213_/C vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__and3_1
XANTENNA__11975__A _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__B1 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10143_/A _10143_/B _09226_/Y vssd1 vssd1 vccd1 vccd1 _10144_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11626__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10977_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12716_ _12716_/A _12716_/B _12716_/C _12716_/D vssd1 vssd1 vccd1 vccd1 _12719_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12647_ reg1_val[6] _12647_/B vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__and2_1
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _12588_/A _12578_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XANTENNA__10773__B _10810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08524__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
X_11529_ hold255/A _11529_/B _11620_/B vssd1 vssd1 vccd1 vccd1 _11529_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12354__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__A1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08740_ _08746_/B _08746_/C _08746_/D vssd1 vssd1 vccd1 vccd1 _08740_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__07781__B2 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08671_ _08670_/A _08670_/B _08670_/C _08672_/B _08581_/X vssd1 vssd1 vccd1 vccd1
+ _08673_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13067__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09286__B2 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _07553_/A _07553_/B vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11125__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ _07387_/A _07387_/B _07386_/A vssd1 vssd1 vccd1 vccd1 _07486_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09223_ _11781_/S _09223_/B vssd1 vssd1 vccd1 vccd1 _09223_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07049__B1 _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _12621_/A reg1_val[30] _09180_/S vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08434__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09085_ _11168_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _09087_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08036_ _08619_/B1 _08096_/B fanout24/X _09403_/S vssd1 vssd1 vccd1 vccd1 _08037_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09265__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__xnor2_1
X_08938_ _08939_/B _08938_/B vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ reg1_val[28] reg1_val[29] _08868_/C _12756_/B _07229_/B vssd1 vssd1 vccd1
+ vccd1 _08870_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _06879_/D _10899_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _10900_/Y sky130_fd_sc_hd__o21ai_1
X_11880_ hold249/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__or2_1
XANTENNA__09204__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__and2_1
XANTENNA__13073__A2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ _10764_/A _10764_/B _10764_/C vssd1 vssd1 vccd1 vccd1 _10765_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12820__A2 _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__a21o_1
X_10693_ _10694_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10870_/A sky130_fd_sc_hd__or2_1
X_12432_ _09196_/S _09217_/Y _12428_/X _12431_/X vssd1 vssd1 vccd1 vccd1 _12432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12364_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11314_ _11205_/A _11205_/B _11206_/Y vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _12347_/B _12345_/B hold251/A vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__a21oi_1
X_11245_ hold331/A _11879_/A2 _11341_/B _11244_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _11249_/B sky130_fd_sc_hd__a311o_1
XANTENNA__12336__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08004__A2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _07031_/X fanout31/X fanout29/X _12143_/A vssd1 vssd1 vccd1 vccd1 _11177_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09752__A2 _09728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10650_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08960__B1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10058_ _10058_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13064__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06981__B _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ fanout46/X _11188_/A _11083_/A fanout44/X vssd1 vssd1 vccd1 vccd1 _09911_/B
+ sky130_fd_sc_hd__o22a_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ _09688_/A _09687_/B _09685_/Y vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__a21o_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _12193_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__xor2_1
X_06984_ reg1_val[5] _06984_/B vssd1 vssd1 vccd1 vccd1 _06984_/Y sky130_fd_sc_hd__xnor2_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08723_/A _08723_/B vssd1 vssd1 vccd1 vccd1 _10541_/C sky130_fd_sc_hd__or2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08654_ _08476_/A _08605_/A _07128_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _09430_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ _07605_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__xor2_1
X_08585_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07536_ _08476_/A _07539_/B vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12802__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__A _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _09202_/X _09205_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__mux2_1
X_07467_ _06973_/A fanout58/X fanout56/X _06973_/Y vssd1 vssd1 vccd1 vccd1 _07468_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07398_ _07398_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07399_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ _09137_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09139_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ fanout67/X _08590_/B _09648_/A fanout64/X vssd1 vssd1 vccd1 vccd1 _09069_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08019_ _10468_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout92_A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A0 _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _09886_/B _12394_/A1 _11030_/S vssd1 vssd1 vccd1 vccd1 _11030_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11972__B _11972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ hold234/A _13143_/B2 _13186_/A2 hold210/X vssd1 vssd1 vccd1 vccd1 hold211/A
+ sky130_fd_sc_hd__a22o_1
X_11932_ _11933_/A _11933_/B _11933_/C vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10588__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07243__A _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _11863_/A _11863_/B vssd1 vssd1 vccd1 vccd1 _11864_/B sky130_fd_sc_hd__nand2_1
X_10814_ _10713_/A _10713_/B _10714_/Y vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11794_ hold225/A _11794_/B vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__or2_1
XANTENNA__10804__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _10745_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ _12395_/A1 _10675_/X _06743_/A vssd1 vssd1 vccd1 vccd1 _10676_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08074__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12415_ _12415_/A _12415_/B vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ _12347_/B _12387_/B hold253/A vssd1 vssd1 vccd1 vccd1 _12346_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12277_ _12280_/B vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__inv_2
XANTENNA__10543__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11228_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11228_/Y sky130_fd_sc_hd__nand2_1
X_11159_ _11158_/B _11159_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07200__A3 _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08370_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12796__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ _07321_/A _07321_/B vssd1 vssd1 vccd1 vccd1 _07325_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12260__A3 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08464__A2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _11070_/A _11071_/A _11169_/A vssd1 vssd1 vccd1 vccd1 _07252_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09413__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07183_ _07171_/X _10222_/A2 _10712_/A _07182_/Y vssd1 vssd1 vccd1 vccd1 _07184_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10023__A2 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09964__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10731__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ _06967_/A _06967_/B vssd1 vssd1 vccd1 vccd1 _06967_/Y sky130_fd_sc_hd__nand2_1
X_09755_ curr_PC[0] curr_PC[1] curr_PC[2] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _10035_/C
+ sky130_fd_sc_hd__and4_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ instruction[5] instruction[6] vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__nand2b_4
X_09686_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__nand2_1
X_08706_ _09670_/A _09553_/B _08656_/B vssd1 vssd1 vccd1 vccd1 _08707_/B sky130_fd_sc_hd__o21ai_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08637_ _08638_/A _08638_/C _08638_/B vssd1 vssd1 vccd1 vccd1 _08637_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout10 _08874_/Y vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__clkbuf_8
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 _11917_/C vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__buf_8
X_08568_ _08650_/A _08568_/B vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__xnor2_2
Xfanout65 _06977_/Y vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__buf_4
XFILLER_0_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout54 fanout55/X vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__clkbuf_8
Xfanout43 _07137_/Y vssd1 vssd1 vccd1 vccd1 _07402_/B sky130_fd_sc_hd__buf_6
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout32 _07181_/X vssd1 vssd1 vccd1 vccd1 fanout32/X sky130_fd_sc_hd__buf_8
X_07519_ _07519_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__nor2_1
X_08499_ _08499_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout87 _11054_/A vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__buf_12
X_10530_ _10263_/X _10403_/X _10404_/X vssd1 vssd1 vccd1 vccd1 _10530_/Y sky130_fd_sc_hd__a21oi_2
Xfanout98 _11386_/A vssd1 vssd1 vccd1 vccd1 fanout98/X sky130_fd_sc_hd__buf_8
Xfanout76 _07251_/Y vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10509_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13200__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12255_/B _12205_/B vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _13180_/A _13180_/B vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10392_ _10390_/A _10390_/B _10393_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12134_/B sky130_fd_sc_hd__xnor2_1
X_12062_ _12257_/A fanout14/X _12309_/A fanout22/X vssd1 vssd1 vccd1 vccd1 _12063_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12172__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _06826_/Y _11012_/X _12025_/S vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10722__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12964_ _12978_/A hold233/X vssd1 vssd1 vccd1 vccd1 _13280_/D sky130_fd_sc_hd__and2_1
X_11915_ _12202_/B fanout22/X fanout14/X _12202_/A vssd1 vssd1 vccd1 vccd1 _11916_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12895_ _12884_/B _13097_/B _12882_/X vssd1 vssd1 vccd1 vccd1 _13101_/B sky130_fd_sc_hd__a21o_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11933_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__and2_1
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11777_/A _11777_/B vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08446__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11450__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10659_ _06820_/Y _10658_/Y _12025_/S vssd1 vssd1 vccd1 vccd1 _10660_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09946__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ instruction[13] vssd1 vssd1 vccd1 vccd1 loadstore_dest[2] sky130_fd_sc_hd__buf_12
XFILLER_0_11_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08532__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _12405_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12374_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10961__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12163__C1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__B2 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A1 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07869_/A _07869_/B _07869_/C vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__a21oi_1
X_06821_ _07213_/A reg1_val[10] vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06752_ reg1_val[8] _07195_/A vssd1 vssd1 vccd1 vccd1 _06752_/Y sky130_fd_sc_hd__nor2_1
X_09540_ _09540_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__xnor2_4
X_09471_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__or3_1
XFILLER_0_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06683_ _11951_/A _11947_/A _06683_/C _11782_/A vssd1 vssd1 vccd1 vccd1 _06884_/B
+ sky130_fd_sc_hd__nor4_1
XANTENNA__09882__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ _08391_/X _08421_/Y _08390_/X vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12229__A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout142_A _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _08353_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07304_ _09670_/A _07304_/B vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__xnor2_2
X_08284_ _08624_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07235_ _10230_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07236_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07166_ reg1_val[14] _07121_/C _07229_/B vssd1 vssd1 vccd1 vccd1 _07167_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09937__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07097_ _12415_/A _07127_/B _07097_/C vssd1 vssd1 vccd1 vccd1 _07113_/B sky130_fd_sc_hd__and3_1
XANTENNA__07948__A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__B2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__A _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 _13209_/A2 vssd1 vssd1 vccd1 vccd1 _13186_/A2 sky130_fd_sc_hd__buf_4
Xfanout222 _06776_/X vssd1 vssd1 vccd1 vccd1 _07097_/C sky130_fd_sc_hd__buf_4
Xfanout211 _09722_/S vssd1 vssd1 vccd1 vccd1 _09724_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout255 _12782_/A vssd1 vssd1 vccd1 vccd1 _13071_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout244 _12504_/S vssd1 vssd1 vccd1 vccd1 _12525_/S sky130_fd_sc_hd__buf_6
Xfanout233 _09232_/Y vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__08373__A1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _13134_/A vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__buf_4
XANTENNA__10180__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ _06991_/B fanout7/X _09301_/A vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__o21ai_1
Xfanout266 _12767_/B vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__buf_8
Xfanout288 _06566_/Y vssd1 vssd1 vccd1 vccd1 _06973_/A sky130_fd_sc_hd__buf_4
XANTENNA__08373__B2 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08057_/A sky130_fd_sc_hd__and2_1
XANTENNA__10180__B2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _10288_/S _09737_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09669_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09669_/Y sky130_fd_sc_hd__nor2_1
X_11700_ _11700_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06823__A_N _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ _12688_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _12682_/C sky130_fd_sc_hd__nand2_1
X_11631_ _11602_/Y _11603_/X _11606_/Y _11946_/A _11630_/X vssd1 vssd1 vccd1 vccd1
+ _11631_/X sky130_fd_sc_hd__o221a_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _11562_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09625__B2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ _13372_/CLK hold244/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__dfxtp_1
X_10513_ _10386_/A _10385_/B _10383_/X vssd1 vssd1 vccd1 vccd1 _10518_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11493_ _11494_/B _11494_/A vssd1 vssd1 vccd1 vccd1 _11493_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11978__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ hold193/X hold149/X hold197/X vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__a21o_1
X_10444_ _10398_/A _10398_/B _10396_/Y vssd1 vssd1 vccd1 vccd1 _10526_/A sky130_fd_sc_hd__a21o_2
X_13163_ hold281/X _06901_/Y _13162_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold282/A
+ sky130_fd_sc_hd__a22o_1
X_10375_ _11734_/A fanout31/X fanout29/X _11568_/A vssd1 vssd1 vccd1 vccd1 _10376_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ hold188/A _12178_/A2 _12176_/B _12113_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12119_/B sky130_fd_sc_hd__a311o_1
XANTENNA__10943__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ hold322/A _13093_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__mux2_1
X_12045_ _06641_/B _06940_/B _09222_/Y _10282_/X _12044_/X vssd1 vssd1 vccd1 vccd1
+ _12045_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08364__A1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__A1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__B2 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__D _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09911__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ _12851_/B _13220_/B _12851_/A vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12878_ hold293/X hold41/X vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08527__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07875__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _11829_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12483__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07020_ _08650_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08971_ _08971_/A _08971_/B _08971_/C _08971_/D vssd1 vssd1 vccd1 vccd1 _08971_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12512__A _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _07922_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07998_/B sky130_fd_sc_hd__xnor2_1
X_07853_ _07853_/A _07853_/B vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__xnor2_1
X_06804_ _09419_/A _09416_/B _06803_/X vssd1 vssd1 vccd1 vccd1 _06804_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09304__B1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__B2 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07853_/B sky130_fd_sc_hd__xnor2_1
X_06735_ _06908_/A _06631_/A _12679_/B _06734_/X vssd1 vssd1 vccd1 vccd1 _07179_/A
+ sky130_fd_sc_hd__a31o_4
X_09523_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__and2_1
X_06666_ _06664_/Y _06600_/Y _06712_/B reg2_val[22] vssd1 vssd1 vccd1 vccd1 _06993_/A
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__10465__A2 _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _09622_/B _09454_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__or2_2
X_09385_ _09170_/X _09172_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__mux2_1
X_08405_ _08566_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08437__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06597_ instruction[41] _06908_/B _06595_/X vssd1 vssd1 vccd1 vccd1 _06767_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07060__B _07060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__A1 _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__B2 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _08336_/A _08336_/B vssd1 vssd1 vccd1 vccd1 _08337_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08267_ _08267_/A _08267_/B vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07218_ _07218_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _07218_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11717__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _07148_/A _07148_/B _07148_/C vssd1 vssd1 vccd1 vccd1 _07150_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08594__A1 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10160_ _07264_/A _06940_/B _09595_/B _06763_/A _10159_/Y vssd1 vssd1 vccd1 vccd1
+ _10160_/X sky130_fd_sc_hd__a221o_1
X_10091_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09207__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _11107_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11980__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ hold15/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ reg1_val[23] _12773_/A vssd1 vssd1 vccd1 vccd1 _12737_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07251__A _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12663_ _12668_/B _12670_/A vssd1 vssd1 vccd1 vccd1 _12664_/B sky130_fd_sc_hd__nand2_2
X_12594_ _12586_/B _12591_/B _12584_/X vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__a21o_1
X_11614_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11615_/B sky130_fd_sc_hd__or2_1
XFILLER_0_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09074__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11545_ _12310_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__A2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11476_ _11988_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11480_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13158__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13215_ _13215_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _13216_/B sky130_fd_sc_hd__nand2_1
X_10427_ hold257/A _10427_/A2 _10425_/X _12433_/A1 vssd1 vssd1 vccd1 vccd1 _10427_/X
+ sky130_fd_sc_hd__a31o_1
Xmax_cap219 _07146_/A vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__buf_4
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13146_ _13146_/A _13146_/B vssd1 vssd1 vccd1 vccd1 _13146_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10358_ _10189_/A _10189_/B _10186_/A vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ hold6/X _13108_/B2 rst vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__a21oi_1
X_10289_ hold232/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10554_/C sky130_fd_sc_hd__or2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12133__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _12420_/A _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06899__A1 _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07560__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__A1 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11644__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ reg1_val[9] reg1_val[22] _09180_/S vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ _09941_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08124_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10080__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _08052_/A _08052_/B _08052_/C vssd1 vssd1 vccd1 vccd1 _08063_/A sky130_fd_sc_hd__or3_1
XFILLER_0_114_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12357__C1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ _07021_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07003_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout105_A _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ _10234_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08956_/B sky130_fd_sc_hd__xnor2_1
X_07905_ _09938_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _07908_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07336__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ _07944_/B _07212_/X _07218_/Y fanout28/X vssd1 vssd1 vccd1 vccd1 _08886_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11883__A1 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _08556_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _07871_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09828__A1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _07737_/Y _07740_/X _07786_/B vssd1 vssd1 vccd1 vccd1 _07767_/X sky130_fd_sc_hd__a21o_1
X_06718_ _06799_/A _06631_/A _12696_/B _06717_/X vssd1 vssd1 vccd1 vccd1 _07251_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__11635__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_2_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07071__A _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07303__A2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ _07171_/X _09450_/B1 _07263_/Y _07182_/Y vssd1 vssd1 vccd1 vccd1 _07699_/B
+ sky130_fd_sc_hd__a22o_1
X_06649_ _06706_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _06649_/Y sky130_fd_sc_hd__nor2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _12053_/A1 _09258_/X _09259_/Y _09436_/X vssd1 vssd1 vccd1 vccd1 dest_val[1]
+ sky130_fd_sc_hd__a31o_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout18_A _08985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ _07593_/A _07593_/B _08633_/B vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _08556_/A _08319_/B vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10071__B1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11228_/A _11226_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _12202_/A fanout46/X fanout44/X _12059_/A vssd1 vssd1 vccd1 vccd1 _11262_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08016__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ _11192_/A _11192_/B vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__and2_1
X_13000_ _13144_/A hold205/X vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__and2_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11626__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10976_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__and3_1
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12715_ reg1_val[20] _12767_/B vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ reg1_val[6] _12647_/B vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _12578_/B vssd1 vssd1 vccd1 vccd1 _12577_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11231__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
X_11528_ hold216/A hold326/A _11528_/C vssd1 vssd1 vccd1 vccd1 _11620_/B sky130_fd_sc_hd__or3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11459_ _11458_/A _11458_/B _11460_/A vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__o21a_1
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13129_ _13134_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13348_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ _08670_/A _08670_/B _08670_/C vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__and3_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07621_ _09766_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07623_/B sky130_fd_sc_hd__xor2_1
X_07552_ _07732_/A _07732_/B _07549_/Y vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__09286__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07483_ _07359_/A _07359_/B _07361_/B _07362_/B _07362_/A vssd1 vssd1 vccd1 vccd1
+ _07486_/A sky130_fd_sc_hd__o32a_2
XANTENNA__08494__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ _12415_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09222_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ _12415_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09153_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08104_ _08104_/A _08104_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09084_ _09659_/B2 fanout77/X fanout73/X _11386_/A vssd1 vssd1 vccd1 vccd1 _09085_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ _08035_/A _08035_/B vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09746__B1 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09986_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__xor2_1
X_08937_ _08937_/A _08937_/B vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__xnor2_1
X_08868_ reg1_val[28] reg1_val[29] _08868_/C _12756_/B vssd1 vssd1 vccd1 vccd1 _08983_/B
+ sky130_fd_sc_hd__or4_2
X_07819_ _08633_/B fanout98/X fanout83/X _09300_/A vssd1 vssd1 vccd1 vccd1 _07820_/B
+ sky130_fd_sc_hd__o22a_1
X_08799_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _12229_/B sky130_fd_sc_hd__xnor2_2
X_10830_ _11052_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10832_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10761_ _10761_/A _10761_/B vssd1 vssd1 vccd1 vccd1 _10764_/C sky130_fd_sc_hd__xor2_1
XANTENNA__12281__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ _10599_/A _10599_/B _10595_/X vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__a21oi_1
X_12500_ _12509_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12502_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ _12417_/A _12431_/A2 _09252_/X _09223_/Y _12430_/X vssd1 vssd1 vccd1 vccd1
+ _12431_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12362_ _08857_/Y _11917_/C _12360_/X _12410_/S vssd1 vssd1 vccd1 vccd1 _12364_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11316_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11986__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ hold242/A _12293_/B vssd1 vssd1 vccd1 vccd1 _12345_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11244_ _11879_/A2 _11341_/B hold331/A vssd1 vssd1 vccd1 vccd1 _11244_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11544__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06799__B _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08360__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ _12065_/A _11175_/B vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__xor2_1
X_10126_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__and2_1
XANTENNA__08960__A1 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08960__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _10058_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap118_A _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10959_ _10959_/A _10959_/B _10959_/C vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__and3_1
XFILLER_0_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08228__B1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ _12629_/A _12629_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold327/X vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__clkbuf_2
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07203__A1 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _09840_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07203__B2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _07402_/B _07212_/X _07218_/Y fanout41/X vssd1 vssd1 vccd1 vccd1 _09772_/B
+ sky130_fd_sc_hd__a22o_1
X_06983_ reg1_val[4] _07063_/C _07093_/A vssd1 vssd1 vccd1 vccd1 _06984_/B sky130_fd_sc_hd__o21a_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08670_/B _08670_/C _08670_/A vssd1 vssd1 vccd1 vccd1 _08723_/B sky130_fd_sc_hd__a21oi_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12520__A _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__B1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _08653_/A _08659_/S vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__xor2_1
X_07604_ _10231_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07605_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07535_ _07541_/B _07541_/C _07541_/A vssd1 vssd1 vccd1 vccd1 _07543_/A sky130_fd_sc_hd__o21a_1
X_07466_ _08650_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _09203_/X _09204_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A1 _11853_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ _07418_/A _07418_/B vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__nor2_1
X_09136_ _09023_/A _09023_/B _09021_/Y vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09067_ _09067_/A _09067_/B vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06796__A3 _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ _08551_/A2 _08400_/B fanout82/X _08551_/B1 vssd1 vssd1 vccd1 vccd1 _08019_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08180__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout85_A _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _11557_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__xnor2_2
X_12980_ _13144_/A hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__and2_1
XANTENNA__09215__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11931_ _12011_/B _11931_/B vssd1 vssd1 vccd1 vccd1 _11933_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11862_ _11862_/A _12020_/C vssd1 vssd1 vccd1 vccd1 _11862_/Y sky130_fd_sc_hd__nor2_1
X_10813_ _10755_/A _10755_/B _10756_/Y vssd1 vssd1 vccd1 vccd1 _10882_/A sky130_fd_sc_hd__o21ai_2
X_11793_ _11793_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _10745_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08355__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10675_ _09886_/B _12394_/A1 _10675_/S vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _12403_/X _12411_/Y _12412_/X _12413_/Y _09149_/X vssd1 vssd1 vccd1 vccd1
+ _12414_/X sky130_fd_sc_hd__a311o_2
XANTENNA__10568__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ hold251/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12276_ _12369_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12280_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11517__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11227_ _06830_/Y _11226_/X _11781_/S vssd1 vssd1 vccd1 vccd1 _11228_/B sky130_fd_sc_hd__mux2_1
X_11158_ _11159_/B _11158_/B vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12190__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__xnor2_4
X_11089_ _11087_/Y _11089_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12796__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ _07321_/A _07321_/B vssd1 vssd1 vccd1 vccd1 _07320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _07251_/A _07251_/B vssd1 vssd1 vccd1 vccd1 _07251_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07182_ _11361_/A _07172_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07182_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09823_ _09823_/A _09823_/B vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06935__B1 _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__B2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ _07016_/A _06994_/A _06966_/C vssd1 vssd1 vccd1 vccd1 _07028_/B sky130_fd_sc_hd__nand3_2
XANTENNA__09543__B _09543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ curr_PC[0] curr_PC[1] curr_PC[2] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06897_ instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1 vccd1 _06897_/Y
+ sky130_fd_sc_hd__a21oi_2
XANTENNA__09885__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09685_/Y sky130_fd_sc_hd__nor2_1
X_08705_ _08705_/A _08705_/B vssd1 vssd1 vccd1 vccd1 _08792_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10495__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08638_/A _08638_/C _08638_/B vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout22 _07347_/B vssd1 vssd1 vccd1 vccd1 fanout22/X sky130_fd_sc_hd__buf_6
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout11 _08858_/Y vssd1 vssd1 vccd1 vccd1 fanout11/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08567_ _07010_/Y _07114_/X _07146_/Y _07018_/X vssd1 vssd1 vccd1 vccd1 _08568_/B
+ sky130_fd_sc_hd__a22o_1
Xfanout55 _07030_/Y vssd1 vssd1 vccd1 vccd1 fanout55/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout44 fanout45/X vssd1 vssd1 vccd1 vccd1 fanout44/X sky130_fd_sc_hd__clkbuf_8
Xfanout33 _07181_/X vssd1 vssd1 vccd1 vccd1 fanout33/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07112__B1 _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ _07518_/A _07518_/B _07518_/C vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__nand3_1
X_08498_ _08499_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout66 fanout67/X vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__clkbuf_8
Xfanout77 _08274_/B vssd1 vssd1 vccd1 vccd1 fanout77/X sky130_fd_sc_hd__buf_6
Xfanout88 _11054_/A vssd1 vssd1 vccd1 vccd1 _11557_/A sky130_fd_sc_hd__clkbuf_16
Xfanout99 _07076_/Y vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__buf_6
XFILLER_0_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07449_ _07451_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07548_/B sky130_fd_sc_hd__or2_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _10461_/B _10461_/A vssd1 vssd1 vccd1 vccd1 _10635_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _11359_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09120_/B sky130_fd_sc_hd__xnor2_1
X_10391_ _10243_/A _10243_/C _10243_/B vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12130_ fanout14/X _12309_/A fanout12/X fanout22/X vssd1 vssd1 vccd1 vccd1 _12131_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _11980_/A _12404_/B _12056_/B _11984_/A vssd1 vssd1 vccd1 vccd1 _12075_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _06879_/D _10898_/B _10918_/S vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10722__B2 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07254__A _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ hold222/X _13095_/B2 _13158_/A2 hold232/X vssd1 vssd1 vccd1 vccd1 hold233/A
+ sky130_fd_sc_hd__a22o_1
X_11914_ _11988_/A _11914_/B vssd1 vssd1 vccd1 vccd1 _11921_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ _13092_/A _13093_/A _13092_/B vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__a21bo_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11776_ _11776_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__or2_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10727_ _10727_/A _10727_/B vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09909__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11738__B1 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ _06747_/Y _10542_/X _06749_/B vssd1 vssd1 vccd1 vccd1 _10658_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589_ _10589_/A _11296_/B _10590_/A vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__or3_1
XANTENNA__12335__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ instruction[12] vssd1 vssd1 vccd1 vccd1 loadstore_dest[1] sky130_fd_sc_hd__buf_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12328_ _11773_/B _12088_/B _12324_/X _12327_/X vssd1 vssd1 vccd1 vccd1 _12329_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10410__B1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10961__B2 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__A1 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ fanout14/X fanout6/X _11813_/A vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07709__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__A3 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06878_/A _06818_/X _06819_/X vssd1 vssd1 vccd1 vccd1 _06820_/Y sky130_fd_sc_hd__a21oi_1
X_06751_ _06799_/A _06631_/A _12662_/B _06750_/X vssd1 vssd1 vccd1 vccd1 _07195_/A
+ sky130_fd_sc_hd__a31o_4
X_06682_ _11797_/S _06682_/B vssd1 vssd1 vccd1 vccd1 _11782_/A sky130_fd_sc_hd__nor2_2
X_09470_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09470_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ _08425_/A _08425_/B vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08352_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _08352_/X sky130_fd_sc_hd__and2_1
XFILLER_0_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11977__B1 _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ _08551_/B2 fanout55/X _12257_/A _06973_/A vssd1 vssd1 vccd1 vccd1 _07304_/B
+ sky130_fd_sc_hd__o22a_1
X_08283_ _08649_/B _08354_/A2 _10585_/B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08284_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _10230_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07236_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout135_A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07165_ reg1_val[11] reg1_val[12] reg1_val[13] _07229_/C _07229_/B vssd1 vssd1 vccd1
+ vccd1 _07246_/B sky130_fd_sc_hd__o41a_2
X_07096_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07096_/X sky130_fd_sc_hd__and2_2
XANTENNA__07948__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout201 _13158_/A2 vssd1 vssd1 vccd1 vccd1 _13209_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout223 _11238_/S vssd1 vssd1 vccd1 vccd1 _11958_/A sky130_fd_sc_hd__clkbuf_8
Xfanout212 _07129_/A vssd1 vssd1 vccd1 vccd1 _09722_/S sky130_fd_sc_hd__buf_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11901__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 _06893_/Y vssd1 vssd1 vccd1 vccd1 _12504_/S sky130_fd_sc_hd__clkbuf_8
Xfanout256 _06564_/A vssd1 vssd1 vccd1 vccd1 _13095_/B2 sky130_fd_sc_hd__buf_4
Xfanout234 _09229_/X vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__buf_4
Xfanout278 _12978_/A vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10180__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09938_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__xnor2_1
Xfanout289 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__clkbuf_16
Xfanout267 _06591_/X vssd1 vssd1 vccd1 vccd1 _12767_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__08373__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ _07998_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07074__A _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _12335_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _06949_/Y sky130_fd_sc_hd__nand2_2
X_09737_ _11235_/S _09736_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _09737_/X sky130_fd_sc_hd__o21a_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09670_/B sky130_fd_sc_hd__xnor2_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A _09599_/B _09598_/X vssd1 vssd1 vccd1 vccd1 _09599_/X sky130_fd_sc_hd__or3b_1
X_08619_ _12785_/A _08619_/A2 _08619_/B1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 _08620_/B
+ sky130_fd_sc_hd__o22a_1
X_11630_ _11630_/A _11630_/B _11630_/C _11630_/D vssd1 vssd1 vccd1 vccd1 _11630_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11561_ _11561_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09625__A2 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ _13372_/CLK hold190/X vssd1 vssd1 vccd1 vccd1 _13300_/Q sky130_fd_sc_hd__dfxtp_1
X_10512_ _10371_/B _10387_/B _10369_/Y vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11494_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11978__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08633__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ hold197/X _12780_/B hold328/X _06564_/A vssd1 vssd1 vccd1 vccd1 _13233_/B
+ sky130_fd_sc_hd__a22o_1
X_10443_ _10402_/A _10401_/B _10401_/A vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ hold320/A _13161_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12393__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _11172_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _12178_/A2 _12176_/B hold188/A vssd1 vssd1 vccd1 vccd1 _12113_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10943__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13093_/Y sky130_fd_sc_hd__xnor2_1
X_12044_ _09595_/B _12043_/X _06642_/B vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08364__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ _13215_/A _13216_/A _13215_/B vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09403__S _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ hold309/X hold29/X vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07875__B2 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07875__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11829_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__or2_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _11760_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12065__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12384__B1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ _09671_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09001__B1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ _07921_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10698__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07852_/A _07852_/B vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ _12621_/A _09725_/S vssd1 vssd1 vccd1 vccd1 _06803_/X sky130_fd_sc_hd__and2_1
X_09522_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08107__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07783_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06734_ reg2_val[11] _06794_/B vssd1 vssd1 vccd1 vccd1 _06734_/X sky130_fd_sc_hd__and2_1
X_06665_ reg2_val[22] _06712_/B _06707_/B1 _06664_/Y vssd1 vssd1 vccd1 vccd1 _06994_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA_fanout252_A _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _09452_/B _09453_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09384_ _09380_/X _09383_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__mux2_1
X_08404_ _06875_/A _10585_/B2 _10067_/A1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08405_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09068__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06596_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06596_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__09607__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ _08335_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08266_ _08776_/B _08687_/B vssd1 vssd1 vccd1 vccd1 _08266_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07217_ _07217_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _10490_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13278__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ _08220_/A _08220_/B _08186_/X vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__a21oi_2
X_07148_ _07148_/A _07148_/B _07148_/C vssd1 vssd1 vccd1 vccd1 _07150_/A sky130_fd_sc_hd__and3_1
XANTENNA__10925__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__A2 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12127__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _09659_/B2 _10233_/B2 fanout98/X _10233_/A1 vssd1 vssd1 vccd1 vccd1 _07080_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10090_ _10091_/B _10091_/A vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10223__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _10213_/A _13072_/A2 hold30/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold31/A
+ sky130_fd_sc_hd__o211a_1
X_10992_ _10992_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10993_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12737_/C _12730_/B _12728_/A vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__11054__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ reg1_val[9] _12662_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__nand2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12593_ _12610_/A _12593_/B vssd1 vssd1 vccd1 vccd1 _12598_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11544_ fanout57/X fanout22/X fanout14/X _11837_/A vssd1 vssd1 vccd1 vccd1 _11545_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ _11645_/A fanout9/X fanout4/X fanout51/X vssd1 vssd1 vccd1 vccd1 _11476_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13158__A2 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ _13226_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13366_/D sky130_fd_sc_hd__and2_1
X_10426_ _10427_/A2 _10425_/X hold257/A vssd1 vssd1 vccd1 vccd1 _10426_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13146_/B sky130_fd_sc_hd__nand2_1
X_10357_ _10357_/A _10357_/B vssd1 vssd1 vccd1 vccd1 _10370_/A sky130_fd_sc_hd__xnor2_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _08872_/B _12797_/B hold25/X vssd1 vssd1 vccd1 vccd1 _13336_/D sky130_fd_sc_hd__a21oi_1
X_10288_ _10285_/X _10287_/X _10288_/S vssd1 vssd1 vccd1 vccd1 _10288_/X sky130_fd_sc_hd__mux2_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ _06655_/B _12025_/X _12026_/Y vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11644__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ hold299/X hold77/X vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07442__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__A _09370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08120_ _08619_/A2 _08354_/A2 fanout71/X _08619_/B2 vssd1 vssd1 vccd1 vccd1 _08121_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08273__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10080__A1 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ _08048_/A _08048_/C _08048_/B vssd1 vssd1 vccd1 vccd1 _08052_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__08025__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ _09668_/A _07002_/B vssd1 vssd1 vccd1 vccd1 _07021_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ fanout56/X _10233_/B2 _10233_/A1 fanout62/X vssd1 vssd1 vccd1 vccd1 _08954_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ _08590_/B fanout75/X fanout71/X _09648_/A vssd1 vssd1 vccd1 vccd1 _07905_/B
+ sky130_fd_sc_hd__o22a_1
X_08884_ _09795_/A _08884_/B vssd1 vssd1 vccd1 vccd1 _08888_/A sky130_fd_sc_hd__xnor2_1
X_07835_ _08507_/A2 _08354_/A2 fanout71/X _08533_/B vssd1 vssd1 vccd1 vccd1 _07836_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13085__B2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _07851_/A _07851_/B _07754_/X vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__12832__A1 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06717_ reg2_val[14] _06767_/A vssd1 vssd1 vccd1 vccd1 _06717_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09828__A2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _09505_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10843__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09377_/Y _09427_/X _09435_/X _12504_/S vssd1 vssd1 vccd1 vccd1 _09436_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08500__A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _10468_/A _07697_/B vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__xnor2_4
X_06648_ instruction[36] _06657_/B vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__and2_4
XFILLER_0_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ instruction[14] _06575_/X _06578_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__o211a_4
X_09367_ _09367_/A _09367_/B vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__xor2_4
XANTENNA_50 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _09671_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08318_ _08533_/B _08553_/A2 _08553_/B1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08319_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10071__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08249_ _08249_/A _08249_/B vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_105_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08016__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _11183_/A _11183_/B _11180_/A vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08016__B2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11192_/B sky130_fd_sc_hd__nand2_1
X_10211_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08567__A2 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10142_ _06812_/X _10141_/Y _12025_/S vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07775__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07527__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10073_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07262__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _10975_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10976_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10834__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12716_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _12644_/A _12641_/Y _12643_/B vssd1 vssd1 vccd1 vccd1 _12649_/A sky130_fd_sc_hd__o21a_2
XANTENNA__13203__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ _12598_/A _12600_/A vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11527_ _11527_/A _11527_/B vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10062__B2 _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _11458_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__nor2_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11390_/C sky130_fd_sc_hd__xnor2_1
X_10409_ _11776_/A _08721_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__o21ai_1
X_13128_ hold308/X _13209_/A2 _13127_/X _13143_/B2 vssd1 vssd1 vccd1 vccd1 _13129_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ hold137/A _13071_/A2 _13071_/B1 hold111/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold112/A sky130_fd_sc_hd__o221a_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08191__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _07101_/Y _07539_/B fanout37/X _07114_/X vssd1 vssd1 vccd1 vccd1 _07621_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ _07551_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07732_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12814__A1 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07482_ _07399_/A _07399_/B _07411_/B _07414_/A vssd1 vssd1 vccd1 vccd1 _07487_/A
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__08494__A1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__B2 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ _11238_/S _09217_/Y _09220_/Y _09243_/B vssd1 vssd1 vccd1 vccd1 _09221_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _11781_/S _09222_/B vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09443__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ _08103_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _08104_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout215_A _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09827__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _08035_/A _08035_/B vssd1 vssd1 vccd1 vccd1 _08034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07757__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07509__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _08832_/A _08832_/B _08830_/Y vssd1 vssd1 vccd1 vccd1 _08937_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08880_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13058__A1 _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _08648_/A _07818_/B _07818_/C vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__nor3_1
X_08798_ _08797_/A _08797_/B _08792_/A _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1
+ _08798_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ _07910_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07808_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10816__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _10761_/B _10761_/A vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout30_A fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ _10637_/A _10637_/B _10638_/Y vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__a21bo_1
X_09419_ _09419_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09419_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _12772_/A _06644_/X _09235_/X _12429_/Y _11446_/B vssd1 vssd1 vccd1 vccd1
+ _12430_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _08857_/Y _12360_/X _12359_/Y vssd1 vssd1 vccd1 vccd1 _12410_/S sky130_fd_sc_hd__o21ai_1
X_11312_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__nand2_1
X_12292_ _11238_/S _12290_/X _12291_/X _06924_/Y vssd1 vssd1 vccd1 vccd1 _12304_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11243_ hold311/A hold319/A _11243_/C vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__or3_1
XANTENNA__11544__B2 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07257__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _11917_/B _07151_/A _07155_/A _06993_/Y vssd1 vssd1 vccd1 vccd1 _11175_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__or2_1
XANTENNA__08960__A2 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _09970_/A _09970_/B _09966_/X vssd1 vssd1 vccd1 vccd1 _10058_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10959_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11242__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _10647_/Y _11112_/A _10887_/Y vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08228__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ _12626_/Y _12628_/B vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08228__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ _12559_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11535__A1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _09773_/A vssd1 vssd1 vccd1 vccd1 _09770_/Y sky130_fd_sc_hd__inv_2
X_06982_ _07093_/A _07063_/C vssd1 vssd1 vccd1 vccd1 _06988_/B sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08721_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__and2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08652_ _08651_/B _08653_/A vssd1 vssd1 vccd1 vccd1 _08652_/X sky130_fd_sc_hd__and2b_1
X_07603_ fanout56/X _08590_/B _09648_/A fanout62/X vssd1 vssd1 vccd1 vccd1 _07604_/B
+ sky130_fd_sc_hd__o22a_1
X_08583_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__or2_1
XANTENNA__09664__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _07692_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _07541_/C sky130_fd_sc_hd__and2_1
XFILLER_0_119_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ fanout62/X _09297_/B2 _09297_/A1 fanout60/X vssd1 vssd1 vccd1 vccd1 _07466_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07630__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ reg1_val[12] reg1_val[19] _09560_/A vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07396_ _10937_/A _07396_/B vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12971__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09066_ _09067_/A _09067_/B vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08017_ _08320_/A _08017_/B vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07077__A _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ fanout51/X fanout27/X fanout25/X _11456_/A vssd1 vssd1 vccd1 vccd1 _09969_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ _08796_/B _08796_/C _09035_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08919_/X
+ sky130_fd_sc_hd__a211o_1
X_11930_ _11930_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__or2_1
X_09899_ _09155_/S _09875_/Y _09881_/X _09882_/X _09898_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10231__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _11862_/A _12020_/C vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ hold299/A _12175_/A2 _11877_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11793_/B
+ sky130_fd_sc_hd__a31o_1
X_10812_ _11776_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__or2_1
X_10743_ _10743_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10745_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11062__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__A1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ hold240/A _11115_/A _10791_/B _12433_/A1 vssd1 vssd1 vccd1 vccd1 _10674_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12413_ _12373_/Y _12374_/X _12411_/Y _12412_/X _06943_/Y vssd1 vssd1 vccd1 vccd1
+ _12413_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _11238_/S _09560_/B _12343_/X _09243_/B vssd1 vssd1 vccd1 vccd1 _12344_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09422__A3 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__A _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07969__B1 _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12275_ _11689_/B _12271_/X _12272_/Y _12274_/X vssd1 vssd1 vccd1 vccd1 _12276_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__A _10406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__A1 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__A1 _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ _06879_/B _11120_/B _11137_/S vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__a21o_1
X_11157_ _12193_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12621__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10108_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09406__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__nand2_1
X_10039_ _09992_/A _09992_/B _09990_/X vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__09930__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12068__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07250_ _07251_/A _07251_/B vssd1 vssd1 vccd1 vccd1 _07250_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12402__C1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07181_ _11361_/A _07172_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12953__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12181__A1 _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _09823_/A _09823_/B vssd1 vssd1 vccd1 vccd1 _09822_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10731__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _09232_/Y _09713_/Y _09714_/X _09752_/X _09712_/X vssd1 vssd1 vccd1 vccd1
+ _09753_/X sky130_fd_sc_hd__a311o_2
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _07016_/A _06994_/A _06966_/C vssd1 vssd1 vccd1 vccd1 _06967_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout282_A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _09035_/A _09371_/A vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__xnor2_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06896_ reg1_idx[2] _06908_/C _06896_/C vssd1 vssd1 vccd1 vccd1 int_return sky130_fd_sc_hd__and3_4
XANTENNA__10051__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__A2_N _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _09684_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10495__A1 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__B2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08635_ _08629_/A _08629_/C _08629_/B vssd1 vssd1 vccd1 vccd1 _08638_/C sky130_fd_sc_hd__o21ai_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08566_ _08566_/A _08566_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout12 _08858_/Y vssd1 vssd1 vccd1 vccd1 fanout12/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07517_ _07475_/A _07475_/B _07474_/X vssd1 vssd1 vccd1 vccd1 _07518_/C sky130_fd_sc_hd__o21bai_1
Xfanout56 _07015_/X vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__buf_8
Xfanout23 _07346_/Y vssd1 vssd1 vccd1 vccd1 _07347_/B sky130_fd_sc_hd__clkbuf_8
Xfanout45 _07117_/X vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__buf_6
XANTENNA__07112__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout34 _07172_/Y vssd1 vssd1 vccd1 vccd1 _08184_/B sky130_fd_sc_hd__buf_6
X_08497_ _09941_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout78 _07249_/Y vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__buf_8
Xfanout67 _06971_/Y vssd1 vssd1 vccd1 vccd1 fanout67/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 _09766_/A vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__buf_8
X_07448_ _07448_/A _07448_/B _07516_/A vssd1 vssd1 vccd1 vccd1 _07449_/B sky130_fd_sc_hd__nor3_1
X_07379_ _07379_/A _07379_/B vssd1 vssd1 vccd1 vccd1 _07380_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09287__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _10222_/A2 _07944_/B fanout28/X _10712_/A vssd1 vssd1 vccd1 vccd1 _09119_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09049_ _07539_/B _10326_/A _09450_/B1 fanout37/X vssd1 vssd1 vccd1 vccd1 _09050_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ _12060_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12077_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12172__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _11776_/A _11011_/B _11011_/C vssd1 vssd1 vccd1 vccd1 _11011_/X sky130_fd_sc_hd__or3_1
XANTENNA__10722__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ _12978_/A hold223/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__and2_1
X_11913_ _12059_/A fanout9/X fanout4/X _11980_/A vssd1 vssd1 vccd1 vccd1 _11914_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12893_ hold48/X hold322/A vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__nand2b_1
X_11844_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__or2_1
XFILLER_0_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07270__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11774_/A _11808_/D _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11435__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10726_/A _10726_/B vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _10657_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _10657_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10588_ _10589_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ instruction[11] vssd1 vssd1 vccd1 vccd1 loadstore_dest[0] sky130_fd_sc_hd__buf_12
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ _12217_/Y _12406_/A _12325_/Y _12326_/X vssd1 vssd1 vccd1 vccd1 _12327_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10961__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12262_/A sky130_fd_sc_hd__xnor2_1
X_11209_ _11209_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08367__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ curr_PC[27] _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__xor2_1
XANTENNA__07445__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__A4 _07089_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ reg2_val[8] _06794_/B vssd1 vssd1 vccd1 vccd1 _06750_/X sky130_fd_sc_hd__and2_1
X_06681_ reg1_val[21] _06681_/B vssd1 vssd1 vccd1 vccd1 _06682_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09660__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ _08420_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08425_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07180__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11977__A1 _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07302_ _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _07302_/X sky130_fd_sc_hd__or2_2
XFILLER_0_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ reg1_val[12] _07233_/B vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12526__A _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ reg1_val[17] _07164_/B vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07095_ reg1_val[23] _07190_/B _07095_/C vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__or3_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout202 _06901_/Y vssd1 vssd1 vccd1 vccd1 _13158_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout213 _06796_/X vssd1 vssd1 vccd1 vccd1 _07129_/A sky130_fd_sc_hd__buf_4
Xfanout246 _06893_/Y vssd1 vssd1 vccd1 vccd1 _12615_/S sky130_fd_sc_hd__clkbuf_8
Xfanout224 _06767_/X vssd1 vssd1 vccd1 vccd1 _11238_/S sky130_fd_sc_hd__buf_4
Xfanout235 _09229_/X vssd1 vssd1 vccd1 vccd1 _12431_/A2 sky130_fd_sc_hd__buf_2
Xfanout279 _13219_/A vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__buf_4
Xfanout268 _06767_/A vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__buf_4
Xfanout257 _06564_/A vssd1 vssd1 vccd1 vccd1 _13108_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09805_ _09648_/A fanout13/X fanout11/X _08590_/B vssd1 vssd1 vccd1 vccd1 _09806_/B
+ sky130_fd_sc_hd__o22a_1
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__xnor2_4
X_09736_ _10148_/S _09198_/X _09249_/B vssd1 vssd1 vccd1 vccd1 _09736_/X sky130_fd_sc_hd__o21a_1
X_06948_ _12335_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07195_/B sky130_fd_sc_hd__and2_2
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _09300_/A fanout11/X fanout7/X _08633_/B vssd1 vssd1 vccd1 vccd1 _09668_/B
+ sky130_fd_sc_hd__o22a_1
X_06879_ _11228_/A _06879_/B _11014_/A _06879_/D vssd1 vssd1 vccd1 vccd1 _06880_/D
+ sky130_fd_sc_hd__or4_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08610_/A _08610_/B _08610_/C vssd1 vssd1 vccd1 vccd1 _08622_/B sky130_fd_sc_hd__a21oi_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09583_/Y _09584_/X _09589_/Y _09597_/X vssd1 vssd1 vccd1 vccd1 _09598_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08549_ _08549_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__xor2_2
X_11560_ _11561_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__or2_1
XFILLER_0_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11968__A1 _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08833__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08833__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11399_/A _11398_/B _11396_/X vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__a21oi_2
X_13230_ hold193/X hold149/X _13236_/A _13229_/X vssd1 vssd1 vccd1 vccd1 hold194/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08633__B _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ _10315_/B _10406_/X _10315_/A vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13161_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _13161_/Y sky130_fd_sc_hd__xnor2_1
X_10373_ fanout58/X fanout35/X fanout33/X fanout56/X vssd1 vssd1 vccd1 vccd1 _10374_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10943__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ hold228/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__or2_1
X_13092_ _13092_/A _13092_/B vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12043_ _11966_/B _09228_/Y _12043_/S vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12171__A _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__B _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ hold129/X hold307/A vssd1 vssd1 vccd1 vccd1 _13215_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08521__B1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ hold313/A hold15/X vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08096__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07875__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11906_/B _11827_/B vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__and2_1
XFILLER_0_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11758_ _11758_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11760_/B sky130_fd_sc_hd__xnor2_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__A1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ _11296_/B _10709_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11689_ _11854_/A _11689_/B vssd1 vssd1 vccd1 vccd1 _11808_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ _13363_/CLK _13359_/D vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09655__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07920_ _07920_/A _07920_/B vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09001__B2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A1 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__B2 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _07851_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _07852_/B sky130_fd_sc_hd__xor2_2
X_06802_ _06875_/A _09396_/S vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nand2_1
X_07782_ _09630_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06733_ _06879_/D vssd1 vssd1 vccd1 vccd1 _06733_/Y sky130_fd_sc_hd__inv_2
X_09521_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__and2b_1
X_06664_ _06706_/A _12652_/B vssd1 vssd1 vccd1 vccd1 _06664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09453_/B _09452_/B vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__and2b_1
X_06595_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06595_/X sky130_fd_sc_hd__o211a_1
X_09383_ _09381_/X _09382_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09383_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09068__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ _08416_/A _08416_/B vssd1 vssd1 vccd1 vccd1 _08403_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout245_A _06893_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _08341_/B _08341_/A vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07079__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08265_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08687_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07216_ _07195_/A _07113_/A _06954_/B _07299_/B vssd1 vssd1 vccd1 vccd1 _07218_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12375__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ reg1_val[24] _07147_/B vssd1 vssd1 vccd1 vccd1 _07148_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _07072_/B _10339_/A _10234_/A vssd1 vssd1 vccd1 vccd1 _07078_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10689__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout60_A _06999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ _10992_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ _09389_/X _09399_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09719_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13372_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12737_/C _12730_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xor2_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ reg1_val[9] _12662_/B vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__or2_1
X_11612_ _11612_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__or3_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12592_ reg1_val[23] curr_PC[23] _12615_/S vssd1 vssd1 vccd1 vccd1 _12593_/B sky130_fd_sc_hd__mux2_2
X_11543_ _11492_/A _11492_/B _11493_/Y vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ _12310_/A _11474_/B vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13213_ hold307/X _13222_/A2 _13212_/X _12781_/A vssd1 vssd1 vccd1 vccd1 _13214_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ hold247/A _10554_/C vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__or2_1
XANTENNA__09231__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13144_ _13144_/A _13144_/B vssd1 vssd1 vccd1 vccd1 _13351_/D sky130_fd_sc_hd__and2_1
XANTENNA__09475__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10357_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12118__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12118__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ hold24/X _13108_/B2 _13222_/A2 hold6/X rst vssd1 vssd1 vccd1 vccd1 hold25/A
+ sky130_fd_sc_hd__a221o_1
X_10287_ _09251_/A _10286_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__mux2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _06655_/B _12025_/X _09227_/X vssd1 vssd1 vccd1 vccd1 _12026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ _13179_/A _13180_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12859_ hold108/X hold289/X vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12054__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08554__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09369__B _09370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10080__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _08050_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08052_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ _08633_/B fanout62/X _09300_/A fanout60/X vssd1 vssd1 vccd1 vccd1 _07002_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06802__A _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _08952_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08955_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11868__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ _07899_/Y _07901_/X _07902_/A vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__a21oi_1
X_08883_ _10859_/A _08096_/B fanout24/X _10327_/B2 vssd1 vssd1 vccd1 vccd1 _08884_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07834_ _07834_/A _07834_/B vssd1 vssd1 vccd1 vccd1 _07837_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13085__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _07765_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07851_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__11155__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06716_ _11246_/S _06716_/B vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__nor2_1
X_09504_ _09505_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09504_/Y sky130_fd_sc_hd__nor2_1
X_07696_ _10585_/B2 _08400_/B fanout82/X _10067_/A1 vssd1 vssd1 vccd1 vccd1 _07697_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__10843__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12832__A2 _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ reg1_val[31] _07127_/B vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__xnor2_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _09560_/A _09434_/Y _09430_/Y _12029_/A vssd1 vssd1 vccd1 vccd1 _09435_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10843__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06578_ instruction[21] _06922_/B vssd1 vssd1 vccd1 vccd1 _06578_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12045__B1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09367_/A _09367_/B vssd1 vssd1 vccd1 vccd1 _09366_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_40 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _09297_/A1 fanout11/X fanout7/X _09297_/B2 vssd1 vssd1 vccd1 vccd1 _09298_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08317_ _08573_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10071__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08248_ _08248_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08249_/B sky130_fd_sc_hd__and2_1
XFILLER_0_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _11645_/B _10210_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__xnor2_1
X_08179_ _08594_/A2 _10067_/A1 _08926_/B1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08180_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08016__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__or2_1
XFILLER_0_113_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07775__A1 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__B1 _06644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _06774_/A _10006_/B _06772_/Y vssd1 vssd1 vccd1 vccd1 _10141_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07775__B2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _12193_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__C1 _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ _10975_/B _10975_/A vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10834__A1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ reg1_val[19] _12767_/B vssd1 vssd1 vccd1 vccd1 _12716_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__10834__B2 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08374__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ _12644_/A _12644_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _12575_/A _12575_/B _12575_/C vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__and3_1
XFILLER_0_93_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ hold295/A _11879_/A2 _11623_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11527_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10062__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11457_ _11457_/A _11576_/A vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11388_/Y sky130_fd_sc_hd__nand2b_1
X_10408_ _10315_/X _10406_/X _10407_/Y vssd1 vssd1 vccd1 vccd1 _10408_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13127_ hold303/X _13126_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__mux2_1
X_10339_ _10339_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10339_/Y sky130_fd_sc_hd__nor2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _11559_/A _13078_/B2 hold138/X vssd1 vssd1 vccd1 vccd1 _13327_/D sky130_fd_sc_hd__o21a_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _12011_/A _12011_/B _12011_/C vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08191__A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ _07550_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09220_ _09411_/A _09219_/X _11958_/A vssd1 vssd1 vccd1 vccd1 _09220_/Y sky130_fd_sc_hd__a21oi_2
X_07481_ _07546_/A _07546_/B _07452_/X vssd1 vssd1 vccd1 vccd1 _07488_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08494__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11703__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08284__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _09233_/A _09229_/B _06872_/Y vssd1 vssd1 vccd1 vccd1 _09151_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__A1 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__B2 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__and2b_1
X_08102_ _08103_/B _08103_/A vssd1 vssd1 vccd1 vccd1 _08102_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08033_ _10081_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08035_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12534__A _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout110_A _07213_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__A1 _10766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07757__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__B _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _09984_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07509__B2 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A1 _07048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ _08935_/A _08935_/B vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13058__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _07818_/B _07818_/C _08648_/A vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__o21a_1
X_08797_ _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__nand2_1
X_07748_ _08533_/B fanout75/X fanout71/X _08507_/A2 vssd1 vssd1 vccd1 vccd1 _07749_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10816__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__B2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _08566_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07685_/A sky130_fd_sc_hd__xnor2_2
X_09418_ _12415_/A _12785_/A _09418_/C vssd1 vssd1 vccd1 vccd1 _09418_/X sky130_fd_sc_hd__or3_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ _11809_/A _10810_/A _11863_/A vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _09349_/A _09349_/B vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__xor2_2
X_12360_ fanout6/X _12360_/B vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _11311_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__xnor2_2
X_12291_ _12421_/B _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _11242_/A _11242_/B _11242_/C vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__or3_1
XANTENNA__07538__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11544__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _11173_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07748__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10957_ _11359_/A _10957_/B vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12619__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10888_ _10888_/A _11001_/A vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06617__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ reg1_val[2] _12627_/B vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09425__B2 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08228__A2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _12575_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__A _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _12178_/A2 _11542_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11509_/Y sky130_fd_sc_hd__a21oi_1
X_12489_ _12495_/B _12489_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12801__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ _12619_/A _12621_/A reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07063_/C
+ sky130_fd_sc_hd__or4_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08720_ _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _08721_/B sky130_fd_sc_hd__xnor2_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08653_/A _08651_/B vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__and2b_1
X_07602_ _10230_/A _07602_/B vssd1 vssd1 vccd1 vccd1 _07605_/A sky130_fd_sc_hd__xnor2_1
X_08582_ _08561_/A _08561_/B _08561_/C vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09664__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ _09795_/A _07533_/B vssd1 vssd1 vccd1 vccd1 _07692_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09664__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ _07477_/B _07520_/A _07477_/A vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ reg1_val[13] reg1_val[18] _09560_/A vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07395_ _07492_/A _07492_/B vssd1 vssd1 vccd1 vccd1 _07418_/A sky130_fd_sc_hd__or2_1
X_09134_ _09134_/A _09134_/B vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_71_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09065_ _09277_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__and2_1
XFILLER_0_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08016_ _08553_/A2 _08274_/B fanout74/X _08553_/B1 vssd1 vssd1 vccd1 vccd1 _08017_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__xor2_2
X_08918_ _09035_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08918_/X sky130_fd_sc_hd__or2_1
XANTENNA__07093__A _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ _09898_/A _09898_/B _09885_/X vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__or3b_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08849_ fanout83/X fanout77/X fanout73/X fanout79/X vssd1 vssd1 vccd1 vccd1 _08850_/B
+ sky130_fd_sc_hd__o22a_1
X_11860_ _12014_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _12020_/C sky130_fd_sc_hd__xnor2_2
X_11791_ _11879_/A2 _11877_/B hold299/A vssd1 vssd1 vccd1 vccd1 _11793_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12439__A _12619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _11809_/A _11041_/A vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__and2b_1
X_10742_ _10742_/A _10742_/B vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__A2 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _11115_/A _10791_/B hold240/A vssd1 vssd1 vccd1 vccd1 _10673_/Y sky130_fd_sc_hd__a21oi_1
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12343_ _12421_/C _12342_/Y _12421_/B vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10422__C1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09467__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ _12153_/Y _12273_/Y _12271_/C vssd1 vssd1 vccd1 vccd1 _12274_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11225_ _11863_/A _08741_/X _08743_/X _11946_/A _11224_/Y vssd1 vssd1 vccd1 vccd1
+ _11253_/B sky130_fd_sc_hd__a311oi_4
X_11156_ _11749_/A _07402_/B fanout41/X _11734_/A vssd1 vssd1 vccd1 vccd1 _11157_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12190__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11087_/Y sky130_fd_sc_hd__nor2_1
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__xor2_4
XANTENNA__12621__B _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _10038_/A _10313_/A vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__or2_1
XFILLER_0_105_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ fanout40/X _07593_/Y _08857_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _11990_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09658__A _10613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _10081_/A _11168_/A _07180_/C vssd1 vssd1 vccd1 vccd1 _07180_/X sky130_fd_sc_hd__or3_4
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07178__A _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10716__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12181__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09823_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _09222_/Y _09728_/X _12291_/B _09155_/S _09751_/X vssd1 vssd1 vccd1 vccd1
+ _09752_/X sky130_fd_sc_hd__a221o_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _06996_/A _06964_/B vssd1 vssd1 vccd1 vccd1 _06966_/C sky130_fd_sc_hd__and2_2
XANTENNA__07117__S _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _08799_/A _08799_/B _08805_/A _07802_/X _07731_/Y vssd1 vssd1 vccd1 vccd1
+ _09371_/A sky130_fd_sc_hd__a32o_2
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06895_ reg1_idx[3] reg1_idx[0] reg1_idx[1] reg1_idx[4] vssd1 vssd1 vccd1 vccd1 _06896_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA_fanout275_A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10495__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _09301_/A _08644_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__mux2_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08605_/A _07101_/Y _07263_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _08566_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout13 _12309_/A vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__clkbuf_8
X_07516_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07518_/B sky130_fd_sc_hd__nor2_1
Xfanout46 _07814_/B vssd1 vssd1 vccd1 vccd1 fanout46/X sky130_fd_sc_hd__clkbuf_8
Xfanout35 _07172_/Y vssd1 vssd1 vccd1 vccd1 fanout35/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11444__B2 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _08619_/B2 _08553_/A2 _08553_/B1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08497_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout24 _07215_/Y vssd1 vssd1 vccd1 vccd1 fanout24/X sky130_fd_sc_hd__buf_6
Xfanout57 _07015_/X vssd1 vssd1 vccd1 vccd1 fanout57/X sky130_fd_sc_hd__buf_4
XFILLER_0_92_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout68 _09930_/A vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__clkbuf_16
Xfanout79 _11188_/A vssd1 vssd1 vccd1 vccd1 fanout79/X sky130_fd_sc_hd__buf_6
X_07447_ _07525_/A _07525_/B _07443_/X vssd1 vssd1 vccd1 vccd1 _07548_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07378_ _07379_/A _07379_/B vssd1 vssd1 vccd1 vccd1 _07385_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08073__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ _09117_/A _09117_/B vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09048_ _09051_/A vssd1 vssd1 vccd1 vccd1 _09048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout90_A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _11776_/A _11011_/B _11011_/C vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09325__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__A1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__B2 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ hold261/A _13095_/B2 _13158_/A2 hold222/X vssd1 vssd1 vccd1 vccd1 hold223/A
+ sky130_fd_sc_hd__a22o_1
X_11912_ _11820_/A _11820_/B _11830_/A vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12892_ _13087_/A _13088_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__a21bo_1
X_11843_ _11843_/A _11843_/B vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__xnor2_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11774_/A _11808_/D vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10726_/A _10726_/B vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _11863_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13375_ _13375_/CLK hold185/X vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__dfxtp_1
X_10587_ _10587_/A _10587_/B vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12326_ _12213_/A _12269_/A _12268_/A vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _12257_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__nor2_1
X_11208_ _11209_/A _11209_/B vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12188_ _12189_/B _12187_/Y _11975_/A _12185_/Y vssd1 vssd1 vccd1 vccd1 dest_val[26]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__08367__A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08367__B2 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__B2 _10171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ hold319/A _11243_/C vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__or2_1
XANTENNA__09316__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06680_ reg1_val[21] _06681_/B vssd1 vssd1 vccd1 vccd1 _11797_/S sky130_fd_sc_hd__and2_1
XFILLER_0_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07180__B _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__xnor2_2
X_07301_ _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _07301_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08281_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08281_/X sky130_fd_sc_hd__or2_1
X_07232_ reg1_val[11] _07229_/C _07229_/B vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07163_ reg1_val[17] _07164_/B vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _07190_/B _07095_/C reg1_val[23] vssd1 vssd1 vccd1 vccd1 _07148_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout203 _06901_/Y vssd1 vssd1 vccd1 vccd1 _13222_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout214 _07152_/A vssd1 vssd1 vccd1 vccd1 _10284_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11901__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout247 _06893_/Y vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__buf_6
Xfanout225 _06600_/Y vssd1 vssd1 vccd1 vccd1 _06707_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07030__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _09227_/X vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__clkbuf_8
X_09804_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__xor2_1
Xfanout269 _06767_/A vssd1 vssd1 vccd1 vccd1 _06712_/B sky130_fd_sc_hd__clkbuf_8
Xfanout258 _13204_/B2 vssd1 vssd1 vccd1 vccd1 _13143_/B2 sky130_fd_sc_hd__buf_4
X_07996_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07996_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13103__B2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _12171_/A _09728_/X _09733_/Y _09734_/X _12107_/B1 vssd1 vssd1 vccd1 vccd1
+ _09735_/X sky130_fd_sc_hd__o221a_1
X_06947_ _12621_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _07009_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _09666_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__xnor2_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06878_ _06878_/A _10280_/A vssd1 vssd1 vccd1 vccd1 _06880_/C sky130_fd_sc_hd__nand2_1
X_08617_ _08622_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08467__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _06793_/Y _09886_/B _09594_/X _09595_/Y _09596_/X vssd1 vssd1 vccd1 vccd1
+ _09597_/X sky130_fd_sc_hd__o2111a_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08548_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11968__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ _08445_/A _08517_/A _08518_/A vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__a21oi_1
X_11490_ _11490_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ _10509_/B _10509_/C _10509_/A vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09298__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06715__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ curr_PC[9] _10686_/C vssd1 vssd1 vccd1 vccd1 _10441_/X sky130_fd_sc_hd__xor2_1
X_13160_ _13160_/A _13160_/B vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10372_ _10372_/A _10372_/B vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09794__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ hold269/A _12175_/A2 _12173_/B _12110_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _12119_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_103_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13091_ _13109_/A hold323/X vssd1 vssd1 vccd1 vccd1 _13340_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12042_ hold314/A _12175_/A2 _12109_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _12042_/X
+ sky130_fd_sc_hd__a31o_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _13211_/A _12943_/B _12853_/X vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11656__A1 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__B2 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ hold283/X hold38/X vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08096__B _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11826_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11827_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11757_ _11757_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__nor2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ _10966_/A fanout9/X fanout4/X _10859_/A vssd1 vssd1 vccd1 vccd1 _10709_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11688_ _11325_/B _11506_/B _11856_/A _11687_/X vssd1 vssd1 vccd1 vccd1 _11689_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10639_ _10639_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13358_ _13364_/CLK _13358_/D vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08840__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ _12309_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13289_ _13352_/CLK hold212/X vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07456__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__B1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07852_/A sky130_fd_sc_hd__xor2_2
X_06801_ reg2_val[0] _06794_/B _06801_/B1 _06799_/X vssd1 vssd1 vccd1 vccd1 _06801_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09671__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ _07153_/Y _07944_/B fanout28/X _07128_/Y vssd1 vssd1 vccd1 vccd1 _07782_/B
+ sky130_fd_sc_hd__a22o_1
X_06732_ _10918_/S _06732_/B vssd1 vssd1 vccd1 vccd1 _06879_/D sky130_fd_sc_hd__nor2_2
X_09520_ _09520_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06663_ instruction[32] _06699_/B vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__and2_4
X_09451_ _10937_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__xor2_1
X_06594_ instruction[25] _06699_/B vssd1 vssd1 vccd1 vccd1 _12619_/B sky130_fd_sc_hd__and2_4
X_09382_ _09165_/X _09169_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09068__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ _10942_/A _08440_/B _08441_/A vssd1 vssd1 vccd1 vccd1 _08416_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _08333_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07079__B2 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _11557_/A _11453_/A _07214_/Y vssd1 vssd1 vccd1 vccd1 _07215_/Y sky130_fd_sc_hd__a21oi_4
X_08195_ _08193_/A _08193_/B _08253_/A vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08028__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _07146_/A _07146_/B vssd1 vssd1 vccd1 vccd1 _07146_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07077_ _11446_/A _07077_/B vssd1 vssd1 vccd1 vccd1 _07077_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07366__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _09386_/X _09388_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__mux2_1
X_07979_ _08049_/A _08049_/B _08049_/C vssd1 vssd1 vccd1 vccd1 _08050_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout53_A _07052_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _10990_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _09650_/B _09650_/C _10231_/A vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__a21o_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12659_/A _12656_/Y _12658_/B vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11611_ _11611_/A _11611_/B _11611_/C vssd1 vssd1 vccd1 vccd1 _11612_/C sky130_fd_sc_hd__and3_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _12598_/B _12591_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11542_ _11542_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11473_ _11837_/A fanout22/X fanout14/X fanout61/X vssd1 vssd1 vccd1 vccd1 _11474_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11070__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ hold301/X _13211_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_1
X_10424_ _10420_/Y _10423_/Y _11958_/A vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__mux2_1
X_13143_ hold319/X _13186_/A2 _13142_/X _13143_/B2 vssd1 vssd1 vccd1 vccd1 _13144_/B
+ sky130_fd_sc_hd__a22o_1
X_10355_ _10355_/A _10355_/B vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__xor2_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13074_ _12310_/A _12797_/B hold45/X vssd1 vssd1 vccd1 vccd1 _13335_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__11326__B1 _11451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ _09722_/X _09725_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _10286_/X sky130_fd_sc_hd__mux2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ _06848_/B _12024_/Y _12025_/S vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13217__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ hold65/X hold302/X vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12858_ hold314/A hold120/X vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12054__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ _11809_/A _11809_/B _11809_/C _11809_/D vssd1 vssd1 vccd1 vccd1 _12020_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12054__B2 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ hold46/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__or2_1
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__A1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ _07000_/A _07000_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__nand2_8
XANTENNA__12357__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08570__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08951_ _08952_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _09064_/A sky130_fd_sc_hd__nor2_1
X_07902_ _07902_/A _07902_/B _07899_/Y vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08882_ _07569_/A _07569_/B _07566_/A vssd1 vssd1 vccd1 vccd1 _08894_/A sky130_fd_sc_hd__a21oi_1
X_07833_ _08573_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07834_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13127__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A _07043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _07760_/Y _07829_/B _07759_/Y vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__a21o_2
X_06715_ _11231_/A _07243_/A vssd1 vssd1 vccd1 vccd1 _06716_/B sky130_fd_sc_hd__nor2_1
X_09503_ _09503_/A _09503_/B vssd1 vssd1 vccd1 vccd1 _09505_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07695_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07695_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10843__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06646_ _12772_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__xnor2_2
X_09434_ _10288_/S _09433_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _09434_/Y sky130_fd_sc_hd__o21ai_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06577_ instruction[13] _06575_/X _06576_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09365_ _09365_/A _09365_/B vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_30 reg2_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_41 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _09462_/B _09296_/B vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__nor2_1
X_08316_ _08594_/A2 _08551_/A2 _08551_/B1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08317_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_52 reg2_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08247_ _08256_/A _08256_/B vssd1 vssd1 vccd1 vccd1 _08247_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09749__B1 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__B2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A1 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _08178_/A _08178_/B vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ _07129_/A _07129_/B vssd1 vssd1 vccd1 vccd1 _07129_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08972__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10315_/A _10140_/B _10140_/C vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__or3_1
XANTENNA__07775__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _07402_/B _10222_/A2 _10712_/A fanout40/X vssd1 vssd1 vccd1 vccd1 _10072_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06983__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _11092_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10975_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10834__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12712_ _12716_/C _12711_/B _12709_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _12641_/Y _12643_/B vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__nand2b_2
X_12574_ _12574_/A _12574_/B _12574_/C vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__or3_1
XFILLER_0_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ _11879_/A2 _11623_/B hold295/A vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11456_ _11456_/A _11988_/A _11566_/A vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__nor3_1
XANTENNA__07215__A1 _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11387_ _11387_/A _11387_/B vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__xnor2_1
X_10407_ _10315_/X _10406_/X _09148_/Y vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13126_ _13126_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13126_/Y sky130_fd_sc_hd__xnor2_1
X_10338_ _07072_/B fanout7/X _10234_/A vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ hold117/X _13071_/A2 _13071_/B1 hold137/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold138/A sky130_fd_sc_hd__o221a_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12008_ _12083_/B _12008_/B vssd1 vssd1 vccd1 vccd1 _12011_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10269_ _09703_/X _09855_/X _09856_/X _10319_/B _10650_/A vssd1 vssd1 vccd1 vccd1
+ _10270_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_0_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08191__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07480_ _07480_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _12339_/A1 _10310_/A _10310_/B _09147_/Y _11889_/A1 vssd1 vssd1 vccd1 vccd1
+ _09150_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09443__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ _08105_/A _08105_/B _08095_/X vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__a21oi_2
X_09081_ _10081_/A _09081_/B vssd1 vssd1 vccd1 vccd1 _09083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _09468_/B2 _08184_/B fanout32/X _08591_/B1 vssd1 vssd1 vccd1 vccd1 _08033_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11538__B1 _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout103_A _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _09836_/A _09836_/B _09834_/X vssd1 vssd1 vccd1 vccd1 _09985_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07757__A2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08934_ _09766_/A _08934_/B vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08706__A1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 _09900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _08865_/A _08865_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10070__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07816_ _08605_/A _07891_/B _07891_/C vssd1 vssd1 vccd1 vccd1 _07818_/C sky130_fd_sc_hd__and3_1
X_08796_ _08803_/A _08796_/B _08796_/C vssd1 vssd1 vccd1 vccd1 _08797_/B sky130_fd_sc_hd__nand3_1
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10816__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _06973_/Y fanout62/X fanout56/X _06973_/A vssd1 vssd1 vccd1 vccd1 _07679_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06629_ _12381_/A _06858_/A vssd1 vssd1 vccd1 vccd1 _06656_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ _12415_/A _12785_/A _09418_/C vssd1 vssd1 vccd1 vccd1 _09417_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _09349_/A _09349_/B vssd1 vssd1 vccd1 vccd1 _09348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11310_ _11311_/B _11311_/A vssd1 vssd1 vccd1 vccd1 _11310_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ reg1_val[28] _12341_/C vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11241_ _11529_/B _11347_/B hold210/A vssd1 vssd1 vccd1 vccd1 _11242_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11172_ _11172_/A _11172_/B vssd1 vssd1 vccd1 vccd1 _11173_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10201__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_30_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07381__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ _06978_/X fanout31/X fanout29/X _07012_/Y vssd1 vssd1 vccd1 vccd1 _10957_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12619__B _12619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ _10646_/A _10763_/X _10765_/B vssd1 vssd1 vccd1 vccd1 _10887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06617__B _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ reg1_val[2] _12627_/B vssd1 vssd1 vccd1 vccd1 _12626_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09425__A2 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ _12610_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__or2_1
XANTENNA__09928__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_11508_ _11686_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__xnor2_4
X_12488_ _12488_/A _12488_/B _12488_/C vssd1 vssd1 vccd1 vccd1 _12489_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ hold281/A _11439_/B vssd1 vssd1 vccd1 vccd1 _11439_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13109_ _13109_/A hold310/X vssd1 vssd1 vccd1 vccd1 _13344_/D sky130_fd_sc_hd__and2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09155__S _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _09670_/A _06980_/B vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__xnor2_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _08650_/A _08659_/S vssd1 vssd1 vccd1 vccd1 _08651_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07601_ fanout50/X _10463_/B2 _10228_/A _09659_/B2 vssd1 vssd1 vccd1 vccd1 _07602_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08581_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08581_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07124__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07532_ _08553_/A2 fanout24/X _07264_/X _08096_/B vssd1 vssd1 vccd1 vccd1 _07533_/B
+ sky130_fd_sc_hd__o22a_1
X_07463_ _07519_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/A sky130_fd_sc_hd__and2_1
XFILLER_0_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09202_ _09200_/X _09201_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _08650_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _07492_/B sky130_fd_sc_hd__xnor2_2
X_09133_ _09134_/A _09134_/B vssd1 vssd1 vccd1 vccd1 _09133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11223__A2 _11258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10431__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ _09064_/A _09064_/B _09064_/C vssd1 vssd1 vccd1 vccd1 _09065_/B sky130_fd_sc_hd__or3_1
XFILLER_0_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08015_ _08445_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13079__C fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12280__A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__and2_1
X_09897_ reg1_val[4] _07097_/C _11966_/B _09890_/X _09896_/X vssd1 vssd1 vccd1 vccd1
+ _09898_/A sky130_fd_sc_hd__a311o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ _07660_/A _07660_/B _08916_/X vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__a21o_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08852_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07363__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _08787_/A _08778_/C _08786_/B vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__a21o_1
X_11790_ hold302/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10810_ _10810_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_39_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10741_ _10742_/A _10742_/B vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__and2_1
XANTENNA__07130__A3 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10670__B1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12411_/Y sky130_fd_sc_hd__nand2_1
X_10672_ hold213/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ reg1_val[28] _12341_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12273_ _12271_/B _12273_/B vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09764__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11224_ _11863_/A _08741_/X _08743_/X vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ _11155_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09591__A1 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__xor2_1
X_10106_ _09927_/A _09926_/B _09924_/X vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__a21o_1
X_10037_ _12490_/S _10033_/X _10034_/X _10036_/Y vssd1 vssd1 vccd1 vccd1 dest_val[5]
+ sky130_fd_sc_hd__a22o_4
X_11988_ _11988_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11992_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ _10939_/A _10939_/B vssd1 vssd1 vccd1 vccd1 _10948_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11989__B1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11253__B _11253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08854__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09004__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10661__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__and2_1
XFILLER_0_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12953__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11913__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10613__A _10613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06963_ _06963_/A _06963_/B _06963_/C vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__nand3_4
X_09751_ _09226_/Y _09742_/X _09743_/Y _09750_/X _09735_/X vssd1 vssd1 vccd1 vccd1
+ _09751_/X sky130_fd_sc_hd__a311o_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _08702_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__xnor2_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06894_ _06922_/B dest_pred_val _06908_/C vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
X_09682_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08633_ _12785_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout268_A _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08564_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _08564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout47 _07111_/Y vssd1 vssd1 vccd1 vccd1 _07814_/B sky130_fd_sc_hd__buf_6
XFILLER_0_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout14 fanout15/X vssd1 vssd1 vccd1 vccd1 fanout14/X sky130_fd_sc_hd__buf_6
Xfanout36 fanout37/X vssd1 vssd1 vccd1 vccd1 _07155_/A sky130_fd_sc_hd__clkbuf_8
Xfanout25 _07215_/Y vssd1 vssd1 vccd1 vccd1 fanout25/X sky130_fd_sc_hd__buf_6
XFILLER_0_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08845__B1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ _08566_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08499_/A sky130_fd_sc_hd__xnor2_1
Xfanout69 _09930_/A vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout58 _07013_/X vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__buf_8
X_07446_ _07446_/A _07446_/B vssd1 vssd1 vccd1 vccd1 _07525_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07377_ _09630_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07379_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08073__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08073__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ _09117_/A _09117_/B vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09047_ _09930_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06720__B _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _11169_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout83_A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__A1 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__B2 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12960_ _12978_/A hold262/X vssd1 vssd1 vccd1 vccd1 _13278_/D sky130_fd_sc_hd__and2_1
XANTENNA__11132__A1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _12001_/B _11911_/B vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__and2_1
XFILLER_0_99_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12891_ hold46/X hold265/X vssd1 vssd1 vccd1 vccd1 _13087_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10669__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A _11842_/B vssd1 vssd1 vccd1 vccd1 _11843_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09089__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11937_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11808_/D sky130_fd_sc_hd__xor2_2
XFILLER_0_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10726_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11199__A1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ _11863_/A _11809_/A _10810_/A _11889_/A1 vssd1 vssd1 vccd1 vccd1 _10655_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _13374_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12324_/X _12325_/B vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__nand2b_1
X_10586_ _11296_/B _10586_/B vssd1 vssd1 vccd1 vccd1 _10587_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12256_ _12256_/A _12256_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12632__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _11207_/A _11207_/B vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__xnor2_2
X_12187_ curr_PC[26] _12124_/C _06908_/C vssd1 vssd1 vccd1 vccd1 _12187_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08367__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _11125_/A _07251_/A _12395_/A1 _11137_/X vssd1 vssd1 vccd1 vccd1 _11138_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09316__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__B2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _11172_/A _11069_/B vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11264__A _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ _07300_/A _07300_/B vssd1 vssd1 vccd1 vccd1 _10466_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11977__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08573__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ _09941_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08282_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12807__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ _08445_/A vssd1 vssd1 vccd1 vccd1 _10735_/A sky130_fd_sc_hd__inv_6
XFILLER_0_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07162_ _11125_/A _11231_/A reg1_val[16] _07121_/C _07093_/A vssd1 vssd1 vccd1 vccd1
+ _07164_/B sky130_fd_sc_hd__o41a_2
XANTENNA__06805__B _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ _07093_/A _07120_/C vssd1 vssd1 vccd1 vccd1 _07095_/C sky130_fd_sc_hd__and2_1
XFILLER_0_42_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 _06901_/Y vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__buf_4
XANTENNA__09555__A1 _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _12175_/A2 vssd1 vssd1 vccd1 vccd1 _11879_/A2 sky130_fd_sc_hd__buf_4
XANTENNA__11362__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__B2 _07211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__and2_1
Xfanout215 _07152_/A vssd1 vssd1 vccd1 vccd1 _10148_/S sky130_fd_sc_hd__buf_2
Xfanout237 _06973_/Y vssd1 vssd1 vccd1 vccd1 _08551_/B2 sky130_fd_sc_hd__buf_6
XFILLER_0_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout259 _06564_/A vssd1 vssd1 vccd1 vccd1 _13204_/B2 sky130_fd_sc_hd__buf_4
Xfanout248 _06908_/C vssd1 vssd1 vccd1 vccd1 _12053_/A1 sky130_fd_sc_hd__clkbuf_16
X_07995_ _07995_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__13103__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _09729_/X _09731_/X _09732_/Y _11958_/A vssd1 vssd1 vccd1 vccd1 _09734_/X
+ sky130_fd_sc_hd__a31o_1
X_06946_ _12621_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07318__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _11611_/A _06877_/B _11428_/A _11333_/A vssd1 vssd1 vccd1 vccd1 _06884_/C
+ sky130_fd_sc_hd__and4_1
X_09665_ _11169_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__xnor2_2
X_08616_ _08616_/A _08616_/B vssd1 vssd1 vccd1 vccd1 _08718_/A sky130_fd_sc_hd__nor2_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _11238_/S _09596_/B vssd1 vssd1 vccd1 vccd1 _09596_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08547_ _08548_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08561_/A sky130_fd_sc_hd__or2_1
XFILLER_0_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11902__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09491__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12717__B _12717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ fanout79/X _10463_/B2 _10228_/A fanout75/X vssd1 vssd1 vccd1 vccd1 _07430_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06715__B _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10440_ _12490_/S _10686_/C _10439_/Y _10437_/X vssd1 vssd1 vccd1 vccd1 dest_val[8]
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ _10369_/Y _10371_/B vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09794__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A1 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12110_ _12175_/A2 _12173_/B hold269/A vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__a21oi_1
X_13090_ hold322/X _13222_/A2 _13089_/X _13095_/B2 vssd1 vssd1 vccd1 vccd1 hold323/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ _12175_/A2 _12109_/B hold314/A vssd1 vssd1 vccd1 vccd1 _12041_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__A1 _09370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 hold329/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__buf_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10561__C1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ _12853_/X _12943_/B vssd1 vssd1 vccd1 vccd1 _13211_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11656__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08521__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ hold303/X hold32/X vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__nand2b_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11826_/A _11826_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__or2_1
XFILLER_0_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ _11756_/A _11756_/B _11756_/C vssd1 vssd1 vccd1 vccd1 _11757_/B sky130_fd_sc_hd__and3_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__or2_1
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12627__B _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ _11503_/X _11856_/A _11685_/X vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11023__S _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _10639_/B _10639_/A vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10919__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13030__A1 _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ _13364_/CLK _13357_/D vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ _12525_/S _10441_/X _10539_/X _10568_/X vssd1 vssd1 vccd1 vccd1 dest_val[9]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_11_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13288_ _13352_/CLK hold236/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__dfxtp_1
X_12308_ _12404_/B _12308_/B vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12239_ hold329/A _12239_/B vssd1 vssd1 vccd1 vccd1 _12296_/B sky130_fd_sc_hd__or2_1
X_06800_ reg2_val[0] _06794_/B _06801_/B1 _06799_/X vssd1 vssd1 vccd1 vccd1 _09101_/A
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__08568__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ _09795_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__xnor2_2
X_06731_ reg1_val[12] _07175_/A vssd1 vssd1 vccd1 vccd1 _06732_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09163__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12844__A1 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _07402_/B _10326_/A _09450_/B1 fanout41/X vssd1 vssd1 vccd1 vccd1 _09451_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06662_ _11966_/A _06662_/B vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__nor2_2
X_08401_ _08440_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08441_/A sky130_fd_sc_hd__nand2_1
X_06593_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06593_/X sky130_fd_sc_hd__or4bb_4
X_09381_ _09162_/X _09164_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09381_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07079__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _08353_/A _08353_/B _08331_/A vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11280__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08263_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08263_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07214_ _07192_/A _07192_/B _07210_/B _11361_/A vssd1 vssd1 vccd1 vccd1 _07214_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout133_A _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__or2_1
XANTENNA__08028__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07145_ _07145_/A _07146_/B vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__xnor2_4
X_07076_ _11446_/A _07077_/B vssd1 vssd1 vccd1 vccd1 _07076_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__11169__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__A0 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ _09630_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _08049_/C sky130_fd_sc_hd__xnor2_1
X_06929_ _09227_/B _09238_/B vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__or2_2
X_09717_ _09715_/X _09716_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07382__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A _08517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout46_A _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _09648_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _09650_/C sky130_fd_sc_hd__or3_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__C1 _12030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09579_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12577_/Y _12598_/C _12600_/B vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__o21ai_4
X_11610_ _11611_/B _11611_/C _11611_/A vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _11718_/C _11540_/Y _12525_/S _11538_/X vssd1 vssd1 vccd1 vccd1 dest_val[18]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_53_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ _13211_/A _13211_/B vssd1 vssd1 vccd1 vccd1 _13211_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12463__A _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _11131_/A _10281_/X _10422_/X vssd1 vssd1 vccd1 vccd1 _10423_/Y sky130_fd_sc_hd__a21oi_2
X_13142_ hold277/X _13141_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__mux2_1
X_10354_ _10933_/A _10354_/B vssd1 vssd1 vccd1 vccd1 _10355_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11326__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ hold44/X _13108_/B2 _13222_/A2 hold24/X rst vssd1 vssd1 vccd1 vccd1 hold45/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10285_ _10283_/X _10284_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10285_/X sky130_fd_sc_hd__mux2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _11951_/A _11949_/X _11966_/A vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09772__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__A1 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ _13175_/A _12925_/B _12863_/X vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ _12855_/X _12857_/B vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12039__C1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ _11808_/A _11808_/B _11808_/C _11808_/D vssd1 vssd1 vccd1 vccd1 _12020_/A
+ sky130_fd_sc_hd__nor4_1
XANTENNA__12054__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ _07128_/Y _13078_/B2 hold166/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13243_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _12065_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09158__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07769__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08950_ _10231_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__xnor2_1
X_07901_ _07897_/A _07897_/B _07897_/C vssd1 vssd1 vccd1 vccd1 _07901_/X sky130_fd_sc_hd__a21o_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__xor2_1
X_07832_ _08594_/A2 fanout79/X fanout75/X _08572_/A2 vssd1 vssd1 vccd1 vccd1 _07833_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09503_/B sky130_fd_sc_hd__xor2_1
X_07763_ _08624_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07829_/B sky130_fd_sc_hd__xor2_1
X_06714_ _11231_/A _07243_/A vssd1 vssd1 vccd1 vccd1 _11246_/S sky130_fd_sc_hd__and2_1
X_07694_ _07789_/A _07789_/B _07691_/Y vssd1 vssd1 vccd1 vccd1 _07715_/B sky130_fd_sc_hd__a21o_1
X_06645_ instruction[41] _06908_/A _06600_/B _06643_/X vssd1 vssd1 vccd1 vccd1 _07127_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout250_A _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _11235_/S _09432_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _09433_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11452__A _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ _09365_/B _09365_/A vssd1 vssd1 vccd1 vccd1 _09364_/Y sky130_fd_sc_hd__nand2b_1
X_06576_ instruction[20] _06922_/B vssd1 vssd1 vccd1 vccd1 _06576_/X sky130_fd_sc_hd__or2_1
XANTENNA__12045__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08315_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__or2_1
XFILLER_0_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 reg2_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 reg2_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09294_/B _09295_/B vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_53 reg2_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 reg1_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08246_ _08271_/A _08271_/B _08235_/Y vssd1 vssd1 vccd1 vccd1 _08256_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _09941_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10359__A2 _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _09725_/S _07129_/B vssd1 vssd1 vccd1 vccd1 _07128_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07377__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07059_ _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__and2_2
X_10070_ _11296_/B _10070_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08185__A0 _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__A1 _07179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ _10972_/A _10972_/B _10972_/C vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__and3_1
XANTENNA__10819__B1 _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _12716_/C _12711_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xor2_4
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ reg1_val[5] _12642_/B vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__B1 _09436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ _12573_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11524_ hold281/A hold320/A _11524_/C vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__or3_1
XFILLER_0_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11455_ _11456_/A _11988_/A _11566_/A vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07053__C_N _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10406_/A _10650_/C vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__xor2_2
X_11386_ _11386_/A _11988_/A vssd1 vssd1 vccd1 vccd1 _11387_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_104_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _13125_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__nand2_1
X_10337_ _10735_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _07192_/C _13078_/B2 hold118/X vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__o21a_1
X_10268_ _09993_/X _10125_/X _10126_/X vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__a21oi_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _12007_/A _12007_/B _12007_/C vssd1 vssd1 vccd1 vccd1 _12008_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08176__B1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08479__A1 _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ hold35/X hold305/X vssd1 vssd1 vccd1 vccd1 _13135_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08846__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _08184_/B _11296_/A _11188_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _09081_/B
+ sky130_fd_sc_hd__o22a_1
X_08100_ _08100_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12815__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08031_ _08083_/A _08083_/B _08027_/X vssd1 vssd1 vccd1 vccd1 _08035_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11538__B2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ _09824_/A _09824_/B _09822_/Y vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08933_ _07539_/B _09450_/B1 _07263_/Y fanout37/X vssd1 vssd1 vccd1 vccd1 _08934_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09903__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__xnor2_2
X_07815_ _07000_/A _07000_/B _06973_/A vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__a21oi_1
X_08795_ _08796_/B _08796_/C _08803_/A vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09667__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11182__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _09419_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09418_/C sky130_fd_sc_hd__xnor2_1
X_07677_ _07687_/B _07687_/A vssd1 vssd1 vccd1 vccd1 _07677_/X sky130_fd_sc_hd__and2b_1
X_06628_ _06626_/X _06628_/B vssd1 vssd1 vccd1 vccd1 _06858_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09347_ _09107_/A _09107_/B _09105_/Y vssd1 vssd1 vccd1 vccd1 _09349_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _09278_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _09941_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08231_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11240_ hold210/A _11529_/B _11347_/B vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ fanout33/X fanout12/X fanout6/X fanout35/X vssd1 vssd1 vccd1 vccd1 _11172_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10201__A1 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__B2 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10122_/X sky130_fd_sc_hd__and2_1
XFILLER_0_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07381__B2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A1 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10955_ _10955_/A _10955_/B vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08330__B1 _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__or2_2
XFILLER_0_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12625_ _12624_/A _12624_/B _12623_/B vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ _12610_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12965__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _11114_/B _11506_/X _11505_/X vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ _12488_/A _12488_/B _12488_/C vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11438_ hold320/A _11524_/C _11879_/A2 vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__o21a_1
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11381_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ hold309/X _13222_/A2 _13107_/X _13108_/B2 vssd1 vssd1 vccd1 vccd1 hold310/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07745__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ hold141/X _13071_/A2 _13053_/B1 hold195/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold196/A sky130_fd_sc_hd__o221a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08580_ _08580_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08584_/B sky130_fd_sc_hd__xor2_1
X_07600_ _07600_/A _07600_/B vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09649__B1 _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _07531_/A _07531_/B vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07124__A1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08321__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07462_ _09795_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07519_/B sky130_fd_sc_hd__xnor2_1
X_09201_ _11125_/A reg1_val[17] _09560_/A vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__mux2_1
X_07393_ _09297_/B2 fanout56/X _09297_/A1 fanout62/X vssd1 vssd1 vccd1 vccd1 _07394_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09132_ _09010_/A _09010_/B _09011_/X vssd1 vssd1 vccd1 vccd1 _09134_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09063_ _09064_/A _09064_/B _09064_/C vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08014_ _08926_/B1 _10227_/B1 _10463_/A1 _08521_/A2 vssd1 vssd1 vccd1 vccd1 _08015_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _11359_/A _09965_/B vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11177__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ _12171_/A _06924_/Y _09895_/X _09595_/B _06780_/A vssd1 vssd1 vccd1 vccd1
+ _09896_/X sky130_fd_sc_hd__a32o_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ _07660_/A _07660_/B _08702_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08916_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09870__A _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08847_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07363__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _08786_/B _08787_/A _08778_/C vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07390__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__xor2_4
X_10740_ _10578_/A _10578_/B _10583_/A vssd1 vssd1 vccd1 vccd1 _10742_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07130__A4 _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _11238_/S _10669_/X _10670_/X _09243_/B vssd1 vssd1 vccd1 vccd1 _10671_/X
+ sky130_fd_sc_hd__a211o_1
X_12410_ _12365_/A _12364_/A _12410_/S vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ reg1_val[28] reg1_val[29] _12341_/C vssd1 vssd1 vccd1 vccd1 _12421_/C sky130_fd_sc_hd__and3_1
XANTENNA__10422__A1 _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ _12324_/B _12323_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12272_/Y sky130_fd_sc_hd__o21ai_1
X_11223_ _11153_/X _11258_/B _11222_/Y vssd1 vssd1 vccd1 vccd1 _11253_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_31_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12471__A _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _11386_/A fanout9/A fanout5/X _11296_/A vssd1 vssd1 vccd1 vccd1 _11155_/B
+ sky130_fd_sc_hd__o22a_1
X_11085_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11085_/Y sky130_fd_sc_hd__nand2b_1
X_10105_ _10105_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10036_ _12490_/S _10172_/B vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11815__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap109_A _10490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ fanout67/X fanout9/X fanout4/X _12059_/A vssd1 vssd1 vccd1 vccd1 _11988_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ _10939_/A _10939_/B vssd1 vssd1 vccd1 vccd1 _11045_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11989__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11989__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08854__A1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08854__B2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10869_ _10743_/A _10743_/B _10741_/X vssd1 vssd1 vccd1 vccd1 _10874_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ reg1_val[26] curr_PC[26] _12615_/S vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12402__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12539_ _11231_/A curr_PC[15] _12615_/S vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__A1 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11913__B2 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06962_ _06963_/A _06963_/B _06963_/C vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__and3_4
X_09750_ _09743_/A _09228_/Y _09237_/Y _09745_/X _09749_/X vssd1 vssd1 vccd1 vccd1
+ _09750_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _09681_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__xnor2_2
X_08701_ _08702_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__xor2_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ instruction[2] _06893_/B _06893_/C vssd1 vssd1 vccd1 vccd1 _06893_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__11725__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _08632_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _08644_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _08586_/A _08563_/B vssd1 vssd1 vccd1 vccd1 _08578_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ _07514_/A _07719_/A vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08845__A1 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ _08551_/B2 _08521_/A2 _08926_/B1 _06875_/A vssd1 vssd1 vccd1 vccd1 _08495_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout15 _07581_/Y vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__clkbuf_8
Xfanout37 _07154_/X vssd1 vssd1 vccd1 vccd1 fanout37/X sky130_fd_sc_hd__clkbuf_8
X_07445_ _10231_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08845__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout26 fanout27/X vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__buf_6
Xfanout59 _07013_/X vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__buf_4
Xfanout48 _11359_/A vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ _07101_/Y fanout28/X _07263_/Y _07944_/B vssd1 vssd1 vccd1 vccd1 _07377_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08073__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09115_ _09827_/A _09115_/B vssd1 vssd1 vccd1 vccd1 _09117_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _09815_/A _07347_/B fanout15/X _09675_/A vssd1 vssd1 vccd1 vccd1 _09047_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12291__A _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09948_ fanout57/X fanout77/X fanout73/X _11837_/A vssd1 vssd1 vccd1 vccd1 _09949_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__10015__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09325__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09191_/X _09213_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__mux2_1
X_11910_ _11910_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__nand2_1
X_12890_ _13083_/A _13083_/B _12887_/X vssd1 vssd1 vccd1 vccd1 _13088_/A sky130_fd_sc_hd__a21o_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _11841_/B _11841_/C vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__nor3_1
XANTENNA__10891__A1 _10406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09089__A1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__B2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11007_/B _11415_/Y _12087_/A _11769_/Y _12088_/A vssd1 vssd1 vccd1 vccd1
+ _11773_/B sky130_fd_sc_hd__o311a_2
XANTENNA__12093__B1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _11557_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10724_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ _11863_/A _11809_/A _10810_/A vssd1 vssd1 vccd1 vccd1 _10654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11199__A2 _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ _13375_/CLK hold156/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
X_10585_ _10859_/A fanout9/A fanout5/X _10585_/B2 vssd1 vssd1 vccd1 vccd1 _10586_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12324_ _12324_/A _12324_/B _12324_/C _12406_/A vssd1 vssd1 vccd1 vccd1 _12324_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _12255_/A _12255_/B _12255_/C vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__and3_1
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11206_ _11207_/B _11207_/A vssd1 vssd1 vccd1 vccd1 _11206_/Y sky130_fd_sc_hd__nand2b_1
X_12186_ curr_PC[25] curr_PC[26] _12186_/C vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__and3_1
X_11137_ _09886_/B _12394_/A1 _11137_/S vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09316__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ fanout33/X fanout13/X fanout12/X fanout35/X vssd1 vssd1 vccd1 vccd1 _11069_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11545__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10019_ hold317/A _10156_/C _10158_/A2 vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_59_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__or2_4
XFILLER_0_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07161_ _11125_/A _11231_/A _07121_/C _07093_/A vssd1 vssd1 vccd1 vccd1 _07168_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12823__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ reg1_val[22] _07092_/B vssd1 vssd1 vccd1 vccd1 _07120_/C sky130_fd_sc_hd__or2_1
XFILLER_0_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13000__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _09385_/S vssd1 vssd1 vccd1 vccd1 _09402_/S sky130_fd_sc_hd__clkbuf_8
Xfanout227 _11029_/A2 vssd1 vssd1 vccd1 vccd1 _12175_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11362__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ _10081_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__xnor2_1
Xfanout216 _06790_/X vssd1 vssd1 vccd1 vccd1 _07152_/A sky130_fd_sc_hd__buf_4
Xfanout238 _09670_/A vssd1 vssd1 vccd1 vccd1 _08566_/A sky130_fd_sc_hd__buf_12
XFILLER_0_1_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout249 _06892_/X vssd1 vssd1 vccd1 vccd1 _06908_/C sky130_fd_sc_hd__buf_6
X_07994_ _07939_/X _08059_/B _07938_/X vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__a21o_2
XANTENNA_fanout280_A _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _09731_/X _09732_/Y _09729_/X vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__a21oi_1
X_06945_ _12619_/A reg1_val[31] _12415_/A vssd1 vssd1 vccd1 vccd1 _06947_/B sky130_fd_sc_hd__and3_4
XANTENNA__07318__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ _09219_/A _09396_/S vssd1 vssd1 vccd1 vccd1 _06876_/Y sky130_fd_sc_hd__nor2_1
X_09664_ fanout60/X fanout77/X fanout73/X fanout52/X vssd1 vssd1 vccd1 vccd1 _09665_/B
+ sky130_fd_sc_hd__o22a_1
X_09595_ _09595_/A _09595_/B vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__nand2_1
X_08615_ _08595_/X _08613_/Y _08612_/Y _08603_/Y vssd1 vssd1 vccd1 vccd1 _08616_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08548_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09491__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09491__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07428_ _07428_/A _07428_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07359_ _07359_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07361_/A sky130_fd_sc_hd__or2_1
XFILLER_0_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10370_ _10370_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09794__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06731__B _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ _09029_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _09030_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ hold289/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12109_/B sky130_fd_sc_hd__or2_1
XANTENNA__09546__A2 _09370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07843__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ hold301/X hold114/X vssd1 vssd1 vccd1 vccd1 _12943_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ hold308/A hold95/X vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _07116_/Y wire8/X _11823_/X _11900_/A vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__a22o_1
X_11755_ _11756_/A _11756_/B _11756_/C vssd1 vssd1 vccd1 vccd1 _11757_/A sky130_fd_sc_hd__a21oi_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10709__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10706_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07493__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__B _06907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ _11686_/A _11767_/A vssd1 vssd1 vccd1 vccd1 _11856_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13030__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356_ _13364_/CLK _13356_/D vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06599__A2 _06591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10568_ _12029_/A _10540_/Y _10541_/X _10567_/X vssd1 vssd1 vccd1 vccd1 _10568_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _10500_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__and2_1
X_13287_ _13287_/CLK _13287_/D vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__dfxtp_1
X_12307_ fanout9/X fanout6/X fanout4/X fanout12/X vssd1 vssd1 vccd1 vccd1 _12308_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12238_ hold242/A _12347_/B _12293_/B vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__11344__A2 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12167_/Y _12169_/B vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07753__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ reg1_val[12] _07175_/A vssd1 vssd1 vccd1 vccd1 _10918_/S sky130_fd_sc_hd__and2_1
XANTENNA__12844__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ reg1_val[23] _07016_/A vssd1 vssd1 vccd1 vccd1 _06662_/B sky130_fd_sc_hd__and2b_1
X_08400_ _09403_/S _08400_/B vssd1 vssd1 vccd1 vccd1 _08440_/B sky130_fd_sc_hd__nor2_1
X_06592_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06908_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09380_ _09378_/X _09379_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09380_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10619__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11280__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__A1 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__xnor2_2
X_07213_ _07213_/A _07213_/B vssd1 vssd1 vccd1 vccd1 _07213_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08028__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11032__A1 _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ _07152_/A _07129_/A _08476_/A _07127_/B _12415_/A vssd1 vssd1 vccd1 vccd1
+ _07146_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10354__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ _07074_/A _06963_/A _06963_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _07077_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07139__S _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07977_ _07975_/Y _07977_/B _08049_/A vssd1 vssd1 vccd1 vccd1 _08049_/B sky130_fd_sc_hd__nand3b_2
X_06928_ _09227_/B _09238_/B vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__nor2_2
X_09716_ _09382_/X _09385_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09716_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12710__A2_N _07089_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06859_ _06852_/Y _06858_/Y _12285_/A vssd1 vssd1 vccd1 vccd1 _06859_/X sky130_fd_sc_hd__a21o_1
X_09647_ _07593_/A _07593_/B _08590_/B vssd1 vssd1 vccd1 vccd1 _09650_/B sky130_fd_sc_hd__a21o_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09576_/Y _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__nand2b_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08529_ _08549_/A _08549_/B _08525_/X vssd1 vssd1 vccd1 vccd1 _08536_/B sky130_fd_sc_hd__o21a_1
XANTENNA__06726__B _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ curr_PC[18] _11539_/B _06908_/C vssd1 vssd1 vccd1 vccd1 _11540_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11471_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ _13226_/A _13210_/B vssd1 vssd1 vccd1 vccd1 _13365_/D sky130_fd_sc_hd__and2_1
X_10422_ _10902_/A _09214_/X _10421_/X _11237_/S vssd1 vssd1 vccd1 vccd1 _10422_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13141_ _13141_/A _13141_/B vssd1 vssd1 vccd1 vccd1 _13141_/Y sky130_fd_sc_hd__xnor2_1
X_10353_ _07151_/A _07237_/Y _07243_/X _07155_/A vssd1 vssd1 vccd1 vccd1 _10354_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _07346_/B _13072_/A2 hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o21a_1
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12023_ _12278_/A _12021_/Y _12022_/X vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__o21a_1
X_10284_ _09719_/X _09724_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12826__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12925_ _12863_/X _12925_/B vssd1 vssd1 vccd1 vccd1 _13175_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10837__B2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__A1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ hold269/X hold98/X vssd1 vssd1 vccd1 vccd1 _12857_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07702__B2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11542__B _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _06908_/C _11803_/X _11806_/X vssd1 vssd1 vccd1 vccd1 dest_val[21] sky130_fd_sc_hd__o21ai_4
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ hold165/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__or2_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11738_ _07155_/Y _12257_/A _12309_/A _07151_/Y vssd1 vssd1 vccd1 vccd1 _11739_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ _11670_/B _11670_/A vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ _13341_/CLK _13339_/D vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__A1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__B2 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07186__C _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10902__A _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ _07897_/A _07897_/B _07897_/C vssd1 vssd1 vccd1 vccd1 _07902_/B sky130_fd_sc_hd__a21oi_1
X_08880_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__xnor2_1
X_07831_ _08445_/A _07831_/B vssd1 vssd1 vccd1 vccd1 _07834_/A sky130_fd_sc_hd__xnor2_1
X_09501_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__nor2_1
X_07762_ _08649_/B fanout52/X fanout50/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _07763_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06713_ _06908_/A _06591_/X _06706_/A _06712_/X vssd1 vssd1 vccd1 vccd1 _07243_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_78_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07693_ _07693_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _07789_/B sky130_fd_sc_hd__xor2_1
X_06644_ _06567_/Y _06600_/Y _06643_/X vssd1 vssd1 vccd1 vccd1 _06644_/X sky130_fd_sc_hd__o21ba_2
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _10148_/S _09431_/X _09249_/B vssd1 vssd1 vccd1 vccd1 _09432_/X sky130_fd_sc_hd__o21a_1
X_06575_ _06893_/C _06893_/B instruction[2] vssd1 vssd1 vccd1 vccd1 _06575_/X sky130_fd_sc_hd__or3b_4
XANTENNA__11452__B _11809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ _09363_/A _09363_/B vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10349__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11789__C1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _08314_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07457__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 reg2_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _07078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _09295_/B _09294_/B vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_54 reg2_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08245_ _08300_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08271_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09749__A2 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _08619_/B2 _08354_/A2 _10585_/B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08177_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10359__A3 _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ _12415_/A _07127_/B _08476_/A vssd1 vssd1 vccd1 vccd1 _07129_/B sky130_fd_sc_hd__and3_2
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _07058_/A _07068_/B _07058_/C vssd1 vssd1 vccd1 vccd1 _07060_/B sky130_fd_sc_hd__or3_4
XFILLER_0_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06735__A2 _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06829__A_N _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10972_/A _10972_/B _10972_/C vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _12767_/B _07089_/C _12716_/A _12716_/B vssd1 vssd1 vccd1 vccd1 _12711_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07696__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ reg1_val[5] _12642_/B vssd1 vssd1 vccd1 vccd1 _12641_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09113__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _12616_/A _12572_/B vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12441__A0 _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ _11034_/X _11522_/Y _12171_/A vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ _07214_/Y wire8/X _11453_/Y _11557_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__a22o_2
XANTENNA__07568__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10650_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11385_ _12310_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__C1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13124_ _13134_/A hold304/X vssd1 vssd1 vccd1 vccd1 _13347_/D sky130_fd_sc_hd__and2_1
X_10336_ _10228_/A fanout13/X fanout11/X _10463_/B2 vssd1 vssd1 vccd1 vccd1 _10337_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__B1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ hold144/A _13055_/A2 _13071_/B1 hold117/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold118/A sky130_fd_sc_hd__o221a_1
X_10267_ _10267_/A _10319_/A _10319_/B _10650_/A vssd1 vssd1 vccd1 vccd1 _10267_/X
+ sky130_fd_sc_hd__or4_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _12007_/A _12007_/B _12007_/C vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11704__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_84_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08479__A2 _08517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _13130_/A _13131_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13136_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ hold71/X _12839_/B vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__B1 _12428_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07439__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08862__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09169__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13364_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__09600__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ _09777_/A _09777_/B _09776_/A vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12831__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11171__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08863_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08863_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08794_ _08789_/A _08789_/B _08789_/C _08790_/A _08705_/A vssd1 vssd1 vccd1 vccd1
+ _08796_/C sky130_fd_sc_hd__a311o_2
X_07814_ _12785_/A _07814_/B vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10778__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ _08445_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09667__B2 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ hold285/A hold321/A _06942_/Y _12433_/A1 _09414_/Y vssd1 vssd1 vccd1 vccd1
+ _09415_/X sky130_fd_sc_hd__a311o_1
X_07676_ _07736_/A _07675_/Y _07671_/Y vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06627_ _07029_/A reg1_val[27] vssd1 vssd1 vccd1 vccd1 _06628_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _09277_/A _09277_/B _09277_/C vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__and3_1
XFILLER_0_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ _08619_/B2 _10585_/B2 _10067_/A1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08229_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__xor2_2
X_11170_ _11170_/A _11170_/B vssd1 vssd1 vccd1 vccd1 _11173_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10201__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _10121_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06651__A_N _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10052_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07381__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10955_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__and3_1
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xor2_4
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12555_ reg1_val[18] curr_PC[18] _12615_/S vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06914__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__and2_1
XFILLER_0_81_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12178__C1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ _12495_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12488_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11437_ _09196_/S _11132_/Y _11143_/Y _09223_/Y _11436_/X vssd1 vssd1 vccd1 vccd1
+ _11437_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11368_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09594__B1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ hold293/X _13106_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
X_10319_ _10319_/A _10319_/B _10650_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _10319_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__12651__B _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _11300_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11299_/X sky130_fd_sc_hd__and2b_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11153__B1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ _10735_/A _13078_/B2 hold142/X vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__o21a_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10900__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07531_/A _07531_/B vssd1 vssd1 vccd1 vccd1 _07541_/B sky130_fd_sc_hd__and2_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07124__A2 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08321__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07461_ _08551_/A2 _08096_/B fanout24/X _07264_/X vssd1 vssd1 vccd1 vccd1 _07462_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ _11231_/A reg1_val[16] _09560_/A vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08592__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07392_ _09670_/A _07392_/B vssd1 vssd1 vccd1 vccd1 _07492_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08085__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ _08999_/A _08999_/B _08997_/Y vssd1 vssd1 vccd1 vccd1 _09134_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _08962_/X _09062_/B vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07832__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_A _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ _08049_/B _08011_/B _08011_/C _08008_/Y vssd1 vssd1 vccd1 vccd1 _08040_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10362__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _07077_/X fanout31/X fanout29/X _07237_/Y vssd1 vssd1 vccd1 vccd1 _09965_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09337__B1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A1 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09895_/X sky130_fd_sc_hd__xor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08915_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _09544_/A sky130_fd_sc_hd__xnor2_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _10081_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08848_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07363__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08777_ _08767_/B _08767_/C _08776_/X vssd1 vssd1 vccd1 vccd1 _08778_/C sky130_fd_sc_hd__a21o_1
X_07728_ _07733_/A _07733_/B _07717_/X vssd1 vssd1 vccd1 vccd1 _07800_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07659_ _07660_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07659_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout21_A _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10665_/Y _10666_/X _12171_/A vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _09329_/A _09329_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__and3_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _12420_/A _08809_/A _08808_/Y _11946_/A _12339_/Y vssd1 vssd1 vccd1 vccd1
+ _12356_/B sky130_fd_sc_hd__a311oi_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07823__B1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ _12271_/A _12271_/B _12271_/C vssd1 vssd1 vccd1 vccd1 _12271_/X sky130_fd_sc_hd__or3_1
XFILLER_0_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _11153_/X _11258_/B _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11153_ _11259_/A _11258_/A _11115_/A vssd1 vssd1 vccd1 vccd1 _11153_/X sky130_fd_sc_hd__o21a_1
X_11084_ _11084_/A _11084_/B vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__xnor2_1
X_10104_ _11052_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__xnor2_4
X_10035_ curr_PC[4] curr_PC[5] _10035_/C vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__and3_1
XANTENNA__08551__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06650__A2_N _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _12131_/A _11986_/B vssd1 vssd1 vccd1 vccd1 _11995_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07106__A2 _12717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10937_ _10937_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11989__A2 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08854__A2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _12607_/A _12607_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _10729_/A _10729_/B _10746_/A vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09301__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12646__B _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10949__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ _07179_/A _06940_/B _10797_/Y _10798_/X vssd1 vssd1 vccd1 vccd1 _10800_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12544_/B _12538_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ reg1_val[5] curr_PC[5] _12504_/S vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07756__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11913__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06961_ _07058_/A _07067_/A _11446_/A _07074_/A vssd1 vssd1 vccd1 vccd1 _06963_/C
+ sky130_fd_sc_hd__and4_1
X_09680_ _09680_/A _09680_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__xnor2_2
X_08700_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__xnor2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ instruction[2] _06893_/B _06893_/C vssd1 vssd1 vccd1 vccd1 _06892_/X sky130_fd_sc_hd__and3_1
XANTENNA__10910__A _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _08630_/B _08638_/A _08630_/A vssd1 vssd1 vccd1 vccd1 _08666_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06618__A2_N _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08562_ _08562_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__xnor2_2
X_07513_ _07718_/B _07718_/C _07718_/A vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__a21o_1
X_08493_ _08493_/A _08493_/B vssd1 vssd1 vccd1 vccd1 _08515_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout38 _07539_/B vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__clkbuf_8
Xfanout16 _07302_/X vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__buf_6
Xfanout27 _07211_/X vssd1 vssd1 vccd1 vccd1 fanout27/X sky130_fd_sc_hd__buf_8
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout156_A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07444_ _08590_/B fanout50/X _09659_/B2 _09648_/A vssd1 vssd1 vccd1 vccd1 _07445_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08845__A2 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 _11740_/A vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__buf_12
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07375_ _11361_/A _07375_/B vssd1 vssd1 vccd1 vccd1 _07379_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _07814_/B _10589_/A _09114_/B1 fanout45/X vssd1 vssd1 vccd1 vccd1 _09115_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09045_ _09062_/B _08968_/B _08981_/B _08982_/B _08982_/A vssd1 vssd1 vccd1 vccd1
+ _09061_/A sky130_fd_sc_hd__a32o_2
XFILLER_0_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__A _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _10736_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11916__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout69_A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09876_/X _09877_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__mux2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08497__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__A1 _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ _07600_/A _07600_/B _07598_/X vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__o21ai_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11841_/A _11841_/B _11841_/C vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09089__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11594_/X _11939_/A _11770_/Y vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11651__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10722_ fanout64/X fanout27/X fanout25/X _11980_/A vssd1 vssd1 vccd1 vccd1 _10723_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _10888_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10810_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13372_ _13372_/CLK _13372_/D vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10584_ _10472_/A _10471_/B _10471_/A vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__09797__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _12323_/A _12369_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _12255_/A _12255_/B _12255_/C vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__a21oi_1
X_11205_ _11205_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12185_ _12158_/Y _12159_/X _12184_/X vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08221__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ hold234/A _11529_/B _11239_/B _11242_/A vssd1 vssd1 vccd1 vccd1 _11136_/X
+ sky130_fd_sc_hd__a31o_1
X_11067_ _11184_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10018_ hold222/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10018_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11969_ _09196_/S _10423_/Y _10434_/Y _09223_/Y _11968_/X vssd1 vssd1 vccd1 vccd1
+ _11969_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_58_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09788__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ _07222_/A vssd1 vssd1 vccd1 vccd1 _07160_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ reg1_val[20] reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07092_/B sky130_fd_sc_hd__or2_1
XANTENNA__12792__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09177__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout228 _12349_/A vssd1 vssd1 vccd1 vccd1 _11029_/A2 sky130_fd_sc_hd__buf_2
Xfanout206 _09385_/S vssd1 vssd1 vccd1 vccd1 _09396_/S sky130_fd_sc_hd__clkbuf_4
X_09801_ fanout52/X _08184_/B fanout32/X fanout50/X vssd1 vssd1 vccd1 vccd1 _09802_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout217 _11021_/S vssd1 vssd1 vccd1 vccd1 _11235_/S sky130_fd_sc_hd__buf_4
XFILLER_0_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09732_/Y sky130_fd_sc_hd__nand2_1
Xfanout239 _07009_/A vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__clkbuf_16
X_07993_ _07993_/A _07993_/B vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__nand2_2
X_06944_ reg1_val[31] _12335_/A vssd1 vssd1 vccd1 vccd1 _06944_/X sky130_fd_sc_hd__and2_1
XANTENNA__07318__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _09663_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__nand2_1
X_06875_ _06875_/A _09403_/S vssd1 vssd1 vccd1 vccd1 _08655_/A sky130_fd_sc_hd__nor2_2
X_09594_ _10286_/S _11446_/B _12394_/A1 _06793_/A _09593_/X vssd1 vssd1 vccd1 vccd1
+ _09594_/X sky130_fd_sc_hd__o221a_1
X_08614_ _08603_/Y _08612_/Y _08613_/Y _08595_/X vssd1 vssd1 vccd1 vccd1 _08616_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08279__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08548_/A sky130_fd_sc_hd__or2_1
XANTENNA__13162__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09491__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _08476_/A _08476_/B vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ _07427_/A _07427_/B vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _07358_/A _07358_/B vssd1 vssd1 vccd1 vccd1 _07359_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09595__B _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ fanout85/X fanout79/X fanout75/X _10466_/A vssd1 vssd1 vccd1 vccd1 _07290_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07396__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ _09029_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _09028_/X sky130_fd_sc_hd__and2_1
XANTENNA__11889__A1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__buf_1
X_12941_ _13206_/A _13207_/A _13206_/B vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ hold305/X hold35/X vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11510__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _11823_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__or2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__A _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ _11841_/B _11754_/B vssd1 vssd1 vccd1 vccd1 _11756_/C sky130_fd_sc_hd__or2_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11500_/Y _11591_/Y _11593_/B vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__o21a_1
X_10705_ _10706_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__and2_1
XANTENNA__07493__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10636_ _10636_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__and2_1
XANTENNA__11026__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06922__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _13364_/CLK _13355_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10567_ _12107_/B1 _10553_/X _10566_/X _10545_/X vssd1 vssd1 vccd1 vccd1 _10567_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10498_ _11359_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__xnor2_1
X_12306_ _08971_/B _06939_/X _12305_/X _11975_/A vssd1 vssd1 vccd1 vccd1 dest_val[28]
+ sky130_fd_sc_hd__o211a_4
X_13286_ _13287_/CLK _13286_/D vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11329__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ _12347_/B _12293_/B hold242/A vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09725__S _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__nand2_1
X_12099_ _12098_/A _12098_/B _11612_/A vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__a21o_1
X_11119_ _11014_/A _11012_/X _11030_/S vssd1 vssd1 vccd1 vccd1 _11120_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11275__B _11275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _07016_/A reg1_val[23] vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06591_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _06591_/X sky130_fd_sc_hd__o311a_4
XFILLER_0_47_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08330_ _08378_/A _08378_/B _08320_/A vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11280__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _08214_/X _08260_/Y _08213_/X vssd1 vssd1 vccd1 vccd1 _08261_/X sky130_fd_sc_hd__a21o_1
X_07212_ _07213_/A _07213_/B vssd1 vssd1 vccd1 vccd1 _07212_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ _10468_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11032__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _07129_/A _08476_/A _12415_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07153_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08433__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07074_ _07074_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _07074_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08984__A1 _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13157__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _07973_/A _07973_/B _07973_/C vssd1 vssd1 vccd1 vccd1 _07977_/B sky130_fd_sc_hd__o21ai_1
X_06927_ _06927_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__nand2_4
X_09715_ _09379_/X _09381_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _10735_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06858_ _06858_/A _06858_/B vssd1 vssd1 vccd1 vccd1 _06858_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12048__A1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ _06799_/A _06801_/B1 _12632_/B _06788_/X vssd1 vssd1 vccd1 vccd1 _10286_/S
+ sky130_fd_sc_hd__a31oi_4
X_09577_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__nand2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ _08459_/A _08459_/B _08459_/C vssd1 vssd1 vccd1 vccd1 _08680_/C sky130_fd_sc_hd__nand3_2
X_11470_ _11470_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06742__B _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _11021_/S _10421_/B vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _13140_/A _13140_/B vssd1 vssd1 vccd1 vccd1 _13141_/B sky130_fd_sc_hd__nand2_1
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08015__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ hold12/X _13071_/A2 _13071_/B1 hold43/A _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold13/A sky130_fd_sc_hd__o221a_1
XANTENNA__06986__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12280_/A _12019_/Y _12374_/D _09148_/Y vssd1 vssd1 vccd1 vccd1 _12022_/X
+ sky130_fd_sc_hd__o31a_1
X_10283_ _09716_/X _09718_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07573__B _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12287__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ hold275/X hold86/X vssd1 vssd1 vccd1 vccd1 _12925_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10837__A2 _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ hold98/X hold269/X vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _12615_/S _11806_/B _11891_/B vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__or3_2
X_12786_ hold3/X _12797_/B _12785_/Y _13109_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11737_ _11737_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10470__B1 _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ _11668_/A _11668_/B vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ _11169_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _11599_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11599_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10222__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ _13343_/CLK _13338_/D vssd1 vssd1 vccd1 vccd1 _13338_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07769__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _13375_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09915__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _10585_/B2 _10227_/B1 _10463_/A1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 _07831_/B
+ sky130_fd_sc_hd__o22a_1
X_07761_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07829_/A sky130_fd_sc_hd__xnor2_1
X_06712_ reg2_val[15] _06712_/B vssd1 vssd1 vccd1 vccd1 _06712_/X sky130_fd_sc_hd__and2_1
X_09500_ _09500_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12829__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07692_ _07692_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__xor2_1
X_06643_ reg2_val[31] _06712_/B vssd1 vssd1 vccd1 vccd1 _06643_/X sky130_fd_sc_hd__and2_1
XFILLER_0_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09197_/X _09250_/B _09722_/S vssd1 vssd1 vccd1 vccd1 _09431_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06574_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06922_/B sky130_fd_sc_hd__and4b_4
XANTENNA__13006__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09362_ _09135_/A _09135_/B _09133_/Y vssd1 vssd1 vccd1 vccd1 _09363_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ _08313_/A _08313_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07457__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__B1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _10234_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__B2 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_33 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 reg1_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08240_/A _08240_/B _08243_/Y vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08175_ _08556_/A _08175_/B vssd1 vssd1 vccd1 vccd1 _08178_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08406__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ reg1_val[27] _07126_/B vssd1 vssd1 vccd1 vccd1 _07126_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _07068_/B _07058_/C _07058_/A vssd1 vssd1 vccd1 vccd1 _07060_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__08709__A1 _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07674__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__A3 _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _07959_/A _07959_/B _07959_/C vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__or3_1
X_10970_ _10836_/A _10836_/B _10833_/A vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10819__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout51_A _07059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _07944_/B _07243_/X _07250_/X fanout28/X vssd1 vssd1 vccd1 vccd1 _09630_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07696__A1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__B2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11229__C1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__B _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ _12639_/A _12636_/Y _12638_/B vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_127_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _12616_/A _12572_/B vssd1 vssd1 vccd1 vccd1 _12573_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10452__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11522_/Y sky130_fd_sc_hd__xnor2_1
X_11453_ _11453_/A wire8/X vssd1 vssd1 vccd1 vccd1 _11453_/Y sky130_fd_sc_hd__nand2_1
X_10404_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__and2_1
X_11384_ fanout61/X fanout22/X fanout14/X _11645_/A vssd1 vssd1 vccd1 vccd1 _11385_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ hold303/X _12780_/B _13122_/X _12781_/A vssd1 vssd1 vccd1 vccd1 hold304/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09070__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ _10235_/B _10235_/C _10235_/A vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07620__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__B2 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ _11557_/A _13078_/B2 hold145/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__o21a_1
X_10266_ _10319_/B _10650_/A vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__nor2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12005_ _12083_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12007_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08176__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _11361_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10199_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11834__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ hold95/X hold308/A vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _12143_/A _12842_/A2 hold99/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold100/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06647__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__A2 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07439__A1 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ _12763_/A _12765_/B _12763_/B vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ _09847_/A _09847_/B _09845_/Y vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09185__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07494__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ _08931_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__nor2_1
X_08862_ _09668_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11171__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _07919_/A _07811_/Y _07809_/Y vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ _07934_/B _07996_/Y _07932_/X vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09667__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ _08354_/A2 _10227_/B1 _10463_/A1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 _07745_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07678__A1 _06973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B2 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _07736_/B vssd1 vssd1 vccd1 vccd1 _07675_/Y sky130_fd_sc_hd__inv_2
X_06626_ reg1_val[27] _07029_/A vssd1 vssd1 vccd1 vccd1 _06626_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ hold321/A _06942_/Y hold285/A vssd1 vssd1 vccd1 vccd1 _09414_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _11359_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _09277_/A _09277_/B _09277_/C vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ _08566_/A _08227_/B vssd1 vssd1 vccd1 vccd1 _08231_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12187__B1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _08104_/A _08104_/B _08102_/X vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09052__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07109_ _07109_/A _07109_/B _07109_/C _07109_/D vssd1 vssd1 vccd1 vccd1 _07116_/B
+ sky130_fd_sc_hd__or4_2
X_08089_ _08092_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08094_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10120_ _10121_/B _10121_/A vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ _11169_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07118__B1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10955_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07669__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10884_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12485__A _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__nand2_2
X_12554_ _12559_/B _12554_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12965__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _11320_/X _11506_/B _11503_/X vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12485_ _12652_/B _12485_/B vssd1 vssd1 vccd1 vccd1 _12486_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _06704_/B _11435_/X _12394_/A1 _06704_/A vssd1 vssd1 vccd1 vccd1 _11436_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11367_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09594__A1 _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13106_/Y sky130_fd_sc_hd__xnor2_1
X_10318_ _10133_/A _10317_/Y _10316_/Y vssd1 vssd1 vccd1 vccd1 _10318_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11298_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11300_/B sky130_fd_sc_hd__and2_1
X_13037_ hold191/A _13055_/A2 _13053_/B1 hold141/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold142/A sky130_fd_sc_hd__o221a_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12350__B1 _09239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _10110_/A _10110_/B _10094_/A vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09897__A2 _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__A _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07124__A3 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08321__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ _07460_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__xor2_1
X_07391_ _06973_/A fanout64/X fanout58/X _06973_/Y vssd1 vssd1 vccd1 vccd1 _07392_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08085__B2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A1 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _08937_/A _08937_/B _08940_/A vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_115_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09061_ _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _08008_/Y _08067_/A vssd1 vssd1 vccd1 vccd1 _08012_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07832__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout101_A _07068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__B2 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__A1 _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _10081_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07596__B1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__and2_1
XANTENNA__08113__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11144__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _09892_/Y _09894_/B vssd1 vssd1 vccd1 vccd1 _09895_/B sky130_fd_sc_hd__nand2b_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10789__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08184_/B _11083_/A _10966_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _08846_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11474__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _08776_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07727_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07733_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10655__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__xnor2_4
X_06609_ instruction[38] _06657_/B vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__and2_4
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07589_ _09671_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07600_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10407__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ _09329_/A _09329_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09328_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout14_A fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09259_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09259_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07823__B2 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07823__A1 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12270_ _12270_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12271_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _11413_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _12053_/A1 _11148_/X _11151_/X vssd1 vssd1 vccd1 vccd1 dest_val[14] sky130_fd_sc_hd__o21ai_4
XANTENNA__09119__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _07111_/Y _11296_/A _11188_/A fanout44/X vssd1 vssd1 vccd1 vccd1 _10104_/B
+ sky130_fd_sc_hd__o22a_2
X_11083_ _11083_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12332__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ curr_PC[4] _10035_/C curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08551__A2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _12257_/A fanout22/X fanout14/X _12202_/B vssd1 vssd1 vccd1 vccd1 _11986_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08839__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _11568_/A fanout42/X fanout40/X _07968_/B vssd1 vssd1 vccd1 vccd1 _10937_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09789__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _10867_/A _10867_/B vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__and2_1
XFILLER_0_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _12610_/A _12597_/B _12601_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _12607_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13104__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10949__B2 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10949__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10798_ hold305/A _11029_/A2 _10915_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09264__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ _12537_/A _12537_/B _12537_/C vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12468_ _12474_/B _12468_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XANTENNA__11559__A _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ _10537_/B _11004_/Y _11415_/Y _11418_/Y vssd1 vssd1 vccd1 vccd1 _11420_/B
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__12662__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _09243_/B _12386_/X _12398_/X vssd1 vssd1 vccd1 vccd1 _12399_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06960_ _11446_/A _07074_/A vssd1 vssd1 vccd1 vccd1 _06960_/X sky130_fd_sc_hd__and2_1
X_06891_ instruction[5] _06891_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xor2_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07772__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ _08630_/A _08630_/B _08638_/A vssd1 vssd1 vccd1 vccd1 _08666_/A sky130_fd_sc_hd__and3_1
XFILLER_0_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _08561_/A _08561_/B _08561_/C vssd1 vssd1 vccd1 vccd1 _08673_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07512_ _07705_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07718_/C sky130_fd_sc_hd__or2_1
X_08492_ _08493_/A _08493_/B vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__or2_1
XFILLER_0_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12837__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout17 _08985_/Y vssd1 vssd1 vccd1 vccd1 _12404_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout28 _07198_/X vssd1 vssd1 vccd1 vccd1 fanout28/X sky130_fd_sc_hd__clkbuf_8
X_07443_ _07446_/A _07446_/B vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06835__B _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout39 _07150_/Y vssd1 vssd1 vccd1 vccd1 _07539_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08108__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09113_ _11054_/A _09113_/B vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__xnor2_1
X_07374_ _07171_/X _07212_/X _07218_/Y _07182_/Y vssd1 vssd1 vccd1 vccd1 _07375_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ _09025_/A _09025_/B _09026_/Y vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11469__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11188__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ fanout55/X _10463_/B2 _10228_/A _12202_/A vssd1 vssd1 vccd1 vccd1 _09947_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__11117__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09182_/X _09206_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__mux2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _07605_/A _07605_/B _07608_/X vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08759_ _08759_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__nand2_1
X_11770_ _11593_/A _11682_/X _11684_/B vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09494__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A _10721_/B vssd1 vssd1 vccd1 vccd1 _10724_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_95_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13042__A1 _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ _09549_/B _10129_/C _10650_/X _10651_/Y _10649_/Y vssd1 vssd1 vccd1 vccd1
+ _10653_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_118_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10602_/A sky130_fd_sc_hd__nand2_1
X_13371_ _13374_/CLK hold194/X vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09797__A1 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _12320_/Y _12322_/B vssd1 vssd1 vccd1 vccd1 _12405_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12404_/B _12253_/B vssd1 vssd1 vccd1 vccd1 _12255_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11205_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12184_ _12164_/X _12165_/Y _12183_/X _12163_/X vssd1 vssd1 vccd1 vccd1 _12184_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08221__B2 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__A1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11135_ _11529_/B _11239_/B hold234/A vssd1 vssd1 vccd1 vccd1 _11135_/Y sky130_fd_sc_hd__a21oi_1
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__or2_1
XANTENNA__07592__A _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ hold261/A _10153_/C _10427_/A2 vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06936__A _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _07016_/A _11446_/B _11967_/X _06662_/B vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09312__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11899_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__and2b_1
X_10919_ _12395_/A1 _10918_/X _06732_/B vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09788__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09788__A1 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ _11125_/A _11231_/A _07121_/C _12717_/B _07229_/B vssd1 vssd1 vccd1 vccd1
+ _07190_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06671__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout229 _10158_/A2 vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__buf_4
Xfanout207 _08476_/A vssd1 vssd1 vccd1 vccd1 _09385_/S sky130_fd_sc_hd__buf_4
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__xnor2_1
Xfanout218 _07145_/A vssd1 vssd1 vccd1 vccd1 _11021_/S sky130_fd_sc_hd__buf_2
XFILLER_0_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07992_ _08000_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _07993_/B sky130_fd_sc_hd__nand2b_1
X_06943_ _12415_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _06943_/Y sky130_fd_sc_hd__nand2_2
X_09731_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09731_/X sky130_fd_sc_hd__or2_1
XANTENNA__09193__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06874_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__or2_4
X_09662_ _09662_/A _09662_/B vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__nand2_1
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__or2_1
X_08613_ _08595_/A _08595_/B _08602_/A _08595_/D vssd1 vssd1 vccd1 vccd1 _08613_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08279__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__and2_1
XANTENNA__11283__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _07424_/Y _07547_/B _07421_/X vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07357_ _07357_/A _07357_/B vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07288_ _11168_/A _07288_/B vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__xnor2_1
X_09027_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__buf_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A1 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _10326_/A _07581_/A _07581_/B _07218_/Y _07345_/X vssd1 vssd1 vccd1 vccd1
+ _09930_/B sky130_fd_sc_hd__a32o_1
XANTENNA__10849__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ hold71/X hold291/X vssd1 vssd1 vccd1 vccd1 _13206_/B sky130_fd_sc_hd__nand2b_1
X_12871_ hold277/X hold56/X vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__nand2b_1
X_11822_ _12065_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__xor2_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11753_ _11753_/A _11753_/B vssd1 vssd1 vccd1 vccd1 _11754_/B sky130_fd_sc_hd__and2_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11684_ _11684_/A _11684_/B vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__or2_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10933_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13015__B2 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07493__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ _10635_/A _10635_/B _10635_/C vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__or3_1
XFILLER_0_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13354_ _13364_/CLK _13354_/D vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _09148_/Y _12280_/X _12281_/Y _12304_/X vssd1 vssd1 vccd1 vccd1 _12305_/X
+ sky130_fd_sc_hd__a31o_1
X_10566_ _09222_/Y _10552_/X _10565_/Y _09155_/S _10563_/Y vssd1 vssd1 vccd1 vccd1
+ _10566_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10497_ _11749_/A fanout31/X fanout29/X _11734_/A vssd1 vssd1 vccd1 vccd1 _10498_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13285_ _13287_/CLK hold209/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11329__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ _13300_/Q _12236_/B vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11837__A _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__nor2_1
X_11118_ _11863_/A _08737_/Y _08739_/X _08740_/Y _11946_/A vssd1 vssd1 vccd1 vccd1
+ _11118_/X sky130_fd_sc_hd__a41o_1
X_12098_ _12098_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _12098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11049_ _11050_/B _11050_/A vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07181__A1 _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06590_/X sky130_fd_sc_hd__or4bb_1
XANTENNA__10188__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08130__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08260_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07211_ _07211_/A _11453_/A vssd1 vssd1 vccd1 vccd1 _07211_/X sky130_fd_sc_hd__or2_2
XFILLER_0_55_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _08553_/B1 _08400_/B fanout82/X _09468_/B2 vssd1 vssd1 vccd1 vccd1 _08192_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09188__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ _07142_/A _07142_/B vssd1 vssd1 vccd1 vccd1 _07356_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08433__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ _06963_/A _06963_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07944__B _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _08650_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _07975_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08121__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__or2_4
X_09714_ _10315_/A _09714_/B _09714_/C vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or3_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06857_ _12162_/A _06856_/X _06853_/X vssd1 vssd1 vccd1 vccd1 _06858_/B sky130_fd_sc_hd__a21o_1
X_09645_ fanout64/X _10463_/B2 _10228_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _09646_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__A1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06788_ reg2_val[2] _06794_/B vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__and2_1
X_09576_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09576_/Y sky130_fd_sc_hd__nor2_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__B2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08624_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08458_ _08459_/A _08459_/B _08459_/C vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__and3_1
XFILLER_0_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11008__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07409_ _07422_/B _07409_/B vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__and2b_1
X_10420_ _10420_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _10420_/Y sky130_fd_sc_hd__xnor2_1
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08423_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _10351_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__nor2_1
X_13070_ _12193_/A _13072_/A2 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__o21a_1
X_10282_ _10288_/S _10281_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10282_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06986__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11657__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ _12280_/A _12374_/D vssd1 vssd1 vccd1 vccd1 _12021_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12923_ _13170_/A _13171_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__10837__A3 _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ hold291/X hold71/X vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__nand2b_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ curr_PC[21] _11892_/C vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__and2_1
X_12785_ _12785_/A _12797_/B vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__nand2_1
X_11736_ _11736_/A _11736_/B vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__or2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12995__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06702__A_N _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _11668_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ _12202_/B fanout74/X _12257_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _10619_/B
+ sky130_fd_sc_hd__o22a_1
X_11598_ _11599_/B vssd1 vssd1 vccd1 vccd1 _11598_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13337_ _13343_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
X_10549_ _10547_/Y _10549_/B vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268_ _13375_/CLK hold100/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09915__A1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199_ hold314/A _13198_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__mux2_1
X_12219_ _11941_/B _12215_/Y _12218_/Y vssd1 vssd1 vccd1 vccd1 _12220_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__09915__B2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07760_/Y sky130_fd_sc_hd__nand2_1
X_06711_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07780__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ _09430_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _09430_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07691_ _07693_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _07691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06642_ _12043_/S _06642_/B vssd1 vssd1 vccd1 vccd1 _06655_/B sky130_fd_sc_hd__nand2_2
X_06573_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06573_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09361_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09363_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11789__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08654__A1 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ fanout64/X _10233_/B2 _10233_/A1 fanout58/X vssd1 vssd1 vccd1 vccd1 _09293_/B
+ sky130_fd_sc_hd__o22a_1
X_08312_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08313_/B sky130_fd_sc_hd__or2_1
XANTENNA__07457__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08302_/B _08302_/A vssd1 vssd1 vccd1 vccd1 _08243_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout229_A _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _07078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08174_ _08533_/B _08521_/A2 _08551_/A2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08175_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08406__A1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__B2 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ reg1_val[26] _07093_/A _07134_/B vssd1 vssd1 vccd1 vccd1 _07126_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07020__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07056_ _07067_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _07058_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10381__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11713__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A1 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _07955_/A _07955_/B _07955_/C vssd1 vssd1 vccd1 vccd1 _07959_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09381__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ instruction[11] _06913_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
X_07889_ _11168_/A _07889_/B vssd1 vssd1 vccd1 vccd1 _07953_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13218__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout44_A fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07696__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _09560_/B vssd1 vssd1 vccd1 vccd1 _09559_/Y sky130_fd_sc_hd__inv_2
X_12570_ reg1_val[20] curr_PC[20] _12615_/S vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12977__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10452__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11521_ _11433_/A _11430_/Y _11432_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06753__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11452_ _11809_/A _11809_/B _11809_/C _11808_/A vssd1 vssd1 vccd1 vccd1 _11542_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__08026__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ _11988_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__xnor2_1
X_10403_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__or2_1
XANTENNA__09070__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ hold283/X _13121_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__mux2_1
X_10334_ _10203_/A _10203_/B _10200_/A vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09070__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07620__A2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11704__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ _13324_/Q _13055_/A2 _13053_/B1 hold144/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold145/A sky130_fd_sc_hd__o221a_1
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10650_/B sky130_fd_sc_hd__xnor2_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12004_ _12004_/A _12004_/B vssd1 vssd1 vccd1 vccd1 _12005_/B sky130_fd_sc_hd__or2_1
X_10196_ fanout57/X fanout35/X fanout32/X _11837_/A vssd1 vssd1 vccd1 vccd1 _10197_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11468__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ _13125_/A _13126_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__a21bo_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ hold98/X _12839_/B vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__or2_1
XANTENNA__07105__A _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12665__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ _12766_/X _12768_/B vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__07439__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ curr_PC[19] _11718_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11720_/C sky130_fd_sc_hd__a21oi_1
X_12699_ _12699_/A _12699_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08930_ _08931_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__and2_1
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ fanout67/X _08633_/B _09300_/A fanout64/X vssd1 vssd1 vccd1 vccd1 _08862_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11171__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10903__C1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07919_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06583__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ _08792_/A _08792_/B vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ _08573_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout179_A _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _07910_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07736_/B sky130_fd_sc_hd__xnor2_4
X_06625_ reg2_val[27] _06712_/B _06600_/Y _06624_/Y vssd1 vssd1 vccd1 vccd1 _07029_/A
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07015__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ _09222_/Y _09412_/X _09408_/A vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__o21a_1
XANTENNA__12959__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ _10222_/A2 fanout28/X _07255_/Y _07944_/B vssd1 vssd1 vccd1 vccd1 _09345_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10376__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11631__B1 _11606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09275_ _09507_/B _09275_/B vssd1 vssd1 vccd1 vccd1 _09277_/C sky130_fd_sc_hd__or2_1
XFILLER_0_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08226_ _06875_/A fanout79/X fanout75/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08227_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08157_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07108_ _07109_/C _07109_/D vssd1 vssd1 vccd1 vccd1 _07108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09052__B2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__A1 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08088_ _08320_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ _07039_/A _07039_/B vssd1 vssd1 vccd1 vccd1 _07082_/B sky130_fd_sc_hd__xor2_2
X_10050_ _11980_/A fanout77/X fanout73/X fanout57/X vssd1 vssd1 vccd1 vccd1 _10051_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07118__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _11054_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10954_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07669__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10673__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ reg1_val[1] _12622_/B vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _12610_/A _12547_/B _12559_/A vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11504_ _11504_/A _11595_/A vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12484_ _12652_/B _12485_/B vssd1 vssd1 vccd1 vccd1 _12495_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _06704_/A _09228_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__or2_1
XFILLER_0_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ _11296_/A _11296_/B _11296_/C vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ _13105_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__nand2_1
X_10317_ _10650_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _10317_/Y sky130_fd_sc_hd__nor2_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10248_ _10248_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__xnor2_4
X_13036_ _07280_/B _13052_/A2 hold192/X vssd1 vssd1 vccd1 vccd1 _13316_/D sky130_fd_sc_hd__a21boi_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11153__A2 _11258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__A3 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _10045_/A _10044_/B _10042_/X vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06658__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13063__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07390_ _10937_/A _07396_/B vssd1 vssd1 vccd1 vccd1 _07413_/A sky130_fd_sc_hd__and2_1
XANTENNA__12810__C1 _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _09061_/B _09061_/A vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__nand2b_1
X_08011_ _08049_/B _08011_/B _08011_/C vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07832__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09196__S _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ fanout60/X _08184_/B fanout32/X fanout52/X vssd1 vssd1 vccd1 vccd1 _09963_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07596__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07596__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__A2 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08913_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09893_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__nand2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _09787_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08848_/A sky130_fd_sc_hd__xnor2_1
X_08775_ _08161_/Y _08214_/X _08160_/Y vssd1 vssd1 vccd1 vccd1 _08787_/A sky130_fd_sc_hd__a21o_1
X_07726_ _07723_/B _07803_/B _07723_/A vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10655__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__xor2_4
X_06608_ _06656_/A vssd1 vssd1 vccd1 vccd1 _06608_/Y sky130_fd_sc_hd__inv_2
X_07588_ fanout67/X _09297_/A1 fanout55/X _09297_/B2 vssd1 vssd1 vccd1 vccd1 _07589_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _09329_/A _09329_/B _09329_/C vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09258_/X sky130_fd_sc_hd__or2_1
XANTENNA__07823__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12525__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ reg1_val[4] reg1_val[27] _09560_/A vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__mux2_1
X_08209_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__xnor2_2
X_11220_ _10772_/B _11219_/Y _11599_/A vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _12525_/S _11255_/B _11151_/C vssd1 vssd1 vccd1 vccd1 _11151_/X sky130_fd_sc_hd__or3_2
XANTENNA__10591__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__nor2_2
X_11082_ _12131_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__xnor2_1
X_10033_ _10001_/X _10002_/Y _10003_/Y _10004_/X _10032_/X vssd1 vssd1 vccd1 vccd1
+ _10033_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_98_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _12004_/A sky130_fd_sc_hd__and2_1
XANTENNA__08839__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ _10935_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10939_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10867_/B sky130_fd_sc_hd__or2_1
XFILLER_0_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12399__A1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09264__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10949__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797_ _11029_/A2 _10915_/B hold305/A vssd1 vssd1 vccd1 vccd1 _10797_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13060__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07275__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09264__B2 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12536_ _12537_/A _12537_/B _12537_/C vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ _12467_/A _12467_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _11002_/X _11415_/A _11769_/B vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12398_ _12392_/Y _12393_/X _12397_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _12398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ hold326/A _12178_/A2 _11528_/C _12433_/A1 vssd1 vssd1 vccd1 vccd1 _11349_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06890_ instruction[3] _06873_/X _06884_/X _06888_/Y _06886_/X vssd1 vssd1 vccd1
+ vccd1 _06891_/B sky130_fd_sc_hd__a221o_2
X_13019_ hold83/X _13055_/A2 _13053_/B1 hold18/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold161/A sky130_fd_sc_hd__o221a_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08884__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ _08561_/A _08561_/B _08561_/C vssd1 vssd1 vccd1 vccd1 _08672_/A sky130_fd_sc_hd__and3_1
XFILLER_0_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07705_/B sky130_fd_sc_hd__xnor2_1
X_08491_ _08491_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08493_/B sky130_fd_sc_hd__xnor2_1
Xfanout18 _08985_/Y vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout29 _07198_/X vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__clkbuf_8
X_07442_ _09668_/A _07442_/B vssd1 vssd1 vccd1 vccd1 _07446_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07373_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09112_ _08096_/B _11083_/A _10966_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _09113_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09030_/A _09030_/B _09028_/X vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10573__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09945_ _10613_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07963__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ _09167_/X _09175_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__mux2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08827_/A _08827_/B vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08758_ _08758_/A _08758_/B _08758_/C vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__nand3_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09494__A1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ _07146_/Y _07944_/B fanout28/X _07153_/Y vssd1 vssd1 vccd1 vccd1 _07710_/B
+ sky130_fd_sc_hd__a22o_1
X_08689_ _07997_/A _07997_/B _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08689_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10721_/A _10721_/B vssd1 vssd1 vccd1 vccd1 _10720_/X sky130_fd_sc_hd__and2_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13042__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10133_/A _10133_/B _10650_/X vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ _10581_/B _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _13374_/CLK hold151/X vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09797__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ _12320_/A _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ fanout12/X fanout9/X fanout4/X _12309_/A vssd1 vssd1 vccd1 vccd1 _12253_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _11204_/B vssd1 vssd1 vccd1 vccd1 _11203_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12183_ _12182_/X _12183_/B _12183_/C _12183_/D vssd1 vssd1 vccd1 vccd1 _12183_/X
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08221__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ hold259/A _11134_/B vssd1 vssd1 vccd1 vccd1 _11239_/B sky130_fd_sc_hd__or2_1
X_11065_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12305__A1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__B _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _10013_/X _10015_/X _10288_/S vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11966_/A _12431_/A2 _11966_/Y _09225_/X vssd1 vssd1 vccd1 vccd1 _11967_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10918_ _09886_/B _12394_/A1 _10918_/S vssd1 vssd1 vccd1 vccd1 _10918_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _12068_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _11083_/A fanout9/X fanout4/X _10966_/A vssd1 vssd1 vccd1 vccd1 _10850_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12954__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12241__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09788__A2 _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ _12679_/B _12520_/B vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12792__A1 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12673__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06671__B _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout208 _06801_/X vssd1 vssd1 vccd1 vccd1 _08476_/A sky130_fd_sc_hd__clkbuf_8
X_07991_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__xnor2_1
X_06942_ _12378_/S _12417_/A vssd1 vssd1 vccd1 vccd1 _06942_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__10413__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09730_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07971__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ instruction[6] _06872_/Y _06864_/X vssd1 vssd1 vccd1 vccd1 _06873_/X sky130_fd_sc_hd__a21bo_1
X_09661_ _09662_/A _09662_/B vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__or2_1
X_09592_ hold322/A _10158_/A2 _09590_/X _09240_/X vssd1 vssd1 vccd1 vccd1 _09593_/B
+ sky130_fd_sc_hd__a31o_1
X_08612_ _08622_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _08612_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__A2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08673_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11283__A1 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_A _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06846__B _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout161_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__B2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B2 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08474_ _08475_/B _08475_/A vssd1 vssd1 vccd1 vccd1 _08474_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13024__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11035__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07356_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07357_/B sky130_fd_sc_hd__or2_1
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07287_ _08354_/A2 fanout73/X fanout71/X fanout77/X vssd1 vssd1 vccd1 vccd1 _07288_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06998__C1 _06964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _09027_/B _09027_/A vssd1 vssd1 vccd1 vccd1 _09026_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__buf_1
X_09928_ _09928_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07962__A1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__B2 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__B2 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _09042_/A _09042_/B _09858_/X vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__a21o_1
X_12870_ hold319/A hold53/X vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__nand2b_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ fanout37/X _07593_/Y _08857_/Y _07151_/A vssd1 vssd1 vccd1 vccd1 _11822_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11753_/A _11753_/B vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__nor2_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _11683_/A _11683_/B _11683_/C vssd1 vssd1 vccd1 vccd1 _11684_/B sky130_fd_sc_hd__and3_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _11568_/A _07151_/A _07155_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _10704_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13015__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10634_ _10635_/A _10635_/B _10635_/C vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13353_ _13363_/CLK _13353_/D vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ _12304_/A _12304_/B _12304_/C _12304_/D vssd1 vssd1 vccd1 vccd1 _12304_/X
+ sky130_fd_sc_hd__or4_1
X_10565_ _10565_/A vssd1 vssd1 vccd1 vccd1 _10565_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10496_ _10933_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13284_ _13287_/CLK _13284_/D vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12235_ _09875_/Y _12234_/Y _12421_/B vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11837__B _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12106_/A _12103_/Y _12105_/B vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__o21a_1
X_11117_ _11863_/A _08737_/Y _08739_/X _08740_/Y vssd1 vssd1 vccd1 vccd1 _11117_/Y
+ sky130_fd_sc_hd__a22oi_2
X_12097_ _06865_/X _12096_/X _12378_/S vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09155__A0 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06947__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ hold204/X _13143_/B2 _13209_/A2 hold228/A vssd1 vssd1 vccd1 vccd1 hold205/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10469__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08130__A1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07469__B1 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08130__B2 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07210_ _07210_/A _07210_/B vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__and2_1
X_08190_ _08320_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08969__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ _10937_/A _07141_/B vssd1 vssd1 vccd1 vccd1 _07142_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08433__A2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ _10339_/A _07072_/B vssd1 vssd1 vccd1 vccd1 _07072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07974_ _08649_/B fanout98/X fanout83/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _07975_/B
+ sky130_fd_sc_hd__o22a_1
X_06925_ instruction[6] instruction[5] _09235_/A vssd1 vssd1 vccd1 vccd1 _06925_/X
+ sky130_fd_sc_hd__or3_4
X_09713_ _10315_/A _09714_/B _09714_/C vssd1 vssd1 vccd1 vccd1 _09713_/Y sky130_fd_sc_hd__o21ai_1
X_06856_ _12098_/A _06855_/X _06854_/X vssd1 vssd1 vccd1 vccd1 _06856_/X sky130_fd_sc_hd__a21o_1
X_09644_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10700__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _09219_/A curr_PC[0] _09411_/B _09409_/X vssd1 vssd1 vccd1 vccd1 _09579_/A
+ sky130_fd_sc_hd__a31oi_2
X_06787_ _06787_/A _06787_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__nor2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ _08641_/A2 _08553_/A2 _08551_/B1 _08649_/B vssd1 vssd1 vccd1 vccd1 _08527_/B
+ sky130_fd_sc_hd__o22a_1
X_08457_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08459_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_108_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07408_ _09766_/A _07408_/B vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_92_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _08420_/A _08420_/B _08352_/X vssd1 vssd1 vccd1 vccd1 _08423_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07339_ _07637_/B _07339_/B vssd1 vssd1 vccd1 vccd1 _07341_/B sky130_fd_sc_hd__and2_1
X_10350_ _10351_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _11021_/S _09199_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06986__A2 _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _09008_/A _08878_/B _09008_/Y vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__a21oi_2
X_12020_ _12020_/A _12020_/B _12020_/C _12020_/D vssd1 vssd1 vccd1 vccd1 _12374_/D
+ sky130_fd_sc_hd__and4_2
XANTENNA__11148__A2_N _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ hold59/X hold295/X vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06767__A _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ hold114/X hold301/X vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__and2b_1
X_12784_ _11917_/C _13072_/A2 hold10/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold11/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ curr_PC[21] _11892_/C vssd1 vssd1 vccd1 vccd1 _11806_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08112__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11735_ _11736_/A _11736_/B vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__nand2_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11666_ _11668_/B vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__inv_2
XFILLER_0_52_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10621_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11597_ _11597_/A _11768_/A vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__and2_1
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ _13344_/CLK _13336_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13267_ _13375_/CLK hold122/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10479_ _12131_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10488_/A sky130_fd_sc_hd__xnor2_1
X_12218_ _12089_/Y _12215_/B _12217_/A vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11707__C1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _13198_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13198_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11722__A2 _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08222__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ _12149_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12151_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06710_ _06711_/B vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06677__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07690_ _07690_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07693_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09053__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06641_ reg1_val[24] _06641_/B vssd1 vssd1 vccd1 vccd1 _06642_/B sky130_fd_sc_hd__or2_1
X_06572_ pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06893_/C sky130_fd_sc_hd__and2_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12435__B1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _09360_/A _09360_/B vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__xor2_1
X_08311_ _08682_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _08311_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_13 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08556_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08302_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_24 reg2_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _10161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__A _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_46 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12738__B2 _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08406__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08173_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__xor2_2
X_07124_ _11125_/A _11231_/A _07121_/C _07123_/X _07093_/A vssd1 vssd1 vccd1 vccd1
+ _07134_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_43_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ _06963_/A _06963_/B _06960_/X _07074_/B vssd1 vssd1 vccd1 vccd1 _07068_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__07090__A1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13163__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07957_ _07957_/A _07957_/B vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__or2_1
XANTENNA__07393__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__A1 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _06908_/A _06908_/B _06908_/C vssd1 vssd1 vccd1 vccd1 _06913_/B sky130_fd_sc_hd__or3_2
XANTENNA__11477__B2 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07888_ _08553_/A2 fanout73/X _08551_/B1 fanout77/X vssd1 vssd1 vccd1 vccd1 _07889_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13218__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06839_ reg1_val[19] _07058_/A vssd1 vssd1 vccd1 vccd1 _06839_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09627_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__and2_1
X_09558_ _10288_/S _09557_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__nor2_1
X_11520_ _11520_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09489_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09490_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10452__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__or2_1
XFILLER_0_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11382_ fanout51/X fanout9/X fanout4/X _11456_/A vssd1 vssd1 vccd1 vccd1 _11383_/B
+ sky130_fd_sc_hd__o22a_1
X_10402_ _10402_/A _10402_/B vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _13121_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13121_/Y sky130_fd_sc_hd__xnor2_1
X_10333_ _10458_/B _10333_/B vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__and2_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09070__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _07210_/B _13052_/A2 hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__a21boi_1
X_10264_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10264_/X sky130_fd_sc_hd__and2_1
X_12003_ _12004_/A _12004_/B vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__nand2_1
X_10195_ _10468_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08977__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__A _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12114__C1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13094__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11468__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ hold32/X hold303/X vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ _06978_/X _12842_/A2 hold121/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold122/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06944__B _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ reg1_val[30] _12767_/B vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__or2_1
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11640__A1 _11559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ curr_PC[19] curr_PC[20] _11718_/C vssd1 vssd1 vccd1 vccd1 _11892_/C sky130_fd_sc_hd__and3_1
XFILLER_0_44_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ _12698_/A _12698_/B _12698_/C vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__and3_2
XFILLER_0_25_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11661_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07121__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06960__A _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13319_ _13324_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11156__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _09669_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08572__A1 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__nor2_1
X_08791_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__or2_1
XANTENNA__12202__A _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07742_ _08594_/A2 fanout83/X fanout79/X _08572_/A2 vssd1 vssd1 vccd1 vccd1 _07743_/B
+ sky130_fd_sc_hd__o22a_2
X_07673_ _08533_/B fanout79/X fanout75/X _08507_/A2 vssd1 vssd1 vccd1 vccd1 _07674_/B
+ sky130_fd_sc_hd__o22a_2
X_06624_ _06706_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _06624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09412_ _11958_/A _09411_/Y _12107_/B1 vssd1 vssd1 vccd1 vccd1 _09412_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13081__B1 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11631__B2 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _09273_/B _09274_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07835__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09588__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08156_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07107_ _07093_/A _07092_/B _07190_/B reg1_val[22] vssd1 vssd1 vccd1 vccd1 _07109_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09052__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ _08553_/B1 _08274_/B fanout74/X _09468_/B2 vssd1 vssd1 vccd1 vccd1 _08088_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _07039_/A _07039_/B vssd1 vssd1 vccd1 vccd1 _07348_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12344__C1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _09324_/A fanout9/A fanout5/X _12785_/A vssd1 vssd1 vccd1 vccd1 _08990_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07118__A2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _12202_/B fanout27/X fanout25/X _12202_/A vssd1 vssd1 vccd1 vccd1 _10952_/B
+ sky130_fd_sc_hd__o22a_1
X_10882_ _10882_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10885_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12621_ _12621_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__or2_1
XFILLER_0_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _12610_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12559_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08037__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12782__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11503_ _11317_/Y _11410_/Y _11412_/B vssd1 vssd1 vccd1 vccd1 _11503_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ reg1_val[7] curr_PC[7] _12525_/S vssd1 vssd1 vccd1 vccd1 _12485_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11434_ _11143_/Y _11433_/Y _12171_/A vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07876__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__A1 _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__xor2_1
X_11296_ _11296_/A _11296_/B _11296_/C vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__or3_1
XFILLER_0_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11138__B1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13104_ _13109_/A hold294/X vssd1 vssd1 vccd1 vccd1 _13343_/D sky130_fd_sc_hd__and2_1
X_10316_ _10125_/X _10263_/X _10264_/X vssd1 vssd1 vccd1 vccd1 _10316_/Y sky130_fd_sc_hd__a21oi_1
X_10247_ _10247_/A _10247_/B vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__nor2_2
X_13035_ hold167/X _13055_/A2 _13053_/B1 hold191/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold192/A sky130_fd_sc_hd__o221a_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10361__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__B2 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _10066_/A _10066_/B _10057_/Y vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07116__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ hold50/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__or2_1
XANTENNA__11072__S _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__B _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ _08049_/A _07977_/B _07975_/Y vssd1 vssd1 vccd1 vccd1 _08011_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13118__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ _09770_/Y _09773_/B _09769_/A vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07596__A2 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__xor2_4
X_09892_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09892_/Y sky130_fd_sc_hd__nor2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout191_A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _09659_/B2 fanout85/X _10466_/A fanout98/X vssd1 vssd1 vccd1 vccd1 _08844_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10151__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _08769_/A _08769_/B _08773_/A _08773_/B _11692_/B vssd1 vssd1 vccd1 vccd1
+ _11863_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__A _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07725_ _07725_/A _07725_/B vssd1 vssd1 vccd1 vccd1 _07803_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10655__A2 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07656_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07656_/X sky130_fd_sc_hd__and2_1
XANTENNA__06584__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ _06605_/X _06607_/B vssd1 vssd1 vccd1 vccd1 _06656_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_48_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07587_ _07587_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _11155_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09329_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ curr_PC[0] _12525_/S _09256_/X vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ _08268_/A _08268_/B _08204_/X vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ reg1_val[5] reg1_val[26] _09560_/A vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _08198_/A _08137_/Y _08127_/X vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__a21o_1
X_11150_ curr_PC[13] _11149_/C curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11151_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10591__A1 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11946__A _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _11456_/A fanout22/X fanout14/X _11386_/A vssd1 vssd1 vccd1 vccd1 _11082_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10850__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11540__B1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _09226_/Y _10008_/Y _12171_/B _09180_/S _10031_/X vssd1 vssd1 vccd1 vccd1
+ _10032_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08320__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__A2 _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13363_/CLK sky130_fd_sc_hd__clkbuf_8
X_11983_ _11983_/A _11983_/B _11983_/C vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__or3_1
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08839__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ _10935_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _11045_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12610_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_94_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12535_ _12544_/A _12535_/B vssd1 vssd1 vccd1 vccd1 _12537_/C sky130_fd_sc_hd__nand2_1
X_10796_ hold308/A _10796_/B vssd1 vssd1 vccd1 vccd1 _10915_/B sky130_fd_sc_hd__or2_1
XANTENNA__09264__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12466_ _12467_/A _12467_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_30_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11417_ _11216_/X _11597_/A _11416_/X vssd1 vssd1 vccd1 vccd1 _11769_/B sky130_fd_sc_hd__a21o_1
X_12397_ _09196_/S _09408_/Y _09434_/Y _09223_/Y _12396_/Y vssd1 vssd1 vccd1 vccd1
+ _12397_/X sky130_fd_sc_hd__o221a_2
XFILLER_0_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11348_ _11529_/B _11528_/C hold326/A vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11279_ _11397_/B _11279_/B vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__or2_1
XANTENNA__11531__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _08648_/A _13078_/B2 hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__o21a_1
XANTENNA__09326__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__A _11593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10098__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _10231_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__xnor2_1
X_08490_ _08490_/A _08490_/B vssd1 vssd1 vccd1 vccd1 _08493_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout19 _11155_/A vssd1 vssd1 vccd1 vccd1 _11296_/B sky130_fd_sc_hd__buf_6
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _08633_/B fanout60/X fanout52/X _09300_/A vssd1 vssd1 vccd1 vccd1 _07442_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07372_ _07372_/A _07372_/B vssd1 vssd1 vccd1 vccd1 _07373_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09111_ _08935_/A _08935_/B _08932_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__a21o_1
X_09042_ _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08405__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout204_A _06901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10022__B1 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10573__B2 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__A1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _12059_/A fanout85/X _10466_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _09945_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _11237_/S _09874_/Y _09252_/A vssd1 vssd1 vccd1 vccd1 _09875_/Y sky130_fd_sc_hd__a21oi_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08825_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08827_/B sky130_fd_sc_hd__and2b_1
X_08757_ _08758_/B _08758_/C _08758_/A vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__a21o_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09494__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ _09795_/A _07708_/B vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__xnor2_4
X_08688_ _08266_/X _08761_/B _08681_/X _08687_/X _08261_/X vssd1 vssd1 vccd1 vccd1
+ _08772_/B sky130_fd_sc_hd__o221a_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _07640_/A _07640_/B vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ _10650_/A _10650_/B _10650_/C _10767_/A vssd1 vssd1 vccd1 vccd1 _10650_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12786__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ fanout60/X fanout85/X _10466_/A fanout52/X vssd1 vssd1 vccd1 vccd1 _09310_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11053__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _10582_/B _10581_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12250__B2 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10680__A2_N _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ _12320_/A _12320_/B _12320_/C vssd1 vssd1 vccd1 vccd1 _12320_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _12404_/B _12204_/A _12203_/B _12202_/X vssd1 vssd1 vccd1 vccd1 _12263_/A
+ sky130_fd_sc_hd__o31a_1
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__xnor2_2
X_12182_ _09222_/Y _12171_/B _10016_/X _09155_/S _12181_/Y vssd1 vssd1 vccd1 vccd1
+ _12182_/X sky130_fd_sc_hd__a221o_1
XANTENNA__06768__B1 _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11958_/A _11132_/Y _11129_/Y _09243_/B vssd1 vssd1 vccd1 vccd1 _11133_/X
+ sky130_fd_sc_hd__a211o_1
X_11064_ _12068_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06783__A3 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _09556_/Y _10014_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _11966_/A _11966_/B vssd1 vssd1 vccd1 vccd1 _11966_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ hold330/A _11029_/A2 _11027_/B _10916_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _10921_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11897_ fanout40/X _07301_/Y _07593_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _11898_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10848_ _12131_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10852_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10779_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09788__A3 _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ reg1_val[12] curr_PC[12] _12525_/S vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12792__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ _12627_/B _12450_/B vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__B1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10555__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10490__A _10490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout209 _12785_/A vssd1 vssd1 vccd1 vccd1 _09403_/S sky130_fd_sc_hd__buf_6
X_07990_ _07990_/A _08154_/A vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__nor2_1
X_06941_ instruction[6] instruction[5] _06940_/B vssd1 vssd1 vccd1 vccd1 _06941_/X
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _11361_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09662_/B sky130_fd_sc_hd__xnor2_1
X_06872_ _06943_/B _06871_/X _06863_/X vssd1 vssd1 vccd1 vccd1 _06872_/Y sky130_fd_sc_hd__o21ai_1
X_08611_ _08611_/A _08611_/B vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__xor2_1
X_09591_ _10158_/A2 _09590_/X hold322/A vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11807__A1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _08542_/A _08542_/B _08542_/C vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__nor3_1
XANTENNA__11283__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__A2 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _08504_/A _08504_/B _08468_/X vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout154_A _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _07547_/A vssd1 vssd1 vccd1 vccd1 _07424_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07355_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08436__B1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07286_ _10230_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10794__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _09025_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _09927_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07962__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _09858_/A _09996_/A _10128_/A _10267_/A vssd1 vssd1 vccd1 vccd1 _09858_/X
+ sky130_fd_sc_hd__or4_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11510__A3 _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ _10234_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09791_/B sky130_fd_sc_hd__xnor2_1
X_08809_ _08809_/A _08809_/B _08809_/C vssd1 vssd1 vccd1 vccd1 _09038_/B sky130_fd_sc_hd__or3_1
X_11820_ _11820_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11829_/A sky130_fd_sc_hd__xnor2_1
X_11751_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__xnor2_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _10702_/A _10702_/B vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__xor2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11682_ _11683_/A _11683_/B _11683_/C vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__a21o_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__B1 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10633_ _10633_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _10635_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11026__A2 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _13352_/CLK _13352_/D vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__dfxtp_1
X_10564_ _11131_/A _10151_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ _12294_/Y _12295_/X _12302_/X vssd1 vssd1 vccd1 vccd1 _12304_/D sky130_fd_sc_hd__o21ai_1
X_10495_ _07077_/X _07151_/A _07155_/A _07237_/Y vssd1 vssd1 vccd1 vccd1 _10496_/B
+ sky130_fd_sc_hd__a22o_1
X_13283_ _13287_/CLK hold215/X vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ _10315_/A _08800_/A _08800_/B _12029_/A vssd1 vssd1 vccd1 vccd1 _12165_/Y
+ sky130_fd_sc_hd__o31ai_2
X_11116_ _11115_/A _11259_/A _11258_/A vssd1 vssd1 vccd1 vccd1 _11116_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06756__A3 _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12096_ _06655_/B _12024_/Y _12043_/S vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__o21a_1
X_11047_ _11045_/A _11045_/B _11048_/B vssd1 vssd1 vccd1 vccd1 _11197_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12998_ _13144_/A hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__and2_1
XANTENNA__07469__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _11947_/A _11865_/X _11883_/S vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08130__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07469__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08969__B2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _07128_/Y _07402_/B fanout41/X _08476_/A vssd1 vssd1 vccd1 vccd1 _07141_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__B1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ _09938_/A _07071_/B vssd1 vssd1 vccd1 vccd1 _07072_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__S _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _09603_/Y _09710_/Y _09711_/Y vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__o21a_1
X_07973_ _07973_/A _07973_/B _07973_/C vssd1 vssd1 vccd1 vccd1 _08049_/A sky130_fd_sc_hd__or3_2
X_06924_ instruction[6] instruction[5] _09235_/A vssd1 vssd1 vccd1 vccd1 _06924_/Y
+ sky130_fd_sc_hd__nor3_2
XANTENNA__10700__A1 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06855_ reg1_val[24] _06975_/A vssd1 vssd1 vccd1 vccd1 _06855_/X sky130_fd_sc_hd__and2_1
X_09643_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10700__B2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _09567_/X _09573_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06786_ reg1_val[3] _07145_/A vssd1 vssd1 vccd1 vccd1 _06787_/B sky130_fd_sc_hd__and2_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08525_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11008__A2 _11041_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _08420_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07407_ _07539_/B _07153_/Y fanout37/X _07128_/Y vssd1 vssd1 vccd1 vccd1 _07408_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07338_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07339_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ _07197_/Y fanout24/X _09114_/B1 _08096_/B vssd1 vssd1 vccd1 vccd1 _07270_/B
+ sky130_fd_sc_hd__o22a_1
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__nand2_1
X_09008_ _09008_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _09008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11716__B1 _11693_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _13165_/B _13166_/A _12865_/X vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09143__B _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ hold307/A hold129/X vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12783_ hold9/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__or2_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _06964_/B _11446_/B _06941_/X _11802_/X vssd1 vssd1 vccd1 vccd1 _11803_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12785__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ _11734_/A _11917_/C _11734_/C vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__and3_1
XFILLER_0_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _11569_/A _11569_/B _11567_/A vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__o21a_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10616_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11596_ _11416_/X _11768_/A _11594_/X vssd1 vssd1 vccd1 vccd1 _11596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13335_ _13344_/CLK _13335_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10547_/Y sky130_fd_sc_hd__nor2_1
X_13266_ _13372_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__dfxtp_1
X_10478_ _10966_/A fanout22/X fanout14/X _10859_/A vssd1 vssd1 vccd1 vccd1 _10479_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12217_ _12217_/A vssd1 vssd1 vccd1 vccd1 _12217_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08179__A2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _13197_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06729__A3 _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _12149_/B _12149_/A vssd1 vssd1 vccd1 vccd1 _12212_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11722__A3 _11809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__B2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _12080_/A _12080_/B _12080_/C vssd1 vssd1 vccd1 vccd1 _12151_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06958__A _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12679__B _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__B _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ reg1_val[24] _06641_/B vssd1 vssd1 vccd1 vccd1 _12043_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ instruction[0] pred_val vssd1 vssd1 vccd1 vccd1 _06893_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12435__A1 _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09290_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__nor2_1
X_08310_ _08682_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _08310_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_14 reg2_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ _08533_/B _08551_/A2 _08551_/B1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08242_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07311__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_25 reg2_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_36 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_47 reg1_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__B _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08172_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08172_/X sky130_fd_sc_hd__and2_1
XFILLER_0_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _07123_/A _07342_/C vssd1 vssd1 vccd1 vccd1 _07123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07090__A2 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ _10231_/A _10061_/A _07053_/X vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__o21a_2
XANTENNA__09509__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__A2 _06901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11174__A1 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B2 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07029__A _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07956_ _07911_/B _07956_/B vssd1 vssd1 vccd1 vccd1 _07957_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09244__A _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ instruction[13] _06907_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
XANTENNA__11477__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ _09787_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__xnor2_2
X_06838_ _06877_/B _11513_/B _06837_/X vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__a21o_1
X_09626_ _09827_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06769_ reg2_val[5] _06794_/B _12421_/B vssd1 vssd1 vccd1 vccd1 _06952_/C sky130_fd_sc_hd__a21o_2
X_09557_ _11021_/S _09556_/Y _09251_/B vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12977__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09490_/A sky130_fd_sc_hd__or2_1
XANTENNA__10437__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07699__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ _08556_/A _08508_/B vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08439_ _08463_/A _08463_/B _08435_/X vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_108_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _12053_/A1 _11445_/Y _11446_/Y _11449_/Y vssd1 vssd1 vccd1 vccd1 dest_val[17]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11381_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10401_ _10401_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_33_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__nand2_1
X_10332_ _10332_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ hold26/X _13055_/A2 _13053_/B1 _13324_/Q _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold27/A sky130_fd_sc_hd__o221a_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _12080_/B _12002_/B vssd1 vssd1 vccd1 vccd1 _12004_/B sky130_fd_sc_hd__and2_1
X_10263_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__or2_1
X_10194_ _12202_/B _08400_/B fanout82/X _12202_/A vssd1 vssd1 vccd1 vccd1 _10195_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12499__B _12499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11468__A2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _13120_/A _13121_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08993__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ hold120/X _12839_/B vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__or2_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10428__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08097__A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__B2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12766_ reg1_val[30] _12773_/A vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__and2_1
XANTENNA__08097__B2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__A2 _07193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _06996_/A _11446_/B _06941_/X _11716_/X vssd1 vssd1 vccd1 vccd1 _11717_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10466__C _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _12698_/A _12698_/B _12698_/C vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07121__B _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06960__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13318_ _13324_/CLK _13318_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08233__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__A1 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__B2 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13249_ _13346_/CLK hold31/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
X_08790_ _08790_/A _08790_/B vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08572__A2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _07810_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07283__S _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _07850_/A _07850_/B _07737_/Y vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__12202__B _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07532__B1 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06623_ instruction[37] _06657_/B vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__and2_4
X_09411_ _09411_/A _09411_/B vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12959__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13081__A1 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _09274_/B _09273_/B vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07835__B2 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__A1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ _08320_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__xnor2_1
X_07106_ _07087_/X _12717_/B _07092_/B _07229_/B reg1_val[22] vssd1 vssd1 vccd1 vccd1
+ _07109_/C sky130_fd_sc_hd__o311a_1
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ _08445_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11147__A1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ _07037_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _07039_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08988_ _08874_/A _11645_/B _12360_/B vssd1 vssd1 vccd1 vccd1 _08988_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__07771__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _07939_/X sky130_fd_sc_hd__or2_1
X_10950_ _11052_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__xnor2_1
X_10881_ _10882_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__nand2_1
X_09609_ _09612_/A vssd1 vssd1 vccd1 vccd1 _09609_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10848__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ _12624_/A _12620_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__and2_4
XFILLER_0_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ reg1_val[17] curr_PC[17] _12615_/S vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__mux2_2
X_11502_ _11500_/Y _11502_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__nand2b_4
X_12482_ _12488_/B _12482_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
XFILLER_0_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11433_ _11433_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11364_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11296_/C sky130_fd_sc_hd__xnor2_1
X_13103_ hold293/X _13222_/A2 _13102_/X _13108_/B2 vssd1 vssd1 vccd1 vccd1 hold294/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13274__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ _10315_/A _10315_/B vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__or2_1
X_10246_ _10245_/B _10245_/C _10245_/A vssd1 vssd1 vccd1 vccd1 _10247_/B sky130_fd_sc_hd__a21oi_1
X_13034_ _10469_/A _13052_/A2 hold168/X vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09200__A0 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__A1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _10119_/A _10119_/B _10120_/X vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__07762__B1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13134__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06955__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ _07237_/Y _12842_/A2 hold75/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold76/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12810__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12749_ _12757_/A _12749_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06971__A _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__B2 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A1 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _10113_/B _09960_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__or2_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08911_ _08912_/B _08912_/A vssd1 vssd1 vccd1 vccd1 _08911_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09891_ _09729_/X _09730_/Y _09732_/Y vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__o21a_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08842_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__xnor2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _11777_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07026__B _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ _07542_/B _07542_/C _07542_/D _07543_/A vssd1 vssd1 vccd1 vccd1 _07725_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07657_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06606_ reg1_val[29] _08971_/A vssd1 vssd1 vccd1 vccd1 _06607_/B sky130_fd_sc_hd__or2_1
XANTENNA__10655__A3 _10810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13054__A1 _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07586_ _07586_/A _07586_/B _07586_/C vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_48_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _09675_/A fanout9/A fanout5/X _09467_/A vssd1 vssd1 vccd1 vccd1 _09326_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _06940_/Y _09255_/X _12053_/A1 vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13297__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09187_ _09185_/X _09186_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08138_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08070_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _11296_/B _11080_/B vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10591__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10031_ _09882_/X _10016_/X _10018_/Y _09237_/Y _10030_/X vssd1 vssd1 vccd1 vccd1
+ _10031_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13219__A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ _11983_/A _11983_/B _11983_/C vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__o21ai_1
X_10933_ _10933_/A _10933_/B vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _10864_/A _10864_/B vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10295__A2_N _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12616_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__and2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10795_ _12395_/A1 _10794_/X _06738_/B vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ _12691_/B _12534_/B vssd1 vssd1 vccd1 vccd1 _12535_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07887__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ _12474_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12467_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11416_ _11213_/Y _11317_/Y _11319_/B vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__o21a_1
X_12396_ _12396_/A _12396_/B vssd1 vssd1 vccd1 vccd1 _12396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11347_ hold210/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11528_/C sky130_fd_sc_hd__or2_1
XANTENNA__10031__B2 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__and2_1
XANTENNA__13129__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _10230_/B _10230_/C _10736_/A vssd1 vssd1 vccd1 vccd1 _10231_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08868__D _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ hold147/A _13055_/A2 _13053_/B1 hold83/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold84/A sky130_fd_sc_hd__o221a_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07127__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06966__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__A1 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06685__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__B2 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ _10234_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07446_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12244__C1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ _07369_/A _07369_/B _07454_/A vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09110_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09041_ _09544_/A _08917_/X _09706_/A _09547_/B _09547_/A vssd1 vssd1 vccd1 vccd1
+ _09042_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09412__B1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10022__A1 _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__A1 _11593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07974__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap197 _06924_/Y vssd1 vssd1 vccd1 vccd1 _12107_/B1 sky130_fd_sc_hd__buf_4
X_09943_ _09943_/A _09943_/B vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09874_ _11021_/S _09723_/X _09251_/B vssd1 vssd1 vccd1 vccd1 _09874_/Y sky130_fd_sc_hd__o21ai_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08826_/B _08825_/B vssd1 vssd1 vccd1 vccd1 _08827_/A sky130_fd_sc_hd__and2b_1
XANTENNA__06876__A _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ _08748_/B _08748_/C _08748_/A _08687_/D vssd1 vssd1 vccd1 vccd1 _08758_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11286__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _09928_/A _08096_/B fanout24/X _09815_/A vssd1 vssd1 vccd1 vccd1 _07708_/B
+ sky130_fd_sc_hd__o22a_2
X_08687_ _08776_/B _08687_/B _08758_/A _08687_/D vssd1 vssd1 vccd1 vccd1 _08687_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _08902_/A _07638_/B vssd1 vssd1 vccd1 vccd1 _07640_/B sky130_fd_sc_hd__nor2_1
X_07569_ _07569_/A _07569_/B vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__xor2_1
X_09308_ _09471_/B _09308_/B vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ _12068_/A _10580_/B vssd1 vssd1 vccd1 vccd1 _10581_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ _09240_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09239_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _12223_/X _12227_/X _12249_/X _12189_/X _11975_/A vssd1 vssd1 vccd1 vccd1
+ dest_val[27] sky130_fd_sc_hd__o32a_4
XFILLER_0_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11201_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__and2_1
X_12181_ _07026_/B _11446_/B _12180_/X vssd1 vssd1 vccd1 vccd1 _12181_/Y sky130_fd_sc_hd__o21ai_1
X_11132_ _11237_/S _09433_/X _11131_/X vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11063_ _11734_/A fanout42/X fanout41/X _11568_/A vssd1 vssd1 vccd1 vccd1 _11064_/B
+ sky130_fd_sc_hd__a22o_1
X_10014_ _09395_/X _09404_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _10014_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11692__A _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ hold289/A _12175_/A2 _12040_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11965_/X
+ sky130_fd_sc_hd__a31o_1
X_10916_ _11029_/A2 _11027_/B hold330/A vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__a21oi_1
X_11896_ _11843_/A _11843_/B _11842_/A vssd1 vssd1 vccd1 vccd1 _11930_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09890__B1 _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ _11296_/A _07347_/B fanout15/X _11188_/A vssd1 vssd1 vccd1 vccd1 _10848_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10778_ _06822_/X _10777_/X _12025_/S vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08506__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12517_ _12523_/B _12517_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
XFILLER_0_82_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ reg1_val[2] curr_PC[2] _12525_/S vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12379_ _12381_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__or2_1
XANTENNA__12462__S _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10490__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06940_ _09396_/S _06940_/B vssd1 vssd1 vccd1 vccd1 _06940_/Y sky130_fd_sc_hd__nand2_1
X_06871_ _12381_/A _06870_/X _06849_/Y vssd1 vssd1 vccd1 vccd1 _06871_/X sky130_fd_sc_hd__a21bo_1
X_08610_ _08610_/A _08610_/B _08610_/C vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__and3_2
X_09590_ hold265/A _13338_/Q vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__or2_1
X_08541_ _08514_/B _08514_/C _08514_/A vssd1 vssd1 vccd1 vccd1 _08675_/B sky130_fd_sc_hd__a21oi_2
X_08472_ _08472_/A _08472_/B vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07423_ _07423_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07547_/A sky130_fd_sc_hd__or2_2
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A _07048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07354_ _07352_/Y _07354_/B vssd1 vssd1 vccd1 vccd1 _07355_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08436__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08987__A2 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ fanout98/X _10463_/B2 _10228_/A fanout83/X vssd1 vssd1 vccd1 vccd1 _07286_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06998__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _08905_/A _08905_/B _08903_/Y vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold331/X vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__buf_1
X_09926_ _09924_/X _09926_/B vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__nand2b_1
X_09857_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__xnor2_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _10233_/B2 _10466_/B _10466_/C _10233_/A1 fanout55/X vssd1 vssd1 vccd1 vccd1
+ _09789_/B sky130_fd_sc_hd__o32a_1
X_08808_ _08808_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _08808_/Y sky130_fd_sc_hd__nand2_1
X_08739_ _08746_/B _08746_/D _08746_/C vssd1 vssd1 vccd1 vccd1 _08739_/X sky130_fd_sc_hd__a21o_1
X_11750_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__nor2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _12068_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10702_/B sky130_fd_sc_hd__xor2_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09872__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ _11683_/A _11683_/B _11683_/C vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__a21oi_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ _10624_/B _10489_/B _10506_/B _10505_/B _10505_/A vssd1 vssd1 vccd1 vccd1
+ _10633_/B sky130_fd_sc_hd__a32o_1
X_13351_ _13352_/CLK _13351_/D vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _10555_/Y _10556_/X _10562_/X vssd1 vssd1 vccd1 vccd1 _10563_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _12297_/Y _12298_/X _12301_/X vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ _10494_/A _10494_/B vssd1 vssd1 vccd1 vccd1 _10505_/A sky130_fd_sc_hd__xor2_2
X_13282_ _13287_/CLK _13282_/D vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ _12231_/Y _12233_/B vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _10315_/A _08800_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__o21a_1
X_12095_ _12278_/B _12094_/B _09149_/X vssd1 vssd1 vccd1 vccd1 _12095_/X sky130_fd_sc_hd__a21o_1
X_11115_ _11115_/A _11259_/A _11258_/A vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__and3_1
X_11046_ _09787_/A _10942_/B _10945_/X vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap112_A _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ hold199/X _13204_/B2 _13186_/A2 hold204/A vssd1 vssd1 vccd1 vccd1 hold200/A
+ sky130_fd_sc_hd__a22o_1
X_11948_ reg1_val[22] _06994_/A _12025_/S vssd1 vssd1 vccd1 vccd1 _11948_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07469__A2 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ hold316/A _11879_/A2 _11963_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11879_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09091__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _09938_/A _07071_/B vssd1 vssd1 vccd1 vccd1 _10339_/A sky130_fd_sc_hd__or2_1
XANTENNA__09091__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10006__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _09603_/Y _09710_/Y _11889_/A1 vssd1 vssd1 vccd1 vccd1 _09711_/Y sky130_fd_sc_hd__a21oi_1
X_07972_ _09941_/A _07972_/B vssd1 vssd1 vccd1 vccd1 _07973_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06923_ instruction[22] _06575_/X _06922_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08354__B1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ reg1_val[25] _06978_/A vssd1 vssd1 vccd1 vccd1 _06854_/X sky130_fd_sc_hd__and2_1
XANTENNA__10161__B1 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10700__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06785_ reg1_val[3] _07145_/A vssd1 vssd1 vccd1 vccd1 _06785_/X sky130_fd_sc_hd__or2_1
X_09573_ _09569_/X _09572_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12989__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _09941_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _08528_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08455_ _08455_/A _08455_/B vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08386_ _08394_/A _08394_/B _08372_/X vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__a21o_1
X_07406_ _07410_/A _07406_/B vssd1 vssd1 vccd1 vccd1 _07422_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10216__A1 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__B2 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07358_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07199_ _06811_/B _11237_/S _06950_/X _06949_/Y vssd1 vssd1 vccd1 vccd1 _07264_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ _09064_/C _09007_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_103_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11716__B2 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _12193_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09705__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _13160_/A _13161_/A _13160_/B vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12131__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__nor2_1
X_11802_ _11774_/Y _11775_/X _11777_/Y _11778_/X _11801_/X vssd1 vssd1 vccd1 vccd1
+ _11802_/X sky130_fd_sc_hd__o221a_1
X_12782_ _12782_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _12782_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ _11733_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__xor2_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10586__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11664_ _11557_/A _11557_/B _11562_/A vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__o21ai_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10615_ _11361_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10617_/B sky130_fd_sc_hd__xnor2_1
X_11595_ _11595_/A _11686_/A vssd1 vssd1 vccd1 vccd1 _11768_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_52_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ _13334_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ _10420_/A _10417_/Y _10419_/B vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_12_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13372_/CLK hold103/X vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
X_10477_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10507_/B sky130_fd_sc_hd__and2_1
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12216_ _12082_/Y _12324_/B _12324_/C vssd1 vssd1 vccd1 vccd1 _12217_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ _13226_/A hold315/X vssd1 vssd1 vccd1 vccd1 _13362_/D sky130_fd_sc_hd__and2_1
XANTENNA__10930__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _12212_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__or2_1
X_12078_ _12151_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12080_/C sky130_fd_sc_hd__nand2_1
X_11029_ hold319/A _11029_/A2 _11243_/C _11028_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _11033_/B sky130_fd_sc_hd__a311o_1
XANTENNA__06958__B _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ rst vssd1 vssd1 vccd1 vccd1 _13219_/A sky130_fd_sc_hd__inv_2
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12435__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07311__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__B2 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 reg2_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08171_ _08171_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08173_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07122_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07342_/C sky130_fd_sc_hd__or2_2
XFILLER_0_15_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07090__A3 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ _09668_/A _07053_/B _09938_/A vssd1 vssd1 vccd1 vccd1 _07053_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_113_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07029__B _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _07955_/A _07955_/B _07955_/C vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__and3_1
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ instruction[12] _06907_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
X_09625_ fanout45/X _10859_/A fanout71/X _07814_/B vssd1 vssd1 vccd1 vccd1 _09626_/B
+ sky130_fd_sc_hd__o22a_1
X_07886_ _08521_/A2 fanout85/X _10466_/A _07201_/X vssd1 vssd1 vccd1 vccd1 _07887_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11882__B1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ reg1_val[18] _07067_/A vssd1 vssd1 vccd1 vccd1 _06837_/X sky130_fd_sc_hd__and2_1
XANTENNA__10685__B2 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ reg2_val[5] _06794_/B _12421_/B vssd1 vssd1 vccd1 vccd1 _06811_/B sky130_fd_sc_hd__a21oi_4
X_09556_ _09556_/A vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__inv_2
X_06699_ instruction[27] _06699_/B vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__and2_4
XANTENNA__12097__S _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _11361_/A _09487_/B vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__xnor2_1
X_08507_ _09403_/S _08507_/A2 _08619_/B1 _08533_/B vssd1 vssd1 vccd1 vccd1 _08508_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ _08438_/A _08438_/B vssd1 vssd1 vccd1 vccd1 _08463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08369_/Y sky130_fd_sc_hd__nor2_1
X_11380_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__and2_1
XFILLER_0_61_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10332_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__or2_1
XANTENNA__09419__B _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _10262_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__xnor2_4
X_13050_ _11172_/A _13078_/B2 hold107/X vssd1 vssd1 vccd1 vccd1 _13323_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _12001_/A _12001_/B _12001_/C vssd1 vssd1 vccd1 vccd1 _12002_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12362__A1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06577__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _10105_/A _10105_/B _10102_/A vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06778__B _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__B1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ hold38/X hold283/X vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10676__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _07012_/Y _12842_/A2 hold109/X _13134_/A vssd1 vssd1 vccd1 vccd1 hold110/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/A _12765_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
XANTENNA__08097__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11716_ _11690_/Y _11691_/X _11693_/Y _11946_/A _11715_/X vssd1 vssd1 vccd1 vccd1
+ _11716_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__B _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__A3 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ reg1_val[15] _12696_/B vssd1 vssd1 vccd1 vccd1 _12698_/C sky130_fd_sc_hd__xnor2_2
X_11647_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__or2_1
XANTENNA__07121__C _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09046__A1 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09046__B2 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11578_ _11579_/B _11579_/A vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07057__B1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09597__A2 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10529_ _10529_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__xnor2_4
X_13317_ _13324_/CLK hold143/X vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11156__A2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ _13343_/CLK _13248_/D vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _13179_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11875__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__or2_1
XANTENNA__12202__C _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07671_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07671_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07532__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06622_ _12415_/B _06622_/B vssd1 vssd1 vccd1 vccd1 _12381_/A sky130_fd_sc_hd__or2_2
X_09410_ _12621_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09411_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07532__B2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__and2_1
XANTENNA__11115__A _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07296__B1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _10937_/A _09272_/B vssd1 vssd1 vccd1 vccd1 _09273_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07835__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ _08619_/B1 _08274_/B fanout74/X _09403_/S vssd1 vssd1 vccd1 vccd1 _08224_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08154_ _08154_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07105_ _11559_/A vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ _08521_/A2 _10227_/B1 _10463_/A1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 _08086_/B
+ sky130_fd_sc_hd__o22a_1
X_07036_ _07037_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _07348_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12344__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08987_ _08874_/A _11645_/B _12360_/B vssd1 vssd1 vccd1 vccd1 fanout5/A sky130_fd_sc_hd__o21a_1
XANTENNA__07771__B2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _07938_/X sky130_fd_sc_hd__and2_1
XANTENNA__11855__B1 _11853_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07869_ _07869_/A _07869_/B _07869_/C vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__and3_1
X_10880_ _10880_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10882_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _09930_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout42_A _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09539_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13072__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12559_/A _12550_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07287__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ _11501_/A _11501_/B _11501_/C vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_109_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12482_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11432_ _11430_/Y _11432_/B vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _11557_/A _11363_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__xnor2_1
X_13102_ hold317/A _13101_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11294_ _11988_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__xnor2_2
X_10314_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10346__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ _10245_/A _10245_/B _10245_/C vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__and3_1
X_13033_ hold178/A _13055_/A2 _13053_/B1 hold167/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold168/A sky130_fd_sc_hd__o221a_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10176_ _10124_/A _10124_/B _10122_/X vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07762__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12099__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _07043_/Y vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__buf_4
X_12817_ hold74/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__or2_1
XFILLER_0_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12810__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12767_/B _07342_/C _12757_/B vssd1 vssd1 vccd1 vccd1 _12749_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ reg1_val[12] _12679_/B vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10585__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09890_ _09888_/Y _09889_/X _07097_/C _06940_/B vssd1 vssd1 vccd1 vccd1 _09890_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08910_ _08910_/A _08910_/B vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08842_/B vssd1 vssd1 vccd1 vccd1 _08841_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09075__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08776_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07723_ _07723_/A _07723_/B vssd1 vssd1 vccd1 vccd1 _07803_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout177_A _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07654_ _07655_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07654_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ reg1_val[29] _08971_/A vssd1 vssd1 vccd1 vccd1 _06605_/X sky130_fd_sc_hd__and2_1
XANTENNA__07323__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13054__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07585_ _07586_/A _07586_/B _07586_/C vssd1 vssd1 vccd1 vccd1 _07587_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09324_ _09324_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07269__B1 _09114_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ _09150_/X _09151_/X _09254_/X _06941_/X vssd1 vssd1 vccd1 vccd1 _09255_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ _08206_/A _08206_/B vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09186_ reg1_val[6] reg1_val[25] _09560_/A vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08137_ _08138_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08137_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07441__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08067_/A _08067_/B _08067_/C vssd1 vssd1 vccd1 vccd1 _08070_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__A1 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ _09297_/B2 fanout58/X fanout56/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _07020_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12404__A wire8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _12171_/A _06924_/Y _10029_/Y _10024_/Y vssd1 vssd1 vccd1 vccd1 _10030_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07744__B2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _12056_/B _11981_/B vssd1 vssd1 vccd1 vccd1 _11983_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _11749_/A _07151_/A _07155_/A _11734_/A vssd1 vssd1 vccd1 vccd1 _10933_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10859__A _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10863_ _10863_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ reg1_val[25] curr_PC[25] _12615_/S vssd1 vssd1 vccd1 vccd1 _12604_/B sky130_fd_sc_hd__mux2_1
X_10794_ _09886_/B _12394_/A1 _10794_/S vssd1 vssd1 vccd1 vccd1 _10794_/X sky130_fd_sc_hd__mux2_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10594__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ _12691_/B _12534_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10803__A1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12793__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06791__B _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12464_ _12637_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07680__B1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ _11415_/A vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__inv_2
X_12395_ _12395_/A1 _12394_/X _06622_/B vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11346_ _06711_/B _11344_/X _11345_/X _11343_/X vssd1 vssd1 vccd1 vccd1 _11346_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11277_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__nor2_1
X_13016_ _13016_/A hold148/X vssd1 vssd1 vccd1 vccd1 _13306_/D sky130_fd_sc_hd__and2_1
XANTENNA__07408__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10228_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _10230_/C sky130_fd_sc_hd__or3_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07127__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06966__B _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12984__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06982__A _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ _09033_/A _09033_/B _08913_/X vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09412__A1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09942_ _09943_/A _09943_/B vssd1 vssd1 vccd1 vccd1 _09942_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07974__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _09886_/A _09871_/X _09872_/Y vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__o21a_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08824_/A _08824_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__xnor2_1
X_08755_ _08348_/Y _08391_/X _08685_/B vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11286__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _07712_/A _07712_/B vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__and2_1
XANTENNA__11286__B2 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07053__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ _08751_/A _08751_/B _08758_/A _08687_/D vssd1 vssd1 vccd1 vccd1 _08761_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07637_ _07637_/A _07637_/B _07637_/C vssd1 vssd1 vccd1 vccd1 _07638_/B sky130_fd_sc_hd__and3_1
XFILLER_0_76_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07568_ _09795_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _07569_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _09306_/B _09306_/C _09306_/A vssd1 vssd1 vccd1 vccd1 _09308_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07499_ _10468_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ _09240_/B _09238_/B vssd1 vssd1 vccd1 vccd1 _09238_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ reg1_val[8] reg1_val[23] _09180_/S vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11200_ _11200_/A vssd1 vssd1 vccd1 vccd1 _11202_/B sky130_fd_sc_hd__inv_2
X_12180_ _09225_/X _12179_/X _06654_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11062_ _12065_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10013_ _10011_/X _10012_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10589__A _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__B _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _12175_/A2 _12040_/B hold289/A vssd1 vssd1 vccd1 vccd1 _11964_/Y sky130_fd_sc_hd__a21oi_1
X_10915_ hold305/A _10915_/B vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__or2_1
X_11895_ _12020_/A _12020_/B _12020_/C _12280_/A vssd1 vssd1 vccd1 vccd1 _11895_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13018__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10846_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12226__B1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12309__A _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10660_/A _10658_/Y _10675_/S vssd1 vssd1 vccd1 vccd1 _10777_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12516_ _12516_/A _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06952__D _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _12453_/B _12447_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XFILLER_0_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12378_ _06870_/X _12381_/B _12378_/S vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08522__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11863_/A _08750_/A _08750_/B _11946_/A vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06870_ _06608_/Y _12335_/B _06850_/X vssd1 vssd1 vccd1 vccd1 _06870_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06696__B _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _08542_/B _08542_/C _08542_/A vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_106_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13009__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ _08471_/A vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__inv_2
XFILLER_0_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07892__B1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _07409_/B _07422_/B vssd1 vssd1 vccd1 vccd1 _07423_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07354_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08436__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07284_ _07281_/A _07281_/B _10230_/A vssd1 vssd1 vccd1 vccd1 _07284_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10962__A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ _09023_/A _09023_/B vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08432__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _09925_/A _09925_/B _09809_/X vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__or3b_1
X_09856_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _09856_/X sky130_fd_sc_hd__and2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _08809_/B _08809_/C vssd1 vssd1 vccd1 vccd1 _08808_/B sky130_fd_sc_hd__nor2_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09787_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__xnor2_1
X_06999_ _07000_/A _07000_/B vssd1 vssd1 vccd1 vccd1 _06999_/X sky130_fd_sc_hd__and2_2
XANTENNA__10202__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _08734_/A _08734_/B _08484_/X _08675_/B vssd1 vssd1 vccd1 vccd1 _08746_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08720_/B sky130_fd_sc_hd__xor2_2
X_10700_ _07077_/X fanout42/X fanout41/X _07237_/Y vssd1 vssd1 vccd1 vccd1 _10701_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11764_/B _11680_/B vssd1 vssd1 vccd1 vccd1 _11683_/C sky130_fd_sc_hd__nand2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__A2 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ _10477_/A _10477_/B _10474_/Y vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__o21ai_2
X_13350_ _13350_/CLK _13350_/D vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__dfxtp_1
X_10562_ _06747_/Y _10557_/Y _10559_/Y _10560_/X _10561_/X vssd1 vssd1 vccd1 vccd1
+ _10562_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _09155_/S _09728_/X _12291_/B _09222_/Y _12300_/X vssd1 vssd1 vccd1 vccd1
+ _12301_/X sky130_fd_sc_hd__a221o_1
X_13281_ _13287_/CLK _13281_/D vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__or2_1
X_12232_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12163_ _12162_/A _12162_/B _12162_/Y _11612_/A vssd1 vssd1 vccd1 vccd1 _12163_/X
+ sky130_fd_sc_hd__a211o_1
X_12094_ _12278_/B _12094_/B vssd1 vssd1 vccd1 vccd1 _12094_/Y sky130_fd_sc_hd__nor2_1
X_11114_ _11321_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__xnor2_4
X_11045_ _11045_/A _11045_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A2 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10170__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12996_ _13144_/A hold219/X vssd1 vssd1 vccd1 vccd1 _13296_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__or2_1
X_11878_ _11879_/A2 _11963_/B hold316/A vssd1 vssd1 vccd1 vccd1 _11878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08517__A _08517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ _11837_/A fanout46/X fanout44/X fanout61/X vssd1 vssd1 vccd1 vccd1 _10830_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09091__A2 _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07971_ _08619_/B2 fanout79/X fanout75/X _08619_/A2 vssd1 vssd1 vccd1 vccd1 _07972_/B
+ sky130_fd_sc_hd__o22a_1
X_06922_ instruction[29] _06922_/B vssd1 vssd1 vccd1 vccd1 _06922_/X sky130_fd_sc_hd__or2_1
X_09710_ _10267_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09710_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__09551__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ reg1_val[26] _07026_/B vssd1 vssd1 vccd1 vccd1 _06853_/X sky130_fd_sc_hd__and2_1
X_09641_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__nand2_1
X_06784_ reg1_val[3] _07145_/A vssd1 vssd1 vccd1 vccd1 _06787_/A sky130_fd_sc_hd__nor2_1
X_09572_ _09570_/X _09571_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09303__B1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ _08619_/B2 _08553_/B1 _09468_/B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08524_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10957__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout257_A _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08455_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08394_/B sky130_fd_sc_hd__xnor2_2
X_07405_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07406_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _09766_/A _07336_/B vssd1 vssd1 vccd1 vccd1 _07338_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07267_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07273_/B sky130_fd_sc_hd__and2_1
X_09006_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07198_ _07193_/B _07193_/A _11559_/A vssd1 vssd1 vccd1 vccd1 _07198_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09908_ fanout42/X _10712_/A _07212_/X fanout40/X vssd1 vssd1 vccd1 vccd1 _09909_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13227__B _13227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _09837_/Y _09839_/B vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__and2b_1
X_12850_ hold287/A hold68/X vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12429__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11801_ _11612_/A _11782_/Y _11789_/X _11800_/X vssd1 vssd1 vccd1 vccd1 _11801_/X
+ sky130_fd_sc_hd__o211a_1
X_12781_ _12781_/A _12781_/B vssd1 vssd1 vccd1 vccd1 _12839_/B sky130_fd_sc_hd__nor2_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__nand2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10614_ _12202_/A fanout35/X fanout33/X fanout64/X vssd1 vssd1 vccd1 vccd1 _10615_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _11410_/Y _11500_/Y _11502_/B vssd1 vssd1 vccd1 vccd1 _11594_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ _13344_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10545_ _06878_/A _10543_/X _10544_/Y vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__o21a_1
X_13264_ _13363_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
X_10476_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13195_ hold314/X _13209_/A2 _13194_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold315/A
+ sky130_fd_sc_hd__a22o_1
X_12215_ _12215_/A _12215_/B vssd1 vssd1 vccd1 vccd1 _12215_/Y sky130_fd_sc_hd__nand2_1
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12147_/B sky130_fd_sc_hd__and2_1
XFILLER_0_20_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ _12077_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__or2_1
X_11028_ _11029_/A2 _11243_/C hold319/A vssd1 vssd1 vccd1 vccd1 _11028_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12979_ hold259/A _13143_/B2 _13186_/A2 hold234/X vssd1 vssd1 vccd1 vccd1 hold235/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08639__A2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07151__A _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__A2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 reg2_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08170_/A _08170_/B vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_82_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07075__A1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _11125_/A _11231_/A _07121_/C _07123_/A vssd1 vssd1 vccd1 vccd1 _08868_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA__06990__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_49 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13148__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ _07891_/B _07891_/C vssd1 vssd1 vccd1 vccd1 _07052_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__07090__A4 _12717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__C1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__A _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07954_ _07954_/A _07954_/B vssd1 vssd1 vccd1 vccd1 _07955_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06905_ instruction[11] _06907_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
X_07885_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07885_/Y sky130_fd_sc_hd__nor2_1
X_06836_ _11428_/A _06834_/X _06835_/X vssd1 vssd1 vccd1 vccd1 _11513_/B sky130_fd_sc_hd__a21o_1
X_09624_ _11054_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09541__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ _06767_/A _06767_/B _12647_/B vssd1 vssd1 vccd1 vccd1 _06767_/X sky130_fd_sc_hd__or3b_2
XANTENNA__12378__S _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ _07152_/A _09397_/X _09249_/B vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06698_ _11531_/S _06698_/B vssd1 vssd1 vccd1 vccd1 _06877_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09486_ _09659_/B2 _08184_/B fanout32/X fanout98/X vssd1 vssd1 vccd1 vccd1 _09487_/B
+ sky130_fd_sc_hd__o22a_1
X_08506_ _08573_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08544_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _08573_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _08463_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08368_ _10468_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07319_ _10231_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _07321_/B sky130_fd_sc_hd__xnor2_2
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__and2_1
X_10330_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__xnor2_1
X_10261_ _10261_/A _10261_/B vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__xor2_4
X_12000_ _12001_/A _12001_/B _12001_/C vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12362__A2 _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _10192_/A _10192_/B vssd1 vssd1 vccd1 vccd1 _10248_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08620__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__B1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _13115_/A _13116_/A _13115_/B vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09451__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ hold108/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__or2_1
XANTENNA__13075__B1 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12764_ _12764_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__or2_2
X_11715_ _11715_/A _11715_/B _11715_/C _11715_/D vssd1 vssd1 vccd1 vccd1 _11715_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12695_ _12698_/B _12695_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
X_11646_ _11734_/C _11646_/B vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07121__D _07123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _11672_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ _10529_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__and2_1
X_13316_ _13324_/CLK _13316_/D vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13247_ _13343_/CLK _13247_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10459_ _10635_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__or2_1
XANTENNA__12353__A2 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _13187_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _13358_/D sky130_fd_sc_hd__and2_1
XANTENNA__09626__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12129_ _12058_/B _12060_/B _12058_/A vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06985__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _08573_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07532__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ reg1_val[30] _08971_/C vssd1 vssd1 vccd1 vccd1 _06622_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _11054_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ _07402_/B _09450_/B1 _07263_/Y fanout41/X vssd1 vssd1 vccd1 vccd1 _09272_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07296__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ _10468_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07296__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout122_A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ _07990_/A _07989_/B _07989_/C vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__o21a_1
X_07104_ _07109_/A _07109_/B vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__nor2_4
X_08084_ _08081_/Y _08140_/B _08080_/Y vssd1 vssd1 vccd1 vccd1 _08100_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ _09668_/A _07035_/B vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _12335_/A _08983_/B _11813_/A reg1_val[30] _12772_/A vssd1 vssd1 vccd1 vccd1
+ _12360_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07771__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _07937_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _07940_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07868_ _07921_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07869_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06819_ reg1_val[9] _07218_/A vssd1 vssd1 vccd1 vccd1 _06819_/X sky130_fd_sc_hd__and2_1
X_09607_ _07201_/X _07347_/B fanout15/X _07264_/X vssd1 vssd1 vccd1 vccd1 _09608_/B
+ sky130_fd_sc_hd__o22a_1
X_07799_ _07797_/A _07797_/B _07798_/Y vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__10210__A _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09538_/X sky130_fd_sc_hd__and2_1
XFILLER_0_109_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout35_A _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07287__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _11501_/A _11501_/B _11501_/C vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _11645_/B _09469_/B vssd1 vssd1 vccd1 vccd1 _09471_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07287__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1_A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10291__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11431_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11432_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09210__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ fanout25/X fanout11/X fanout7/A _07211_/X vssd1 vssd1 vccd1 vccd1 _11363_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _13101_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13101_/Y sky130_fd_sc_hd__xnor2_1
X_10313_ _10313_/A _10313_/B _10313_/C _10313_/D vssd1 vssd1 vccd1 vccd1 _10570_/B
+ sky130_fd_sc_hd__or4_1
X_11293_ _11456_/A fanout9/X fanout4/X _11386_/A vssd1 vssd1 vccd1 vccd1 _11294_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__A1 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10243_/B _10243_/C _10243_/A vssd1 vssd1 vccd1 vccd1 _10245_/C sky130_fd_sc_hd__o21ai_1
X_13032_ _07071_/B _12797_/B hold179/X vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09446__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10346__B2 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ _10137_/B _10137_/C _12420_/A vssd1 vssd1 vccd1 vccd1 _10175_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09880__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout180 _12847_/B vssd1 vssd1 vccd1 vccd1 _12797_/B sky130_fd_sc_hd__buf_4
Xfanout191 _08650_/A vssd1 vssd1 vccd1 vccd1 _08624_/A sky130_fd_sc_hd__buf_12
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _07243_/X _12842_/A2 hold81/X _13187_/A vssd1 vssd1 vccd1 vccd1 hold82/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12757_/B sky130_fd_sc_hd__or2_1
XFILLER_0_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10774__B _10810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ reg1_val[12] _12679_/B vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _11624_/Y _11625_/X _11628_/X vssd1 vssd1 vccd1 vccd1 _11630_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10585__A1 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__B2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06699__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _10234_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08776_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__or2_1
X_07722_ _07721_/A _07721_/C _07721_/B vssd1 vssd1 vccd1 vccd1 _07723_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07604__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06604_ _06602_/Y _06707_/B1 _06794_/B reg2_val[29] vssd1 vssd1 vccd1 vccd1 _08971_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12798__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09334_/A sky130_fd_sc_hd__xnor2_1
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07586_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08466__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__A1 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07269__B2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ instruction[5] _06864_/X _09240_/A _09221_/X _09253_/X vssd1 vssd1 vccd1
+ vccd1 _09254_/X sky130_fd_sc_hd__o311a_1
XANTENNA__10273__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09185_ reg1_val[7] reg1_val[24] _09560_/A vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__mux2_1
X_08205_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08206_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08136_ _08134_/A _08134_/B _08206_/A vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07441__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08067_/A _08067_/B _08067_/C vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__and3_1
XFILLER_0_31_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__A2 _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__A3 _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ _07010_/A _07010_/B _09671_/A vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__mux2_2
XANTENNA__12404__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _09297_/A1 _12257_/A fanout13/X _09297_/B2 vssd1 vssd1 vccd1 vccd1 _08970_/B
+ sky130_fd_sc_hd__o22a_2
X_11980_ _11980_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _11981_/B sky130_fd_sc_hd__nor2_1
X_10931_ _12131_/A _10931_/B vssd1 vssd1 vccd1 vccd1 _10935_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10859__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _10862_/A _10862_/B _10862_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__or3_1
XFILLER_0_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12601_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ hold207/A _11115_/A _10912_/B _10792_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _10800_/A sky130_fd_sc_hd__a311o_1
XFILLER_0_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _11125_/A curr_PC[14] _12615_/S vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__mux2_1
X_12463_ _12637_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07680__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _11414_/A _11597_/A vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__and2_1
XANTENNA__07680__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ _12431_/A2 _12394_/A1 _12415_/B vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10567__A1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__A2 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _06711_/A _11966_/B _11446_/B _07074_/A vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11276_ _11367_/A _11276_/B vssd1 vssd1 vccd1 vccd1 _11278_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ _07593_/A _07593_/B _10227_/B1 vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__a21o_1
X_13015_ hold147/X _13222_/A2 _13052_/A2 _09219_/A vssd1 vssd1 vccd1 vccd1 hold148/A
+ sky130_fd_sc_hd__a22o_1
X_10158_ hold309/A _10158_/A2 _10292_/B _09240_/X vssd1 vssd1 vccd1 vccd1 _10159_/B
+ sky130_fd_sc_hd__a31o_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__buf_1
XANTENNA__07127__C _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12244__A1 _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__S _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09948__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12505__A _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09943_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__06777__A3 _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07974__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09872_ _09886_/A _09871_/X _11612_/A vssd1 vssd1 vccd1 vccd1 _09872_/Y sky130_fd_sc_hd__a21oi_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A _08823_/B vssd1 vssd1 vccd1 vccd1 _08824_/B sky130_fd_sc_hd__xor2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _08749_/A _08749_/B _08753_/A _08753_/B _08750_/A vssd1 vssd1 vccd1 vccd1
+ _11511_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07705_ _07705_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07712_/B sky130_fd_sc_hd__xor2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11286__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08685_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08687_/D sky130_fd_sc_hd__or2_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07636_ _07637_/A _07637_/B _07637_/C vssd1 vssd1 vccd1 vccd1 _08902_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__12386__S _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ _10327_/B2 _08096_/B _10589_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _07568_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12786__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09306_/A _09306_/B _09306_/C vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__and3_1
XFILLER_0_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09240_/B _09238_/B vssd1 vssd1 vccd1 vccd1 _09237_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ _08354_/A2 _08400_/B fanout82/X _10585_/B2 vssd1 vssd1 vccd1 vccd1 _07499_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09939__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ _09160_/X _09167_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _08556_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08124_/A sky130_fd_sc_hd__xnor2_1
X_09099_ _09099_/A _09099_/B vssd1 vssd1 vccd1 vccd1 _09100_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12415__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ _10148_/X _10150_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__mux2_1
X_11061_ _06993_/Y _07151_/A _07155_/A _11749_/A vssd1 vssd1 vccd1 vccd1 _11062_/B
+ sky130_fd_sc_hd__a22o_1
X_10012_ _09390_/X _09401_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10589__B _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ hold316/A _11963_/B vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10914_ hold220/A _11115_/A _11024_/B _10913_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _10921_/A sky130_fd_sc_hd__a311o_1
X_11894_ _06908_/C _11890_/X _11893_/X vssd1 vssd1 vccd1 vccd1 dest_val[22] sky130_fd_sc_hd__o21ai_4
X_10845_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10776_ _10776_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12515_ _12516_/A _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12377_ _06607_/B _12334_/X _06605_/X vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11328_ _11863_/A _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _11328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11259_ _11259_/A _11809_/C vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12701__A2 _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06993__A _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _08573_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07892__A1 _07060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07421_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ _07282_/A _07282_/B _10230_/A vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11728__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13350_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout202_A _06901_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 hold330/X vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__buf_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_09924_ _09925_/A _09925_/B _09809_/X vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09855_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__A1 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10703__B2 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _08805_/B _08805_/C _08805_/A vssd1 vssd1 vccd1 vccd1 _08809_/C sky130_fd_sc_hd__a21oi_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06998_ _07299_/B _07050_/A _07050_/B _06964_/B vssd1 vssd1 vccd1 vccd1 _07000_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__07580__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ fanout58/X fanout85/X _10466_/A fanout57/X vssd1 vssd1 vccd1 vccd1 _09787_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07064__A _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ _08731_/X _10896_/B _11011_/C vssd1 vssd1 vccd1 vccd1 _08737_/Y sky130_fd_sc_hd__nand3b_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10467__B1 _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _08669_/A _08669_/B _08720_/A vssd1 vssd1 vccd1 vccd1 _08670_/C sky130_fd_sc_hd__a21o_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ _08891_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__and2_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10518_/A _10518_/B _10516_/X vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08599_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08599_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ _07218_/A _11446_/B _09235_/X _06749_/B _12504_/S vssd1 vssd1 vccd1 vccd1
+ _10561_/X sky130_fd_sc_hd__o221a_1
X_10492_ _10491_/A _10491_/B _10491_/C vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__a21oi_1
X_12300_ _06613_/X _11966_/B _12299_/Y _06615_/B _06940_/B vssd1 vssd1 vccd1 vccd1
+ _12300_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ _13287_/CLK _13280_/D vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12162_ _12162_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12093_ _12019_/Y _12374_/D _12280_/A vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__a21oi_1
X_11113_ _10653_/B _11112_/Y _11111_/Y vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__o21ai_4
X_11044_ _10958_/A _10958_/B _10955_/A vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12799__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12995_ hold218/X _13143_/B2 _13186_/A2 hold199/X vssd1 vssd1 vccd1 vccd1 hold219/A
+ sky130_fd_sc_hd__a22o_1
X_11946_ _11946_/A _11946_/B vssd1 vssd1 vccd1 vccd1 _11972_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ hold299/A _11877_/B vssd1 vssd1 vccd1 vccd1 _11963_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10828_ _12068_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _10759_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11422__A2 _11451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A3 _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08533__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12055__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ reg1_val[31] _07127_/B _09595_/B vssd1 vssd1 vccd1 vccd1 _12429_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07970_ _08566_/A _07970_/B _07970_/C vssd1 vssd1 vccd1 vccd1 _07973_/B sky130_fd_sc_hd__and3_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06921_ instruction[21] _06575_/X _06920_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08354__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06852_ reg1_val[27] _07029_/A vssd1 vssd1 vccd1 vccd1 _06852_/Y sky130_fd_sc_hd__nand2_1
X_09640_ _09517_/A _09517_/B _09514_/A vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07562__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06783_ _06799_/A _06801_/B1 _12637_/B _06781_/X vssd1 vssd1 vccd1 vccd1 _07145_/A
+ sky130_fd_sc_hd__a31o_4
X_09571_ _09187_/X _09212_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ _08566_/A _08522_/B vssd1 vssd1 vccd1 vccd1 _08528_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08453_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08461_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout152_A _06995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07404_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _08384_/A _08428_/A vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08814__B1 _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ _07114_/X _07539_/B fanout37/X _07146_/Y vssd1 vssd1 vccd1 vccd1 _07336_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _09630_/A _07266_/B vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09064_/C sky130_fd_sc_hd__and2_1
XFILLER_0_103_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07197_ _07195_/A _07194_/X _07195_/Y _06963_/A vssd1 vssd1 vccd1 vccd1 _07197_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__10924__A1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07059__A _07060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09907_ _09814_/A _09814_/B _09813_/A vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10213__A _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__nand2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10432__A1_N _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _09769_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__or2_1
X_11800_ _11795_/Y _11796_/X _11799_/X _11793_/X vssd1 vssd1 vccd1 vccd1 _11800_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12780_ rst _12780_/B _12780_/C vssd1 vssd1 vccd1 vccd1 _13240_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07305__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _11730_/B _11731_/B vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _11562_/A _11562_/B _11570_/B _11571_/B _11571_/A vssd1 vssd1 vccd1 vccd1
+ _11675_/A sky130_fd_sc_hd__a32oi_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11593_ _11593_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__nand2_4
X_10613_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10612__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ _13344_/CLK hold128/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_10544_ _06878_/A _10543_/X _11612_/A vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13263_ _13363_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13277__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ hold289/X _13193_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_1
X_12214_ _12324_/A _12270_/A vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_102_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12145_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12212_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ _12077_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12151_/A sky130_fd_sc_hd__nand2_1
X_11027_ hold330/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11243_/C sky130_fd_sc_hd__or2_1
XANTENNA__11876__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12978_ _12978_/A hold260/X vssd1 vssd1 vccd1 vccd1 _13287_/D sky130_fd_sc_hd__and2_1
XANTENNA__09297__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07432__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _11930_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09049__B1 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_17 reg2_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 reg2_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_39 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07120_ reg1_val[23] _12717_/B _07120_/C vssd1 vssd1 vccd1 vccd1 _07123_/A sky130_fd_sc_hd__or3_4
XFILLER_0_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__B2 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13148__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ _07891_/B _07891_/C vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__and2_4
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12513__A _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07953_ _07953_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _07954_/B sky130_fd_sc_hd__and2_1
XANTENNA__07607__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06904_ instruction[2] instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _06907_/B sky130_fd_sc_hd__and4b_4
XANTENNA__11129__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ _07985_/A _07985_/B _07881_/A vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__a21oi_1
X_06835_ reg1_val[17] _11446_/A vssd1 vssd1 vccd1 vccd1 _06835_/X sky130_fd_sc_hd__and2_1
X_09623_ _11386_/A fanout27/X fanout25/X fanout83/X vssd1 vssd1 vccd1 vccd1 _09624_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11619__C1 _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06766_ _06567_/Y _06593_/X _06596_/Y _12647_/B _06908_/A vssd1 vssd1 vccd1 vccd1
+ _06766_/X sky130_fd_sc_hd__o2111a_1
X_09554_ _08656_/B _08708_/B _09554_/S vssd1 vssd1 vccd1 vccd1 _09554_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09541__B _09543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06697_ _11531_/S _06698_/B vssd1 vssd1 vccd1 vccd1 _06697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09485_ _09787_/A _09485_/B vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ _08594_/A2 _09468_/B2 _08591_/B1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08506_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08436_ _08594_/A2 _08553_/A2 _08553_/B1 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08437_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08367_ _08619_/B1 _08400_/B fanout82/X _09403_/S vssd1 vssd1 vccd1 vccd1 _08368_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07318_ fanout62/X _08590_/B _09648_/A fanout60/X vssd1 vssd1 vccd1 vccd1 _07319_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08298_ _08298_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__xnor2_2
X_07249_ _11071_/A _11070_/A vssd1 vssd1 vccd1 vccd1 _07249_/Y sky130_fd_sc_hd__nand2_1
X_10260_ _10261_/A _10261_/B vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__and2_1
XFILLER_0_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09763__A1 _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10373__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__B2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10192_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09208__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__A1 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ hold15/X hold313/A vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07526__B1 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _11917_/B _12782_/Y hold102/X _13226_/A vssd1 vssd1 vccd1 vccd1 hold103/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12822__A1 _07067_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A _12763_/B vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__nand2_2
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11709_/Y _11710_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11715_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ _12694_/A _12694_/B _12694_/C vssd1 vssd1 vccd1 vccd1 _12695_/B sky130_fd_sc_hd__nand3_1
X_11645_ _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _11576_/A _11576_/B _11574_/Y vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__or3b_1
X_10527_ _10529_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or2_1
X_13315_ _13324_/CLK hold169/X vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10458_ _10458_/A _10458_/B _10458_/C vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__and3_1
X_13246_ _13341_/CLK _13246_/D vssd1 vssd1 vccd1 vccd1 hold104/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07214__C1 _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13177_ hold302/X _13209_/A2 _13176_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 _13178_/B
+ sky130_fd_sc_hd__a22o_1
X_10389_ _10192_/A _10192_/B _10190_/X vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10552__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _12075_/A _12075_/B _12074_/A vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__a21o_1
X_12059_ _12059_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06620_ reg1_val[30] _08971_/C vssd1 vssd1 vccd1 vccd1 _12415_/B sky130_fd_sc_hd__and2_1
XANTENNA__13066__A1 _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _09507_/A _09270_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__or2_1
XANTENNA__07296__A2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11115__C _11258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _09468_/B2 _08400_/B fanout82/X _08591_/B1 vssd1 vssd1 vccd1 vccd1 _08222_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08150_/A _08150_/B _08151_/Y vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07103_ reg1_val[20] _07229_/B _07190_/B reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07109_/B
+ sky130_fd_sc_hd__a211oi_4
X_08083_ _08083_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ fanout62/X _09300_/A fanout56/X _08633_/B vssd1 vssd1 vccd1 vccd1 _07035_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _12378_/S _08983_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _08985_/Y sky130_fd_sc_hd__o21ai_4
X_07936_ _07936_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07940_/A sky130_fd_sc_hd__nor2_1
X_07867_ _07867_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__and2_1
X_06818_ _10414_/A _06816_/X _06817_/X vssd1 vssd1 vccd1 vccd1 _06818_/X sky130_fd_sc_hd__a21o_1
X_09606_ _09503_/A _09503_/B _09501_/Y vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__a21o_2
X_07798_ _07860_/B _07860_/A vssd1 vssd1 vccd1 vccd1 _07798_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11068__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__A1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _06747_/Y _06749_/B vssd1 vssd1 vccd1 vccd1 _06878_/A sky130_fd_sc_hd__nand2b_1
X_09537_ _09537_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09815_/A fanout9/A fanout5/X _09468_/B2 vssd1 vssd1 vccd1 vccd1 _09469_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07287__A2 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _09201_/X _09203_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09399_/X sky130_fd_sc_hd__mux2_1
X_08419_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08425_/A sky130_fd_sc_hd__nor2_1
X_11430_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11430_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08236__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10043__A1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13100_ _13109_/A hold318/X vssd1 vssd1 vccd1 vccd1 _13342_/D sky130_fd_sc_hd__and2_1
X_10312_ _10136_/A _10136_/B _09710_/Y vssd1 vssd1 vccd1 vccd1 _10313_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11292_ _11173_/A _11173_/B _11170_/A vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10346__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _10243_/A _10243_/B _10243_/C vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__or3_1
X_13031_ hold186/A _13055_/A2 _13053_/B1 hold178/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold179/A sky130_fd_sc_hd__o221a_1
XANTENNA__07247__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10438_/C _10173_/Y _12490_/S _10171_/X vssd1 vssd1 vccd1 vccd1 dest_val[6]
+ sky130_fd_sc_hd__a2bb2o_4
Xfanout170 _09152_/Y vssd1 vssd1 vccd1 vccd1 _09155_/S sky130_fd_sc_hd__clkbuf_8
Xfanout181 _12847_/B vssd1 vssd1 vccd1 vccd1 _13052_/A2 sky130_fd_sc_hd__buf_2
Xfanout192 _08650_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__buf_8
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12815_ hold80/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__or2_1
XANTENNA__06708__A_N _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ _12744_/X _12746_/B vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__07710__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12682_/B _12677_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
XFILLER_0_127_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _09196_/S _10904_/Y _10922_/Y _09223_/Y _11627_/X vssd1 vssd1 vccd1 vccd1
+ _11628_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _11559_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11561_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10585__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ hold193/X _12780_/B _12774_/Y _06564_/A vssd1 vssd1 vccd1 vccd1 _13229_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12063__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__A1 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07157__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06996__A _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _11604_/B _11604_/C _11693_/A vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__and3_1
XFILLER_0_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07721_ _07721_/A _07721_/B _07721_/C vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__and3_1
X_07652_ _07487_/A _07487_/B _07485_/Y vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ reg2_val[29] _06794_/B _06707_/B1 _06602_/Y vssd1 vssd1 vccd1 vccd1 _06850_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_07583_ _11813_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09322_ _09322_/A vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07269__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__A1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__B2 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout232_A _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _09217_/Y _09223_/Y _09252_/X _09196_/S _09242_/Y vssd1 vssd1 vccd1 vccd1
+ _09253_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09415__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09184_ _09168_/X _10421_/B _11235_/S vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _08204_/A _08204_/B _08207_/B vssd1 vssd1 vccd1 vccd1 _08204_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11222__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__or2_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07441__A2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _08066_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08067_/C sky130_fd_sc_hd__and2_1
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ _07011_/A _07011_/B _09671_/A vssd1 vssd1 vccd1 vccd1 _07017_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08968_ _09062_/B _08968_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__nand2_1
X_08899_ _07644_/A _07644_/B _07643_/A vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__a21o_1
X_07919_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__xnor2_1
X_10930_ _11386_/A fanout22/X fanout15/X _11296_/A vssd1 vssd1 vccd1 vccd1 _10931_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _12600_/A _12600_/B _12600_/C _12600_/D vssd1 vssd1 vccd1 vccd1 _12601_/B
+ sky130_fd_sc_hd__and4_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10861_ _10862_/A _10862_/B _10862_/C vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10792_ _11115_/A _10912_/B hold207/A vssd1 vssd1 vccd1 vccd1 _10792_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09654__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11461__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12537_/B _12531_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
XFILLER_0_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11052__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ reg1_val[4] curr_PC[4] _12504_/S vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11413_ _11413_/A _11504_/A vssd1 vssd1 vccd1 vccd1 _11597_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07680__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ hold324/A _12349_/A _12391_/X _12393_/B1 vssd1 vssd1 vccd1 vccd1 _12393_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11344_ _06711_/A _09886_/B _12395_/A1 vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12961__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11276_/B sky130_fd_sc_hd__and2_1
X_13014_ _13226_/A hold163/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__and2_1
X_10226_ _10055_/A _10053_/Y _10052_/Y vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07196__A1 _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _10158_/A2 _10292_/B hold309/A vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__a21oi_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10088_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12244__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _12721_/Y _12725_/B _12723_/B vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__o21a_2
XANTENNA__07440__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09948__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A1 _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09948__B2 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap112 _10213_/A vssd1 vssd1 vccd1 vccd1 _09450_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12505__B _12506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09940_ _10234_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__xnor2_4
X_09871_ _12025_/S _06808_/Y _09870_/Y vssd1 vssd1 vccd1 vccd1 _09871_/X sky130_fd_sc_hd__o21a_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _09766_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08823_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06767__C_N _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout182_A _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _07739_/A _07739_/B _07700_/X vssd1 vssd1 vccd1 vccd1 _07712_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08684_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08751_/C sky130_fd_sc_hd__nor2_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11691__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _08831_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07637_/C sky130_fd_sc_hd__or2_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _09670_/A _09305_/B _09305_/C vssd1 vssd1 vccd1 vccd1 _09306_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _12029_/A _11966_/B _08655_/A vssd1 vssd1 vccd1 vccd1 _09236_/X sky130_fd_sc_hd__o21a_1
X_07497_ _07500_/A _07500_/B vssd1 vssd1 vccd1 vccd1 _07497_/X sky130_fd_sc_hd__or2_1
XANTENNA__09939__A1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09167_ _09163_/X _09166_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09098_ _09329_/B _09098_/B vssd1 vssd1 vccd1 vccd1 _09099_/B sky130_fd_sc_hd__and2_2
X_08118_ _08507_/A2 _08521_/A2 _08926_/B1 _08533_/B vssd1 vssd1 vccd1 vccd1 _08119_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ _08049_/A _08049_/B _08049_/C vssd1 vssd1 vccd1 vccd1 _08050_/B sky130_fd_sc_hd__nand3_1
X_11060_ _11060_/A _11060_/B vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _09383_/X _09387_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10011_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08375__B1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11962_ hold204/A _12178_/A2 _12037_/B _11961_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _11971_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10913_ _11115_/A _11024_/B hold220/A vssd1 vssd1 vccd1 vccd1 _10913_/Y sky130_fd_sc_hd__a21oi_1
X_11893_ _12615_/S _11893_/B _12051_/C vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__or3_2
XFILLER_0_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844_ _11557_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__B2 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__A1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ _12523_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12516_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10775_ _10541_/B _10541_/C _10657_/A _11776_/A vssd1 vssd1 vccd1 vccd1 _10776_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12445_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12453_/B sky130_fd_sc_hd__or2_1
X_12376_ _12280_/A _12373_/Y _12374_/X _09148_/Y vssd1 vssd1 vccd1 vccd1 _12376_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08091__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _11115_/A _11259_/X _11451_/A _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11327_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _11258_/A _11258_/B vssd1 vssd1 vccd1 vccd1 _11809_/C sky130_fd_sc_hd__or2_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _11189_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__xnor2_1
X_10209_ _07218_/Y _08873_/X _08988_/Y _10326_/A vssd1 vssd1 vccd1 vccd1 _10210_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10173__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07435__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08118__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09650__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07892__A2 _07060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _07425_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07170__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ _07351_/A _07351_/B vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11976__A1 _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07282_ _07282_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11728__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__B2 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10951__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold326/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold325/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _09793_/A _09793_/B _09792_/A vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__xnor2_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__A _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _08805_/A _08805_/B _08805_/C vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__and3_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _06996_/A _06967_/A _07074_/B _06681_/B vssd1 vssd1 vccd1 vccd1 _07000_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__07580__A1 _12193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ _10230_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__xnor2_1
X_08736_ _08736_/A _08736_/B vssd1 vssd1 vccd1 vccd1 _11011_/C sky130_fd_sc_hd__xnor2_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09560__A _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _08616_/A _08718_/B _08616_/B vssd1 vssd1 vccd1 vccd1 _08720_/A sky130_fd_sc_hd__o21ba_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ _07618_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07619_/B sky130_fd_sc_hd__or2_1
XFILLER_0_119_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__or2_1
XANTENNA__07080__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07549_ _07550_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _07549_/Y sky130_fd_sc_hd__nand2_1
X_10560_ hold303/A _12349_/A _10677_/B _12393_/B1 vssd1 vssd1 vccd1 vccd1 _10560_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ _10491_/A _10491_/B _10491_/C vssd1 vssd1 vccd1 vccd1 _10493_/A sky130_fd_sc_hd__and3_1
X_09219_ _09219_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09219_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12170_/A _12167_/Y _12169_/B vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _06866_/X _12160_/X _12378_/S vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__mux2_1
X_12092_ _12324_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__xnor2_2
X_11112_ _11112_/A _11322_/A vssd1 vssd1 vccd1 vccd1 _11112_/Y sky130_fd_sc_hd__nand2_1
X_11043_ _10990_/A _10990_/B _10988_/Y vssd1 vssd1 vccd1 vccd1 _11105_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07255__A _07255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _13144_/A hold250/X vssd1 vssd1 vccd1 vccd1 _13295_/D sky130_fd_sc_hd__and2_1
X_11945_ _11945_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ _11958_/A _10565_/A _11875_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _11876_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08086__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ _07968_/B _07402_/B fanout41/X _07077_/X vssd1 vssd1 vccd1 vccd1 _10828_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10758_ _10759_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12428_ hold174/A _12426_/X _12427_/Y vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _12053_/A1 _10685_/X _10688_/X vssd1 vssd1 vccd1 vccd1 dest_val[10] sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08533__B _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _08874_/A fanout6/X _12404_/B vssd1 vssd1 vccd1 vccd1 _12359_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06920_ instruction[28] _06922_/B vssd1 vssd1 vccd1 vccd1 _06920_/X sky130_fd_sc_hd__or2_1
X_06851_ reg1_val[28] _06851_/B vssd1 vssd1 vccd1 vccd1 _06851_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07562__A1 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__B2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ _06799_/A _06801_/B1 _12637_/B _06781_/X vssd1 vssd1 vccd1 vccd1 _07146_/A
+ sky130_fd_sc_hd__a31oi_4
X_09570_ _09205_/X _09209_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__mux2_1
X_08521_ _06875_/A _08521_/A2 _08551_/A2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08522_/B
+ sky130_fd_sc_hd__o22a_1
X_08452_ _08477_/A _08477_/B _08490_/B _08451_/B _08451_/A vssd1 vssd1 vccd1 vccd1
+ _08461_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07403_ _10937_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout145_A _07054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08428_/A sky130_fd_sc_hd__or2_1
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07334_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08814__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08814__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ _07944_/B _09450_/B1 _07263_/Y fanout28/X vssd1 vssd1 vccd1 vccd1 _07266_/B
+ sky130_fd_sc_hd__a22o_1
X_09004_ _09630_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ _07195_/A _07194_/X _07195_/Y _06963_/A vssd1 vssd1 vccd1 vccd1 _10326_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07059__B _07060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09906_ _09849_/A _09849_/B _09850_/Y vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__10213__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09837_/Y sky130_fd_sc_hd__nor2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12429__A2 _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _09767_/B _09768_/B vssd1 vssd1 vccd1 vccd1 _09769_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11637__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__C1 _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _10276_/B _10276_/C vssd1 vssd1 vccd1 vccd1 _08721_/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout58_A _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ _11731_/B _11730_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__xnor2_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07305__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07305__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11661_/A _11661_/B vssd1 vssd1 vccd1 vccd1 _11677_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11592_ _11592_/A _11592_/B _11592_/C vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12062__B1 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ fanout82/X fanout13/X fanout12/X _07236_/Y vssd1 vssd1 vccd1 vccd1 _10613_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10612__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13331_ _13334_/CLK hold133/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
X_10543_ _06818_/X _10542_/X _12025_/S vssd1 vssd1 vccd1 vccd1 _10543_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _13364_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
X_10474_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08569__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ _13193_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__xnor2_1
X_12213_ _12213_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__and2_1
XANTENNA__09230__A1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _12202_/D _12144_/B vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07241__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _12075_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12077_/B sky130_fd_sc_hd__xor2_1
X_11026_ hold259/A _11115_/A _11134_/B _11025_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _11033_/A sky130_fd_sc_hd__a311o_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12977_ hold220/X _13095_/B2 _13158_/A2 hold259/X vssd1 vssd1 vccd1 vccd1 hold260/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09297__A1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__B2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11928_ _11928_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ _11114_/B _11506_/X _11857_/Y _11858_/X vssd1 vssd1 vccd1 vccd1 _11860_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__09049__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 reg2_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 reg2_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07050_ _07050_/A _07050_/B vssd1 vssd1 vccd1 vccd1 _07891_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08272__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09221__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__A _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _07902_/A _07902_/B _07899_/Y vssd1 vssd1 vccd1 vccd1 _07955_/B sky130_fd_sc_hd__o21bai_1
X_06903_ hold184/A _12780_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
X_07883_ _09795_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13069__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ _11333_/A _06832_/Y _06833_/X vssd1 vssd1 vccd1 vccd1 _06834_/X sky130_fd_sc_hd__a21o_1
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__or2_1
X_09553_ _12420_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09554_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06765_ _06765_/A _06765_/B vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09288__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__xnor2_1
X_06696_ reg1_val[18] _07068_/A vssd1 vssd1 vccd1 vccd1 _06698_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ fanout62/X fanout85/X _10466_/A fanout60/X vssd1 vssd1 vccd1 vccd1 _09485_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _08438_/A _08438_/B vssd1 vssd1 vccd1 vccd1 _08435_/X sky130_fd_sc_hd__or2_1
X_08366_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08366_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07317_ _10230_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07321_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08297_ _08333_/A _08333_/B _08286_/Y vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ _09787_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07179_ _07179_/A _07179_/B vssd1 vssd1 vccd1 vccd1 _07179_/X sky130_fd_sc_hd__xor2_4
X_10190_ _10191_/B _10191_/A vssd1 vssd1 vccd1 vccd1 _10190_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09515__A2 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _13110_/A _13111_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08869__A4 _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ hold101/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07533__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__A2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12822__A2 _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12762_ reg1_val[29] _12767_/B vssd1 vssd1 vccd1 vccd1 _12763_/B sky130_fd_sc_hd__nand2_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ _09196_/S _10789_/X _10801_/Y _09223_/Y _11712_/X vssd1 vssd1 vccd1 vccd1
+ _11713_/X sky130_fd_sc_hd__o221a_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12693_ _12694_/A _12694_/B _12694_/C vssd1 vssd1 vccd1 vccd1 _12698_/B sky130_fd_sc_hd__a21o_1
X_11644_ _11837_/A fanout9/X fanout4/X fanout61/X vssd1 vssd1 vccd1 vccd1 _11734_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11575_ _11576_/A _11576_/B _11574_/Y vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__10597__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _10526_/A _10526_/B vssd1 vssd1 vccd1 vccd1 _10529_/B sky130_fd_sc_hd__xor2_4
X_13314_ _13324_/CLK hold180/X vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10457_ _10458_/A _10458_/B _10458_/C vssd1 vssd1 vccd1 vccd1 _10635_/A sky130_fd_sc_hd__a21oi_1
X_13245_ _13341_/CLK _13245_/D vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07708__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ hold275/X _13175_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__mux2_1
X_10388_ _10248_/A _10247_/B _10247_/A vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12127_ _12374_/D _12279_/B _12280_/A vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__a21o_1
X_12058_ _12058_/A _12058_/B vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11009_ _10929_/X _11041_/C _11008_/Y vssd1 vssd1 vccd1 vccd1 _11009_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13066__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ _08212_/B _08212_/A vssd1 vssd1 vccd1 vccd1 _08151_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07102_ reg1_val[20] _07087_/X _12717_/B reg1_val[21] _07229_/B vssd1 vssd1 vccd1
+ vccd1 _07109_/A sky130_fd_sc_hd__o311a_2
XFILLER_0_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08082_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08140_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07033_ _09670_/A _07033_/B vssd1 vssd1 vccd1 vccd1 _07037_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout108_A _09114_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08984_ _12378_/S _08983_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _11917_/C sky130_fd_sc_hd__o21a_4
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08953__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ _07935_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__and2_1
XFILLER_0_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07866_ _07826_/A _07825_/B _07825_/C vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__a21o_1
X_09605_ _09535_/A _09535_/B _09536_/Y vssd1 vssd1 vccd1 vccd1 _09702_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__08449__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06817_ _07195_/A reg1_val[8] vssd1 vssd1 vccd1 vccd1 _06817_/X sky130_fd_sc_hd__and2b_1
X_07797_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07860_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11068__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__A2 _12782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06748_ reg1_val[9] _07217_/A vssd1 vssd1 vccd1 vccd1 _06749_/B sky130_fd_sc_hd__nand2_1
X_09536_ _09537_/B _09537_/A vssd1 vssd1 vccd1 vccd1 _09536_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _09467_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__nor2_1
X_06679_ _06964_/B vssd1 vssd1 vccd1 vccd1 _06681_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ _08426_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ _09395_/X _09397_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _09398_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08184__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__B1 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08236__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08349_ _08311_/Y _08348_/Y _08310_/Y vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__a21o_1
X_11360_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__and2_1
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__A2 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__C _11041_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07444__B1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _09864_/A _09864_/B _09440_/C vssd1 vssd1 vccd1 vccd1 _10313_/C sky130_fd_sc_hd__o21bai_1
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__xnor2_2
X_13030_ _09938_/A _12797_/B hold187/X vssd1 vssd1 vccd1 vccd1 _13313_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10242_ _10372_/B _10241_/C _10241_/A vssd1 vssd1 vccd1 vccd1 _10243_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07247__B _07248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ curr_PC[6] _10172_/B _12053_/A1 vssd1 vssd1 vccd1 vccd1 _10173_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout182 _12839_/B vssd1 vssd1 vccd1 vccd1 _12847_/B sky130_fd_sc_hd__buf_2
Xfanout160 _06942_/Y vssd1 vssd1 vccd1 vccd1 _10427_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout171 _07910_/A vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__buf_12
Xfanout193 _06987_/Y vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__clkbuf_16
X_12814_ _07250_/X _12842_/A2 hold54/X _13187_/A vssd1 vssd1 vccd1 vccd1 hold55/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ reg1_val[26] _12773_/A vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07683__B1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11627_ _12395_/A1 _11626_/X _06690_/B vssd1 vssd1 vccd1 vccd1 _11627_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ fanout29/X _08857_/Y wire8/X _07193_/Y vssd1 vssd1 vccd1 vccd1 _11559_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10509_ _10509_/A _10509_/B _10509_/C vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__and3_1
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08822__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _11489_/A _11489_/B vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13228_ hold149/X _12781_/A _13236_/A hold150/X vssd1 vssd1 vccd1 vccd1 hold151/A
+ sky130_fd_sc_hd__o211a_1
X_13159_ _13187_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13354_/D sky130_fd_sc_hd__and2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _07522_/A _07522_/C _07522_/B vssd1 vssd1 vccd1 vccd1 _07721_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__xnor2_4
X_06602_ _06706_/A _12691_/B vssd1 vssd1 vccd1 vccd1 _06602_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06713__A2 _06591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07582_ _09324_/A _07347_/B fanout15/X _12785_/A vssd1 vssd1 vccd1 vccd1 _07583_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12798__A1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09322_/A sky130_fd_sc_hd__and2_1
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09112__B1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__A _12679_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08466__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _09252_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__or2_2
XANTENNA__10273__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ _09175_/X _09182_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__mux2_1
X_08203_ _08203_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__and2_1
X_08134_ _08134_/A _08134_/B vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09179__A0 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__nand2_1
X_07016_ _07016_/A _07016_/B vssd1 vssd1 vccd1 vccd1 _11917_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08926__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _08967_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _08968_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08898_ _08898_/A _08898_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__xor2_2
X_07918_ _07918_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07925_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07849_ _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__and2b_1
X_10860_ _10860_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10862_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout40_A fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _09520_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09103__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ hold240/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10912_/B sky130_fd_sc_hd__or2_1
XANTENNA__09654__A1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__B2 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11461__B2 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A1 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ _12530_/A _12530_/B _12530_/C vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _12467_/B _12461_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11412_ _11410_/Y _11412_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12392_ _12349_/A _12391_/X hold324/A vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08642__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11343_ hold320/A _11879_/A2 _11524_/C _11342_/Y _12175_/C1 vssd1 vssd1 vccd1 vccd1
+ _11343_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08090__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__nor2_1
X_13013_ hold263/A _06564_/A _13222_/A2 hold162/X vssd1 vssd1 vccd1 vccd1 hold163/A
+ sky130_fd_sc_hd__a22o_1
X_10225_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__xnor2_1
X_10156_ hold293/A hold317/A _10156_/C vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__or3_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _09936_/A _09936_/B _09933_/A vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06825__A_N _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08817__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _10989_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09645__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08448__A2 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12728_ _12728_/A _12728_/B vssd1 vssd1 vccd1 vccd1 _12737_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12659_ _12659_/A _12659_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
XFILLER_0_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09648__A _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08552__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap102 _07067_/Y vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__buf_4
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _12025_/S _09870_/B vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06919__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _07101_/Y fanout37/X _07263_/Y _07539_/B vssd1 vssd1 vccd1 vccd1 _08822_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08751_/A _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__a21oi_1
X_08683_ _08683_/A _08683_/B _08683_/C vssd1 vssd1 vccd1 vccd1 _08685_/B sky130_fd_sc_hd__and3_1
X_07703_ _08320_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__xnor2_4
X_07634_ _07634_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _07565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__A1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _09305_/B _09305_/C _09670_/A vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__a21o_1
X_07496_ _11168_/A _07496_/B vssd1 vssd1 vccd1 vccd1 _07500_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09235_ _09235_/A instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09235_/X
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09939__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09164_/X _09165_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09097_ _09097_/A _09097_/B vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__or2_1
X_08117_ _08200_/A _08200_/B _08109_/X vssd1 vssd1 vccd1 vccd1 _08138_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08048_ _08048_/A _08048_/B _08048_/C vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__and3_1
XANTENNA_fanout88_A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _11237_/S _10009_/Y _09252_/A vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__09293__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__B2 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _09375_/B _09996_/Y _09998_/X vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__a21boi_2
X_11961_ _12178_/A2 _12037_/B hold204/A vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07017__S _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10912_ hold207/A _10912_/B vssd1 vssd1 vccd1 vccd1 _11024_/B sky130_fd_sc_hd__or2_1
XANTENNA__09875__A1 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11892_ curr_PC[21] curr_PC[22] _11892_/C vssd1 vssd1 vccd1 vccd1 _12051_/C sky130_fd_sc_hd__and3_1
XANTENNA__07886__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10843_ _12202_/A fanout27/X fanout25/X fanout64/X vssd1 vssd1 vccd1 vccd1 _10844_/B
+ sky130_fd_sc_hd__o22a_1
X_10774_ _10774_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10774_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11985__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _12673_/B _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__or2_1
XFILLER_0_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12444_ _12453_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _12446_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _12280_/A _12374_/X _12373_/Y vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ _11115_/A _11259_/X _11451_/A vssd1 vssd1 vccd1 vccd1 _11326_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _12490_/S _11253_/X _11254_/X _11256_/Y vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__a22o_4
X_11188_ _11188_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _11189_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11370__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__xnor2_1
X_10139_ _10315_/A _10140_/B _10140_/C vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08118__B2 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07877__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07629__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ _07574_/A _07350_/B vssd1 vssd1 vccd1 vccd1 _07351_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07281_ _07281_/A _07281_/B vssd1 vssd1 vccd1 vccd1 _08476_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09022_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_127_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11728__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold279 hold324/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xor2_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _12202_/A _10463_/B2 _10228_/A fanout64/X vssd1 vssd1 vccd1 vccd1 _09785_/B
+ sky130_fd_sc_hd__o22a_1
X_08804_ _08796_/B _08796_/C _08803_/A _08803_/B vssd1 vssd1 vccd1 vccd1 _08805_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout292_A _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _06996_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _07050_/B sky130_fd_sc_hd__nor2_1
X_08735_ _08731_/X _10896_/B vssd1 vssd1 vccd1 vccd1 _11011_/B sky130_fd_sc_hd__and2b_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11664__A1 _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08666_ _08666_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _08716_/B sky130_fd_sc_hd__or2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08597_ _08597_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__xnor2_2
X_07617_ _07618_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07548_ _07548_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07550_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07479_ _07551_/A _07551_/B _07478_/A vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _10490_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _10491_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09218_ _09219_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08192__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _09235_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__or2_2
XFILLER_0_17_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12098_/A _12096_/X _12115_/S vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10927__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _10887_/Y _11322_/A _11109_/X vssd1 vssd1 vccd1 vccd1 _11111_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _11420_/B _12087_/Y _12088_/Y _12325_/B vssd1 vssd1 vccd1 vccd1 _12092_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12442__A _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ _11809_/A _11809_/B vssd1 vssd1 vccd1 vccd1 _11259_/A sky130_fd_sc_hd__or2_1
XANTENNA__09545__B1 _09370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ hold225/X _13143_/B2 _13186_/A2 hold218/X vssd1 vssd1 vccd1 vccd1 hold250/A
+ sky130_fd_sc_hd__a22o_1
X_11944_ _11776_/B _11777_/A _11864_/A _11776_/A vssd1 vssd1 vccd1 vccd1 _11945_/B
+ sky130_fd_sc_hd__a31o_1
X_11875_ _11958_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10826_ _10826_/A _10826_/B vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10757_ _10757_/A _10757_/B vssd1 vssd1 vccd1 vccd1 _10759_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13212__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _12490_/S _10926_/C _10688_/C vssd1 vssd1 vccd1 vccd1 _10688_/X sky130_fd_sc_hd__or3_2
X_12427_ hold174/A _12426_/X _09239_/Y vssd1 vssd1 vccd1 vccd1 _12427_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09784__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _12310_/A _12310_/B _12313_/A vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__xnor2_2
X_12289_ _12234_/A _12231_/Y _12233_/B vssd1 vssd1 vccd1 vccd1 _12341_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06850_ reg1_val[29] _06850_/B vssd1 vssd1 vccd1 vccd1 _06850_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11894__A1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1_N _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06781_ reg2_val[3] _06794_/B vssd1 vssd1 vccd1 vccd1 _06781_/X sky130_fd_sc_hd__and2_1
X_08520_ _08520_/A _08520_/B vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__xnor2_1
X_08451_ _08451_/A _08451_/B vssd1 vssd1 vccd1 vccd1 _08490_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _08476_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07403_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08382_ _08384_/A _08382_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12527__A _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07333_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08814__A2 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13122__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A _10613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07264_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _10712_/A _07944_/B fanout28/X _07212_/X vssd1 vssd1 vccd1 vccd1 _09004_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10047__A _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _07195_/A _07195_/B vssd1 vssd1 vccd1 vccd1 _07195_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _09854_/A _09854_/B _09852_/X vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11885__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ _09836_/A _09836_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__xnor2_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _09768_/B _09767_/B vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__and2b_1
X_06979_ _06973_/A fanout67/X _08551_/B2 fanout64/X vssd1 vssd1 vccd1 vccd1 _06980_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11637__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ _09699_/B _09699_/A vssd1 vssd1 vccd1 vccd1 _09698_/Y sky130_fd_sc_hd__nand2b_1
X_08718_ _08718_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _10276_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _09403_/S _08649_/B vssd1 vssd1 vccd1 vccd1 _08659_/S sky130_fd_sc_hd__nor2_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07305__A2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11748_/B _11660_/B vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__or2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11591_ _11593_/A vssd1 vssd1 vccd1 vccd1 _11591_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12062__A1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ _10494_/A _10493_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _10626_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10612__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ _13334_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
X_10542_ _06752_/Y _10412_/X _06754_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__o21a_1
X_13261_ _13364_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08018__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__B1 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ _10355_/A _10355_/B _10352_/A vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__a21o_1
X_12212_ _12212_/A _12212_/B _12212_/C vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__or3_1
XANTENNA__08569__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ _13226_/A hold290/X vssd1 vssd1 vccd1 vccd1 _13361_/D sky130_fd_sc_hd__and2_1
XANTENNA__08650__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12143_ _12143_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07241__A1 _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _12074_/A _12074_/B vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07266__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _11115_/A _11134_/B hold259/A vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10404__B _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__A1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__B1 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11628__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ _12978_/A hold221/X vssd1 vssd1 vccd1 vccd1 _13286_/D sky130_fd_sc_hd__and2_1
XANTENNA__09297__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ _11928_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__nand2_1
X_11858_ _11505_/X _11856_/A _12016_/A _11855_/X vssd1 vssd1 vccd1 vccd1 _11858_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09049__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _11238_/S _10682_/Y _11788_/Y _09243_/B vssd1 vssd1 vccd1 vccd1 _11789_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_19 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12053__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _12490_/S _10805_/X _10806_/X _10808_/Y vssd1 vssd1 vccd1 vccd1 dest_val[11]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07951_ _07951_/A _08046_/A vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__or2_1
XFILLER_0_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06902_ _12782_/A _12781_/B vssd1 vssd1 vccd1 vccd1 _13227_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ _09675_/A _08096_/B fanout24/X _09467_/A vssd1 vssd1 vccd1 vccd1 _07883_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06833_ reg1_val[16] _07074_/A vssd1 vssd1 vccd1 vccd1 _06833_/X sky130_fd_sc_hd__and2_1
X_09621_ _09621_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13117__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11619__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06764_ reg1_val[6] _07264_/A vssd1 vssd1 vccd1 vccd1 _06765_/B sky130_fd_sc_hd__and2_1
X_09552_ _09552_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09552_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09288__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ _08520_/A _08502_/Y _08498_/X vssd1 vssd1 vccd1 vccd1 _08510_/A sky130_fd_sc_hd__o21a_1
XANTENNA_fanout255_A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ reg1_val[18] _07068_/A vssd1 vssd1 vccd1 vccd1 _11531_/S sky130_fd_sc_hd__and2_1
XANTENNA__12292__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07342__C _07342_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__B1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ _09941_/A _08434_/B vssd1 vssd1 vccd1 vccd1 _08438_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12044__A1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ _10735_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08370_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12257__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07316_ _09659_/B2 _10463_/B2 _10228_/A fanout98/X vssd1 vssd1 vccd1 vccd1 _07317_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ _09787_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _11071_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07178_ _07179_/A _07179_/B vssd1 vssd1 vccd1 vccd1 _07178_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09748__B1 _09239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09819_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07814__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _06993_/Y _12842_/A2 hold78/X _13187_/A vssd1 vssd1 vccd1 vccd1 hold79/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12761_ reg1_val[29] _12767_/B vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__or2_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ _12395_/A1 _11711_/X _06675_/B vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__a21o_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12692_ _12698_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _12694_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11643_ _11753_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10046__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11574_ _11470_/A _11470_/B _11467_/A vssd1 vssd1 vccd1 vccd1 _11574_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10597__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10597__B2 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10525_ _10525_/A _10525_/B vssd1 vssd1 vccd1 vccd1 _10526_/B sky130_fd_sc_hd__nand2_2
X_13313_ _13324_/CLK _13313_/D vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _10608_/B _10456_/B vssd1 vssd1 vccd1 vccd1 _10458_/C sky130_fd_sc_hd__nand2_1
X_13244_ _13341_/CLK _13244_/D vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13175_/A _13175_/B vssd1 vssd1 vccd1 vccd1 _13175_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12126_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__nor2_1
X_10387_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12057_ _12056_/B _12057_/B vssd1 vssd1 vccd1 vccd1 _12058_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11008_ _10929_/X _11041_/C _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06740__A3 _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ hold230/X _13095_/B2 _13158_/A2 hold261/X vssd1 vssd1 vccd1 vccd1 hold262/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__B _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__xnor2_2
X_07101_ _07101_/A _07101_/B vssd1 vssd1 vccd1 vccd1 _07101_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07032_ fanout67/X _08551_/B2 fanout55/X _06973_/A vssd1 vssd1 vccd1 vccd1 _07033_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08290__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11537__B1 _11512_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10325__A _11296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08953__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ reg1_val[30] _08983_/B vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08953__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _07932_/X _07934_/B vssd1 vssd1 vccd1 vccd1 _08705_/A sky130_fd_sc_hd__nand2b_4
X_07865_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__nand2_1
X_09604_ _09540_/A _09540_/B _09538_/X vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10060__A _10234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _10280_/A _06814_/Y _06815_/X vssd1 vssd1 vccd1 vccd1 _06816_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07796_ _07794_/A _07794_/B _07795_/Y vssd1 vssd1 vccd1 vccd1 _07860_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11068__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06747_ reg1_val[9] _07217_/A vssd1 vssd1 vccd1 vccd1 _06747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08469__B1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06678_ reg2_val[21] _06712_/B _06600_/Y _06677_/Y vssd1 vssd1 vccd1 vccd1 _06964_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_09466_ _09466_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08465__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08417_ _08429_/A _08429_/B _08403_/Y vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__o21a_1
X_09397_ _09246_/X _09396_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09397_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08184__B _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08348_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08641__B1 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07444__B2 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07444__A1 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _08619_/B2 _10067_/A1 _08926_/B1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08280_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _11290_/A _11290_/B vssd1 vssd1 vccd1 vccd1 _11291_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ _10310_/A _10310_/B _10310_/C vssd1 vssd1 vccd1 vccd1 _10313_/B sky130_fd_sc_hd__or3_1
XFILLER_0_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10241_ _10241_/A _10372_/B _10241_/C vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__and3_1
X_10172_ curr_PC[6] _10172_/B vssd1 vssd1 vccd1 vccd1 _10438_/C sky130_fd_sc_hd__and2_1
XFILLER_0_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12450__A _12627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 _09238_/X vssd1 vssd1 vccd1 vccd1 _12433_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout172 _07066_/Y vssd1 vssd1 vccd1 vccd1 _10234_/A sky130_fd_sc_hd__buf_12
Xfanout161 _06942_/Y vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__buf_4
Xfanout150 _07011_/Y vssd1 vssd1 vccd1 vccd1 _08649_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout194 _09941_/A vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__buf_12
XFILLER_0_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ hold53/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ reg1_val[26] _12773_/A vssd1 vssd1 vccd1 vccd1 _12744_/X sky130_fd_sc_hd__and2_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10019__B1 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07683__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ _09886_/B _12394_/A1 _11626_/S vssd1 vssd1 vccd1 vccd1 _11626_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09424__A2 _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11557_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__xnor2_1
X_10508_ _10507_/A _10507_/B _10507_/C vssd1 vssd1 vccd1 vccd1 _10509_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__06789__A3 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _11486_/A _11486_/B _11489_/B vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13227_ hold149/X _13227_/B vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__nand2_1
X_10439_ curr_PC[7] _10438_/C curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ hold320/X _13158_/A2 _13157_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 _13159_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12109_ hold314/A _12109_/B vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__or2_1
XANTENNA__12360__A fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13089_ hold265/X _13088_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__mux2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07650_ _07650_/A _07650_/B vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__xnor2_4
X_06601_ instruction[39] _06657_/B vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__and2_4
XANTENNA__12247__A1 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__A3 _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07581_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12798__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09320_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09112__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A1 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _09251_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_118_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09178_/X _09181_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__A2 _11258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08623__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08133_ _10468_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout218_A _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _08049_/B _08011_/C _08011_/B vssd1 vssd1 vccd1 vccd1 _08067_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07016_/A _07016_/B vssd1 vssd1 vccd1 vccd1 _07015_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08926__B2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__B2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _08967_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _09062_/B sky130_fd_sc_hd__or2_1
X_08897_ _08897_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__nor2_1
X_07917_ _07941_/A _07941_/B _07885_/Y vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10497__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07848_ _07918_/A _07918_/B _07828_/Y vssd1 vssd1 vccd1 vccd1 _07856_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06627__A_N _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ _09324_/A _11155_/A _09330_/B _09328_/X vssd1 vssd1 vccd1 vccd1 _09520_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__09103__A1 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__B2 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _08553_/B1 _08096_/B fanout24/X _09468_/B2 vssd1 vssd1 vccd1 vccd1 _07780_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10790_ _12171_/A _10789_/X _10786_/X vssd1 vssd1 vccd1 vccd1 _10790_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout33_A _07181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11461__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09449_ _09622_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12460_/A _12460_/B _12460_/C vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11411_/A _11411_/B _11411_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12391_ hold287/A _12391_/B vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _11879_/A2 _11524_/C hold320/A vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07539__A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12961__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__B2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273_ _07180_/X fanout7/X _11272_/Y vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ _13219_/A hold264/X vssd1 vssd1 vccd1 vccd1 _13304_/D sky130_fd_sc_hd__and2_1
X_10224_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__nand2b_1
X_10155_ hold232/A _10427_/A2 _10289_/B _10154_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _10155_/Y sky130_fd_sc_hd__a311oi_1
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__and2_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_10988_ _10989_/A _10989_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09645__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ reg1_val[22] _12773_/A vssd1 vssd1 vccd1 vccd1 _12728_/B sky130_fd_sc_hd__or2_1
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _12656_/Y _12658_/B vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ instruction[7] _11609_/B vssd1 vssd1 vccd1 vccd1 _11611_/C sky130_fd_sc_hd__or2_1
XFILLER_0_53_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12589_ _12589_/A vssd1 vssd1 vccd1 vccd1 _12598_/C sky130_fd_sc_hd__inv_2
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09648__B _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12165__B1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09581__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08820_ _08820_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _08751_/A _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__and3_1
X_07702_ _08926_/B1 _08274_/B fanout74/X _08521_/A2 vssd1 vssd1 vccd1 vccd1 _07703_/B
+ sky130_fd_sc_hd__o22a_2
X_08682_ _08682_/A _08682_/B vssd1 vssd1 vccd1 vccd1 _08758_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07895__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _07634_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07895__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07564_ _07565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__and2_1
X_09303_ _09305_/B _09305_/C _09670_/A vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__a21oi_1
X_07495_ _10067_/A1 _08274_/B fanout74/X _09114_/B1 vssd1 vssd1 vccd1 vccd1 _07496_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ instruction[4] instruction[6] instruction[5] instruction[3] vssd1 vssd1 vccd1
+ vccd1 _11966_/B sky130_fd_sc_hd__and4bb_4
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ reg1_val[7] reg1_val[24] _09180_/S vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__mux2_1
X_08116_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09096_ _09097_/A _09097_/B vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08047_ _07959_/A _07959_/C _07959_/B vssd1 vssd1 vccd1 vccd1 _08048_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13096__A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__A2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10182__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _10267_/A _09707_/X _10319_/A _09997_/X vssd1 vssd1 vccd1 vccd1 _09998_/X
+ sky130_fd_sc_hd__o31a_1
X_08949_ fanout64/X _08590_/B _09648_/A fanout58/X vssd1 vssd1 vccd1 vccd1 _08950_/B
+ sky130_fd_sc_hd__o22a_1
X_11960_ hold199/A _11960_/B vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__or2_1
X_10911_ _12171_/A _10904_/Y _10908_/X _10910_/Y vssd1 vssd1 vccd1 vccd1 _10911_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07335__B1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11891_ curr_PC[22] _11891_/B vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10659__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__B2 _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A1 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10842_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10773_ _10774_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10773_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08835__B1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _12673_/B _12513_/B vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07102__A3 _12717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _12622_/B _12443_/B vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _12330_/A _12330_/B _12374_/C _12374_/D vssd1 vssd1 vccd1 vccd1 _12374_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _11504_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11256_ _12490_/S _11448_/C vssd1 vssd1 vccd1 vccd1 _11256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06901__A _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12622__B _12622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__A1 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _11060_/A _11060_/B _11057_/A vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__a21bo_1
X_10207_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11370__B2 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _12420_/A _10137_/B _10137_/C vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__a21o_1
X_10069_ _10326_/A _08873_/X _08988_/Y _10213_/A vssd1 vssd1 vccd1 vccd1 _10070_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08118__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07877__A1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__B2 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07629__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__B2 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ _10469_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07282_/B sky130_fd_sc_hd__or2_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07179__A _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__B2 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__A1 _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _09920_/B _09921_/B vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07907__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09003__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__and2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__xnor2_1
X_08803_ _08803_/A _08803_/B vssd1 vssd1 vccd1 vccd1 _08803_/X sky130_fd_sc_hd__or2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout285_A _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06995_ _06991_/A _06991_/B _09301_/A vssd1 vssd1 vccd1 vccd1 _06995_/X sky130_fd_sc_hd__mux2_2
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _10896_/B sky130_fd_sc_hd__xnor2_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11113__A1 _10653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _08666_/B _08716_/A _08666_/A vssd1 vssd1 vccd1 vccd1 _08718_/B sky130_fd_sc_hd__o21ba_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08596_ _08588_/A _08588_/B _08588_/C _08595_/X vssd1 vssd1 vccd1 vccd1 _08669_/A
+ sky130_fd_sc_hd__a31o_2
X_07616_ _09827_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07618_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ _07547_/A _07547_/B vssd1 vssd1 vccd1 vccd1 _07550_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07551_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _09217_/A vssd1 vssd1 vccd1 vccd1 _09217_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _09235_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09148_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ _09787_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11110_/A _11217_/A vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06815__A_N _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12090_ _11936_/Y _12215_/A _12089_/Y vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11339__A _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11041_/A _11041_/B _11041_/C vssd1 vssd1 vccd1 vccd1 _11809_/B sky130_fd_sc_hd__nand3_2
XANTENNA__09545__B2 _09370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__B _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ _13144_/A hold226/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__and2_1
XFILLER_0_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11943_ _11895_/X _12020_/D _11942_/Y vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__o21a_1
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10825_ _10826_/B _10826_/A vssd1 vssd1 vccd1 vccd1 _10825_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10756_ _10757_/B _10757_/A vssd1 vssd1 vccd1 vccd1 _10756_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09481__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10687_ curr_PC[9] _10686_/C curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10688_/C sky130_fd_sc_hd__a21oi_1
X_12426_ hold324/A _12391_/X _12349_/A vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11013__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__B2 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09784__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12357_ _08971_/A _11446_/B _12333_/X _12356_/X _11975_/A vssd1 vssd1 vccd1 vccd1
+ dest_val[29] sky130_fd_sc_hd__o221a_4
XANTENNA__09784__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08830__B _08831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11308_ _11204_/A _11203_/Y _11201_/X vssd1 vssd1 vccd1 vccd1 _11309_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06631__A _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12288_ _10315_/A _08808_/A _08808_/B _09232_/Y _12287_/Y vssd1 vssd1 vccd1 vccd1
+ _12304_/B sky130_fd_sc_hd__o311a_1
X_11239_ hold234/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__or2_1
X_06780_ _06780_/A _06780_/B vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07462__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08450_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08490_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08381_ _08410_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08382_/B sky130_fd_sc_hd__nand2_1
X_07401_ _09827_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07332_ _09827_/A _07332_/B vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08293__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__A1 _11645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07263_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12359__B1 _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _07113_/A _06954_/B _07195_/B vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _09795_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout200_A _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _09904_/A _09904_/B vssd1 vssd1 vccd1 vccd1 _10038_/A sky130_fd_sc_hd__nand2_1
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09836_/B sky130_fd_sc_hd__xnor2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06978_ _06978_/A _06978_/B vssd1 vssd1 vccd1 vccd1 _06978_/X sky130_fd_sc_hd__xor2_4
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09767_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11637__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__A1 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09697_ _09697_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__xnor2_2
X_08717_ _10140_/B _10140_/C vssd1 vssd1 vccd1 vccd1 _10276_/B sky130_fd_sc_hd__and2_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08648_ _08648_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _08653_/A sky130_fd_sc_hd__xnor2_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08579_ _08577_/Y _08597_/B _08564_/Y vssd1 vssd1 vccd1 vccd1 _08584_/A sky130_fd_sc_hd__o21ai_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _11592_/A _11592_/B _11592_/C vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10610_ _10610_/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12062__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _11776_/A _10541_/B _10541_/C vssd1 vssd1 vccd1 vccd1 _10541_/X sky130_fd_sc_hd__or3_1
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _13364_/CLK _13260_/D vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08018__A1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12213_/A vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__inv_2
X_10472_ _10472_/A _10472_/B vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08569__A2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08018__B2 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ hold289/X _13209_/A2 _13190_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold290/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12142_ _07301_/Y _08873_/X _08988_/Y _07031_/X vssd1 vssd1 vccd1 vccd1 _12202_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11069__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _12073_/A _12073_/B _12073_/C vssd1 vssd1 vccd1 vccd1 _12074_/B sky130_fd_sc_hd__nor3_1
XANTENNA__09518__A1 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ hold220/A _11024_/B vssd1 vssd1 vccd1 vccd1 _11134_/B sky130_fd_sc_hd__or2_1
XANTENNA__10701__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13078__B2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12286__C1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ hold207/X _13095_/B2 _13158_/A2 hold220/X vssd1 vssd1 vccd1 vccd1 hold221/A
+ sky130_fd_sc_hd__a22o_1
X_11926_ _11926_/A _11926_/B vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13297_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ _11857_/A vssd1 vssd1 vccd1 vccd1 _11857_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ _11958_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10808_ _12490_/S _10808_/B vssd1 vssd1 vccd1 vccd1 _10808_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11261__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ _10862_/B _10739_/B vssd1 vssd1 vccd1 vccd1 _10742_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09002__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12409_ _12409_/A _12409_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _08045_/B _07950_/B vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06901_ _12781_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _06901_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07881_ _07881_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06832_ _11228_/A _06830_/Y _06831_/X vssd1 vssd1 vccd1 vccd1 _06832_/Y sky130_fd_sc_hd__o21bai_1
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08288__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__A1 _07243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ _06763_/A vssd1 vssd1 vccd1 vccd1 _06765_/A sky130_fd_sc_hd__inv_2
X_09551_ _12339_/A1 _09758_/A _10310_/C _11889_/A1 vssd1 vssd1 vccd1 vccd1 _09552_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10827__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08502_ _08520_/B vssd1 vssd1 vccd1 vccd1 _08502_/Y sky130_fd_sc_hd__inv_2
X_06694_ _06692_/Y _06707_/B1 _06712_/B reg2_val[18] vssd1 vssd1 vccd1 vccd1 _07068_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_09482_ _10469_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09483_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08496__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08619_/B2 _08551_/A2 _08551_/B1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08434_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06660__A_N _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09445__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _09468_/B2 _10227_/B1 _10463_/A1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 _08365_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12257__B _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07315_ _07372_/A _07372_/B vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ _08291_/A _08291_/B _08294_/Y vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ reg1_val[14] _07246_/B vssd1 vssd1 vccd1 vccd1 _07248_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11555__A1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ _07213_/A _07113_/A _06954_/B _06958_/C _07299_/B vssd1 vssd1 vccd1 vccd1
+ _07179_/B sky130_fd_sc_hd__o41a_4
XANTENNA__09748__A1 _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09818_ _11155_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07814__B _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A _06994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _06785_/X _09595_/B _11966_/B _06787_/B _09748_/X vssd1 vssd1 vccd1 vccd1
+ _09749_/X sky130_fd_sc_hd__a221o_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12764_/B _12760_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__nor2_8
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11711_ _09886_/B _12394_/A1 _11711_/S vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ reg1_val[14] _12691_/B vssd1 vssd1 vccd1 vccd1 _12692_/B sky130_fd_sc_hd__or2_1
X_11642_ _11641_/B _11642_/B vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__and2b_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09436__B1 _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11071__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__B2 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11573_ _11482_/A _11482_/B _11481_/A vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10597__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13312_ _13324_/CLK _13312_/D vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10525_/B sky130_fd_sc_hd__or2_1
XFILLER_0_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10455_ _10454_/B _10455_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand2b_1
X_13243_ _13341_/CLK _13243_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11546__B2 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13187_/A hold276/X vssd1 vssd1 vccd1 vccd1 _13357_/D sky130_fd_sc_hd__and2_1
XANTENNA__11546__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07277__A _10469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__xor2_1
X_12125_ _06908_/C _12121_/X _12124_/X vssd1 vssd1 vccd1 vccd1 dest_val[25] sky130_fd_sc_hd__o21ai_4
XFILLER_0_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12056_ _12057_/B _12056_/B vssd1 vssd1 vccd1 vccd1 _12058_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09492__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _11217_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11041_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _12978_/A hold231/X vssd1 vssd1 vccd1 vccd1 _13277_/D sky130_fd_sc_hd__and2_1
XFILLER_0_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08836__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _11910_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__or2_1
XFILLER_0_90_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12889_ hold273/X hold3/X vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11262__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _07101_/A _07101_/B vssd1 vssd1 vccd1 vccd1 _07100_/X sky130_fd_sc_hd__and2_1
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08080_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08080_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12805__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07299_/B _07025_/X _08971_/D _07029_/Y vssd1 vssd1 vccd1 vccd1 _07031_/X
+ sky130_fd_sc_hd__a31o_4
XANTENNA__11537__B2 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06803__B _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08402__A1 _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08953__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07933_ _07932_/A _07932_/B _07932_/C vssd1 vssd1 vccd1 vccd1 _07934_/B sky130_fd_sc_hd__a21o_1
X_07864_ _07864_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07928_/B sky130_fd_sc_hd__xnor2_4
X_06815_ _07202_/A reg1_val[7] vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__and2b_1
X_09603_ _09758_/A _10310_/C _12420_/A vssd1 vssd1 vccd1 vccd1 _09603_/Y sky130_fd_sc_hd__o21ai_1
X_07795_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07795_/Y sky130_fd_sc_hd__nand2b_1
X_06746_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07218_/A sky130_fd_sc_hd__inv_2
X_09534_ _09534_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08469__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06677_ _06706_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _06677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _09466_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11172__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08416_ _08416_/A _08416_/B vssd1 vssd1 vccd1 vccd1 _08429_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09396_ _09193_/X _09195_/X _09396_/S vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11225__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10579__A2 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08683_/A _08683_/B _08683_/C vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11900__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12973__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__B2 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__A1 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07444__A2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _08566_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__xnor2_2
X_07229_ reg1_val[11] _07229_/B _07229_/C vssd1 vssd1 vccd1 vccd1 _07230_/B sky130_fd_sc_hd__and3_1
XFILLER_0_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10240_ _10372_/A _10239_/C _10086_/A vssd1 vssd1 vccd1 vccd1 _10241_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__07097__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _09148_/Y _10137_/Y _10138_/X _10170_/X vssd1 vssd1 vccd1 vccd1 _10171_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout140 _09467_/A vssd1 vssd1 vccd1 vccd1 _08591_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout173 _07066_/Y vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__clkbuf_4
Xfanout162 _06942_/Y vssd1 vssd1 vccd1 vccd1 _12339_/A1 sky130_fd_sc_hd__buf_2
Xfanout151 _07011_/Y vssd1 vssd1 vccd1 vccd1 _09297_/B2 sky130_fd_sc_hd__buf_4
Xfanout184 _09238_/X vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout195 _06984_/Y vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__buf_12
XANTENNA__07904__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _07255_/Y _12842_/A2 hold57/X _13144_/A vssd1 vssd1 vccd1 vccd1 hold58/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ _12743_/A _12747_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
XANTENNA__11082__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12682_/A _12674_/B vssd1 vssd1 vccd1 vccd1 _12676_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07683__A2 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ hold275/A _11879_/A2 _11708_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11625_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09424__A3 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _11900_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11557_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09487__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _10507_/A _10507_/B _10507_/C vssd1 vssd1 vccd1 vccd1 _10509_/B sky130_fd_sc_hd__or3_1
XFILLER_0_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11487_ _11379_/A _11379_/B _11376_/A vssd1 vssd1 vccd1 vccd1 _11489_/B sky130_fd_sc_hd__a21oi_2
X_13226_ _13226_/A hold175/X vssd1 vssd1 vccd1 vccd1 _13369_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ curr_PC[7] curr_PC[8] _10438_/C vssd1 vssd1 vccd1 vccd1 _10686_/C sky130_fd_sc_hd__and3_2
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13157_ hold297/X _13156_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
X_10369_ _10370_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _10369_/Y sky130_fd_sc_hd__nor2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _11238_/S _12106_/Y _12107_/X vssd1 vssd1 vccd1 vccd1 _12108_/Y sky130_fd_sc_hd__o21ai_1
X_13088_ _13088_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _13088_/Y sky130_fd_sc_hd__xnor2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ hold228/A _12178_/A2 _12112_/B _12038_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12039_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09896__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06600_ _06908_/A _06600_/B vssd1 vssd1 vccd1 vccd1 _06600_/Y sky130_fd_sc_hd__nand2_4
X_07580_ _12193_/A _07346_/B _11813_/A vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__08566__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__B1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07470__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A2 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _10902_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _09251_/B sky130_fd_sc_hd__or2_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08201_ _08204_/A _08204_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__or2_1
XFILLER_0_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09179_/X _09180_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11720__A _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__A3 _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08132_ _08553_/A2 _08400_/B fanout82/X _08553_/B1 vssd1 vssd1 vccd1 vccd1 _08133_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _08063_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_113_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07014_ _06994_/A _06967_/A _06966_/C _07074_/B vssd1 vssd1 vccd1 vccd1 _07016_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA_fanout113_A _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10194__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A2 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _11168_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11167__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__xor2_1
X_08896_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10497__B2 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A1 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _07847_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__xnor2_2
X_07778_ _07784_/B _07784_/A vssd1 vssd1 vccd1 vccd1 _07778_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08476__A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06729_ _06908_/A _06801_/B1 _12685_/B _06728_/X vssd1 vssd1 vccd1 vccd1 _07175_/A
+ sky130_fd_sc_hd__a31o_4
X_09517_ _09517_/A _09517_/B vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09103__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _09447_/B _09448_/B vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout26_A fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _09158_/X _09161_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09379_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _11411_/A _11411_/B _11411_/C vssd1 vssd1 vccd1 vccd1 _11410_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _12390_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ hold331/A _11341_/B vssd1 vssd1 vccd1 vccd1 _11524_/C sky130_fd_sc_hd__or2_1
XFILLER_0_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08090__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__B _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ _07172_/B fanout7/X _10081_/A vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13011_ hold253/X _06564_/A _13222_/A2 hold263/X vssd1 vssd1 vccd1 vccd1 hold264/A
+ sky130_fd_sc_hd__a22o_1
X_10223_ _12193_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10225_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10427_/A2 _10289_/B hold232/A vssd1 vssd1 vccd1 vccd1 _10154_/Y sky130_fd_sc_hd__a21oi_1
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__or2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07290__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _10989_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ reg1_val[22] _12773_/A vssd1 vssd1 vccd1 vccd1 _12728_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12657_ reg1_val[8] _12657_/B vssd1 vssd1 vccd1 vccd1 _12658_/B sky130_fd_sc_hd__nand2_1
X_11608_ _06697_/Y _11515_/B _11531_/S vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__a21oi_1
X_12588_ _12588_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__C _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ curr_PC[18] _11539_/B vssd1 vssd1 vccd1 vccd1 _11718_/C sky130_fd_sc_hd__and2_2
Xmax_cap115 _07179_/X vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__buf_6
XFILLER_0_13_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09945__A _10613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ hold301/X _13209_/A2 _13208_/X _12781_/A vssd1 vssd1 vccd1 vccd1 _13210_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__S _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _08760_/A sky130_fd_sc_hd__nor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ _07701_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__xnor2_4
X_08681_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08681_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _11168_/A _07632_/B vssd1 vssd1 vccd1 vccd1 _07634_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07895__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _09301_/B _09301_/C _09301_/A vssd1 vssd1 vccd1 vccd1 _09305_/C sky130_fd_sc_hd__a21o_1
X_07563_ _09630_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07494_ _08445_/A _07494_/B vssd1 vssd1 vccd1 vccd1 _07500_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09233_ _09233_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _11946_/A sky130_fd_sc_hd__or2_4
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13343_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ reg1_val[6] reg1_val[25] _09180_/S vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09095_ _09095_/A _09095_/B vssd1 vssd1 vccd1 vccd1 _09097_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08046_ _08046_/A _08046_/B vssd1 vssd1 vccd1 vccd1 _08048_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07032__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ _09703_/X _09855_/X _09856_/X vssd1 vssd1 vccd1 vccd1 _09997_/X sky130_fd_sc_hd__a21o_1
X_08948_ _10230_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _08952_/A sky130_fd_sc_hd__xnor2_1
X_08879_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08879_/X sky130_fd_sc_hd__or2_1
X_10910_ _12171_/A _10910_/B vssd1 vssd1 vccd1 vccd1 _10910_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07335__A1 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__B2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _06994_/A _11446_/B _06941_/X _11889_/X vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06719__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _11001_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10810_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08835__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ reg1_val[11] curr_PC[11] _12525_/S vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11360__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12456__A _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12442_ _12622_/B _12443_/B vssd1 vssd1 vccd1 vccd1 _12453_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12395__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11324_ _10406_/A _10890_/X _11322_/X _11323_/X vssd1 vssd1 vccd1 vccd1 _11325_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ curr_PC[15] _11255_/B vssd1 vssd1 vccd1 vccd1 _11448_/C sky130_fd_sc_hd__and2_1
XANTENNA__10704__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__B1 _09240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07023__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _11186_/A _11186_/B vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11370__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _12420_/A _10137_/B _10137_/C vssd1 vssd1 vccd1 vccd1 _10137_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _12131_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08523__B1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07877__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07629__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _12709_/A _12709_/B vssd1 vssd1 vccd1 vccd1 _12716_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__A _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12813__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _09921_/B _09920_/B vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09003__A1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07195__A _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09003__B2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__B1 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ _06994_/A _06994_/B vssd1 vssd1 vccd1 vccd1 _06994_/Y sky130_fd_sc_hd__xnor2_4
X_09782_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09782_/X sky130_fd_sc_hd__and2b_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _07801_/Y _08696_/B _08698_/Y vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__a21o_1
X_08733_ _08673_/A _08726_/A _08726_/B _08726_/C _08732_/X vssd1 vssd1 vccd1 vccd1
+ _08734_/B sky130_fd_sc_hd__a41o_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout278_A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08664_ _08637_/X _08714_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__a21o_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08595_/A _08595_/B _08602_/A _08595_/D vssd1 vssd1 vccd1 vccd1 _08595_/X
+ sky130_fd_sc_hd__and4_1
X_07615_ _07814_/B _07201_/X _07264_/X fanout45/X vssd1 vssd1 vccd1 vccd1 _07616_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07546_ _07546_/A _07546_/B vssd1 vssd1 vccd1 vccd1 _07553_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11821__B1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _09184_/X _09215_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__mux2_1
X_07477_ _07477_/A _07477_/B _07520_/A vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ _12339_/A1 _10310_/A _10310_/B vssd1 vssd1 vccd1 vccd1 _09147_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ fanout52/X fanout85/X _10466_/A fanout50/X vssd1 vssd1 vccd1 vccd1 _09079_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _08624_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout93_A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__A2 _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _12525_/S _11037_/X _11038_/X _11039_/Y vssd1 vssd1 vccd1 vccd1 dest_val[13]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10560__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ hold237/A _13143_/B2 _13186_/A2 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12301__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__B1 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _11895_/X _12020_/D _09149_/X vssd1 vssd1 vccd1 vccd1 _11942_/Y sky130_fd_sc_hd__a21oi_1
X_11873_ _11785_/B _11787_/B _11785_/A vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__a21bo_1
X_10824_ _10824_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10826_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ _10755_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10757_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11812__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ curr_PC[9] curr_PC[10] _10686_/C vssd1 vssd1 vccd1 vccd1 _10926_/C sky130_fd_sc_hd__and3_1
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ hold162/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12425_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08036__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12356_/A _12356_/B _12356_/C _12344_/X vssd1 vssd1 vccd1 vccd1 _12356_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__09784__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09495__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__A1 _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07244__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11307_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08992__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06631__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _12280_/A _08808_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _12287_/Y sky130_fd_sc_hd__o21ai_1
X_11238_ _11234_/Y _11237_/X _11238_/S vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__mux2_1
X_11169_ _11169_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07743__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08380_ _08380_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__xnor2_1
X_07400_ _07814_/B _09815_/A fanout45/X _09675_/A vssd1 vssd1 vccd1 vccd1 _07401_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07331_ _09928_/A fanout45/X _08551_/B1 _07814_/B vssd1 vssd1 vccd1 vccd1 _07332_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10082__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _11361_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__xnor2_1
X_07193_ _07193_/A _07193_/B vssd1 vssd1 vccd1 vccd1 _07193_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09001_ _10859_/A fanout24/X _10966_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _09002_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11031__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13020__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _12053_/A1 _09901_/Y _09902_/X _09900_/X vssd1 vssd1 vccd1 vccd1 dest_val[4]
+ sky130_fd_sc_hd__a31o_4
X_09834_ _09954_/A _09834_/B _09835_/B vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11175__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06977_ _06978_/A _06978_/B vssd1 vssd1 vccd1 vccd1 _06977_/Y sky130_fd_sc_hd__xnor2_2
X_09765_ _07539_/B _10222_/A2 _10712_/A fanout37/X vssd1 vssd1 vccd1 vccd1 _09766_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12834__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12295__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _08716_/A _08716_/B vssd1 vssd1 vccd1 vccd1 _10140_/C sky130_fd_sc_hd__xor2_1
X_09696_ _09534_/A _09534_/B _09532_/X vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__a21oi_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ _08605_/A _07128_/Y _07153_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _08648_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__xnor2_2
X_07529_ _09630_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07531_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ _11776_/A _10541_/B _10541_/C vssd1 vssd1 vccd1 vccd1 _10540_/Y sky130_fd_sc_hd__o21ai_1
X_10471_ _10471_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08018__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13011__A2 _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _12212_/A _12212_/B _12212_/C vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ hold316/A _13189_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__mux2_1
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08974__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ _12073_/A _12073_/B _12073_/C vssd1 vssd1 vccd1 vccd1 _12074_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09518__A2 _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _11020_/Y _11022_/X _11958_/A vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07563__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__A2 _13227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ _12978_/A hold208/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__and2_1
XFILLER_0_63_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11925_ _11926_/A _11926_/B vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11856_/A _12016_/A vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__nand2_1
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06626__B _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ curr_PC[11] _10926_/C vssd1 vssd1 vccd1 vccd1 _10808_/B sky130_fd_sc_hd__and2_1
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11261__B2 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10738_ _10738_/A _10738_/B vssd1 vssd1 vccd1 vccd1 _10739_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07465__B1 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _12220_/B _12406_/Y _12407_/Y _12368_/B vssd1 vssd1 vccd1 vccd1 _12409_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_70_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10669_ _10009_/Y _10668_/Y _11237_/S vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09757__A2 _09753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ _12339_/A1 _08808_/Y _08809_/A vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06900_ _06767_/A _06593_/X _09240_/B instruction[4] _06897_/Y vssd1 vssd1 vccd1
+ vccd1 _12781_/B sky130_fd_sc_hd__a221o_1
XANTENNA__09164__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__nor2_1
X_06831_ _07243_/A _11231_/A vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06762_ reg1_val[6] _07264_/A vssd1 vssd1 vccd1 vccd1 _06763_/A sky130_fd_sc_hd__or2_1
X_09550_ _12339_/A1 _09758_/A _10310_/C vssd1 vssd1 vccd1 vccd1 _09552_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10827__B2 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__A1 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ fanout67/X _10233_/B2 _10233_/A1 fanout64/X vssd1 vssd1 vccd1 vccd1 _09482_/B
+ sky130_fd_sc_hd__o22a_1
X_08501_ _08624_/A _08501_/B vssd1 vssd1 vccd1 vccd1 _08520_/B sky130_fd_sc_hd__xnor2_2
X_06693_ reg2_val[18] _06712_/B _06707_/B1 _06692_/Y vssd1 vssd1 vccd1 vccd1 _07067_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ _08556_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08438_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08496__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09445__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A1 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _08413_/A _08413_/B _08358_/X vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11252__A1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07314_ _10234_/A _07314_/B vssd1 vssd1 vccd1 vccd1 _07372_/B sky130_fd_sc_hd__xnor2_1
X_08294_ _08338_/B _08338_/A vssd1 vssd1 vccd1 vccd1 _08294_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ _09787_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07259_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__B1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _07113_/A _06954_/B _06958_/C _07299_/B vssd1 vssd1 vccd1 vccd1 _07213_/B
+ sky130_fd_sc_hd__o31a_4
XANTENNA__09748__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11555__A2 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ _07264_/X fanout9/A fanout5/X _09928_/A vssd1 vssd1 vccd1 vccd1 _09818_/B
+ sky130_fd_sc_hd__o22a_1
X_09748_ _07145_/A _06940_/B _09239_/Y _09747_/X vssd1 vssd1 vccd1 vccd1 _09748_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout56_A _07015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ hold302/A _11879_/A2 _11790_/B _12175_/C1 vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07144__C1 _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _09680_/A _09680_/B vssd1 vssd1 vccd1 vccd1 _09679_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ reg1_val[14] _12691_/B vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ _11642_/B _11641_/B vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__and2b_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _11483_/A _11483_/B _11471_/Y vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__10046__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10523_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13324_/CLK hold159/X vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12464__A _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10454_ _10455_/B _10454_/B vssd1 vssd1 vccd1 vccd1 _10608_/B sky130_fd_sc_hd__nand2b_1
X_13242_ _13341_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11546__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ hold275/X _13209_/A2 _13172_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold276/A
+ sky130_fd_sc_hd__a22o_1
X_10385_ _10383_/X _10385_/B vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08947__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _12504_/S _12124_/B _12124_/C vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__or3_1
XANTENNA__10712__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _12404_/B _12055_/B vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__xnor2_1
X_11006_ _10000_/B _10534_/Y _11004_/Y _11005_/Y vssd1 vssd1 vccd1 vccd1 _11007_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__12259__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ hold325/X _13095_/B2 _13158_/A2 hold230/X vssd1 vssd1 vccd1 vccd1 hold231/A
+ sky130_fd_sc_hd__a22o_1
X_11908_ _12001_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06637__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12888_ _13338_/Q hold165/X vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11839_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11841_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10037__A2 _10033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07030_ _07299_/B _07025_/X _08971_/D _07029_/Y vssd1 vssd1 vccd1 vccd1 _07030_/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__09159__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10606__B _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__xnor2_2
X_07932_ _07932_/A _07932_/B _07932_/C vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__and3_1
X_07863_ _07863_/A _07863_/B vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__nor2_2
X_06814_ _10143_/A _06812_/X _06813_/Y vssd1 vssd1 vccd1 vccd1 _06814_/Y sky130_fd_sc_hd__o21ai_1
X_09602_ _12053_/A1 _09438_/Y _09439_/X _09601_/X vssd1 vssd1 vccd1 vccd1 dest_val[2]
+ sky130_fd_sc_hd__a31o_4
X_09533_ _09533_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__xor2_2
X_07794_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout260_A _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06745_ _06799_/A _06801_/B1 _12666_/B _06744_/X vssd1 vssd1 vccd1 vccd1 _07217_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__08469__A2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06676_ instruction[0] instruction[1] instruction[2] instruction[31] pred_val vssd1
+ vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__o311a_4
XANTENNA__11473__A1 _11837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _09464_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09395_ _09393_/X _09394_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__mux2_1
X_08415_ _08414_/A _08460_/A _08414_/B _08411_/X vssd1 vssd1 vccd1 vccd1 _08429_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11225__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08683_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07429__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__B1 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__A2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ _06875_/A fanout75/X fanout71/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08278_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ _07229_/B _07229_/C reg1_val[11] vssd1 vssd1 vccd1 vccd1 _07230_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07097__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ _07142_/A _07142_/B _07357_/A vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_30_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _12029_/A _10139_/Y _10140_/X _10169_/X vssd1 vssd1 vccd1 vccd1 _10170_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07601__B1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _07100_/X vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__buf_4
Xfanout163 _12178_/A2 vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__buf_4
Xfanout174 _06949_/Y vssd1 vssd1 vccd1 vccd1 _07074_/B sky130_fd_sc_hd__clkbuf_8
Xfanout152 _06995_/X vssd1 vssd1 vccd1 vccd1 _08619_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout141 _09675_/A vssd1 vssd1 vccd1 vccd1 _09468_/B2 sky130_fd_sc_hd__buf_6
XANTENNA__11161__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _06925_/X vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__clkbuf_8
Xfanout185 _09235_/X vssd1 vssd1 vccd1 vccd1 _12394_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__07904__B2 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A1 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ hold56/X _12841_/B vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09657__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ reg1_val[25] _12773_/A vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__xnor2_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12673_ reg1_val[11] _12673_/B vssd1 vssd1 vccd1 vccd1 _12674_/B sky130_fd_sc_hd__or2_1
X_11624_ _11879_/A2 _11708_/B hold275/A vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ fanout44/X _12257_/A fanout13/X fanout46/X vssd1 vssd1 vccd1 vccd1 _11556_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__nand2_1
X_10506_ _10506_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10507_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07288__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07840__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13225_ hold324/X _12781_/A _13224_/Y _12780_/B hold174/X vssd1 vssd1 vccd1 vccd1
+ hold175/A sky130_fd_sc_hd__a32o_1
X_10437_ _10408_/X _10411_/Y _10415_/X _10436_/X _12053_/A1 vssd1 vssd1 vccd1 vccd1
+ _10437_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07199__A2 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _13156_/A _13156_/B vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10368_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__xor2_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12641__B _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ _12171_/A _10146_/X _12107_/B1 vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__o21a_1
X_13087_ _13087_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__nand2_1
X_10299_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__nor2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12038_ _12178_/A2 _12112_/B hold228/A vssd1 vssd1 vccd1 vccd1 _12038_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09896__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11455__A1 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08204_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09678__A _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _11231_/A reg1_val[16] _09180_/S vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10415__C1 _11612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__A2 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _08320_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08134_/B sky130_fd_sc_hd__xnor2_1
X_08062_ _08052_/A _08052_/C _08052_/B vssd1 vssd1 vccd1 vccd1 _08063_/B sky130_fd_sc_hd__o21ai_1
X_07013_ _06975_/A _06974_/X _06975_/Y _06967_/Y vssd1 vssd1 vccd1 vccd1 _07013_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10718__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10194__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08964_ fanout98/X fanout77/X fanout73/X _11296_/A vssd1 vssd1 vccd1 vccd1 _08965_/B
+ sky130_fd_sc_hd__o22a_1
X_07915_ _07953_/A _07953_/B _07913_/B _07914_/Y vssd1 vssd1 vccd1 vccd1 _07941_/A
+ sky130_fd_sc_hd__o31ai_2
X_08895_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__and2_1
XANTENNA__10497__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__B1 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _07921_/A _07921_/B _07839_/X vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__a21o_1
X_07777_ _07810_/A _07810_/B _07773_/Y vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06728_ reg2_val[12] _06767_/A vssd1 vssd1 vccd1 vccd1 _06728_/X sky130_fd_sc_hd__and2_1
X_09516_ _09630_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09517_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08476__B _08476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09448_/B _09447_/B vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__and2b_1
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06659_ reg2_val[23] _06767_/A _06600_/Y _06658_/Y vssd1 vssd1 vccd1 vccd1 _07016_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _09154_/X _09157_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout19_A _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08075__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _08380_/A _08380_/B _08325_/X vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__o21a_2
X_11340_ _12171_/A _11338_/Y _11339_/Y _06925_/X vssd1 vssd1 vccd1 vccd1 _11340_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _11557_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__xnor2_1
X_13010_ _13134_/A hold254/X vssd1 vssd1 vccd1 vccd1 _13303_/D sky130_fd_sc_hd__and2_1
XANTENNA__06673__A_N _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ fanout40/X _10222_/A2 _07255_/Y _07137_/Y vssd1 vssd1 vccd1 vccd1 _10223_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07836__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11382__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ hold222/A hold261/A _10153_/C vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__or3_1
XFILLER_0_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13123__B2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nand2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11437__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__A1 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _10987_/B _10987_/A vssd1 vssd1 vccd1 vccd1 _11098_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _12737_/B _12725_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XFILLER_0_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ reg1_val[8] _12657_/B vssd1 vssd1 vccd1 vccd1 _12656_/Y sky130_fd_sc_hd__nor2_1
X_12587_ _12572_/B _12580_/B _12610_/A vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__o21ai_2
X_11607_ _11781_/S _11607_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__or2_1
XFILLER_0_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12636__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11538_ _06941_/X _11537_/X _07068_/A _06940_/B vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11469_ _11900_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ hold291/X _13207_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _13144_/A hold278/X vssd1 vssd1 vccd1 vccd1 _13350_/D sky130_fd_sc_hd__and2_1
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _07701_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07700_/X sky130_fd_sc_hd__or2_1
X_08680_ _08748_/A _08746_/A _08680_/C _08680_/D vssd1 vssd1 vccd1 vccd1 _08751_/B
+ sky130_fd_sc_hd__nand4b_2
XANTENNA__09172__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ fanout79/X fanout77/X fanout75/X fanout73/X vssd1 vssd1 vccd1 vccd1 _07632_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06809__B _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _10326_/A fanout28/X _07218_/Y _07944_/B vssd1 vssd1 vccd1 vccd1 _07563_/B
+ sky130_fd_sc_hd__a22o_1
X_09301_ _09301_/A _09301_/B _09301_/C vssd1 vssd1 vccd1 vccd1 _09305_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07493_ fanout75/X _10227_/B1 _10463_/A1 fanout71/X vssd1 vssd1 vccd1 vccd1 _07494_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ _09233_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09232_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09163_ _09161_/X _09162_/X _09385_/S vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10347__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_A _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _08183_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ _09095_/A _09095_/B vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08045_ _07950_/B _08045_/B vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10167__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07032__A1 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07032__B2 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09996_ _09996_/A _10128_/A _10267_/A _10319_/A vssd1 vssd1 vccd1 vccd1 _09996_/Y
+ sky130_fd_sc_hd__nor4_1
XANTENNA__09309__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__B1 _11258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ fanout60/X _10463_/B2 _10228_/A fanout52/X vssd1 vssd1 vccd1 vccd1 _08948_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10810__A _10810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _09008_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07829_ _07829_/A _07829_/B vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07335__A2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _11359_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06719__B _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _09710_/B _10267_/X _10769_/Y _10770_/Y _10768_/Y vssd1 vssd1 vccd1 vccd1
+ _10772_/B sky130_fd_sc_hd__o311a_4
XANTENNA__07099__A1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A2 _07048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _12516_/B _12510_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ _12621_/A curr_PC[1] _12525_/S vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12372_ _12405_/B _12372_/B vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08950__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ _11109_/X _11506_/A _11322_/X _10889_/X _11320_/X vssd1 vssd1 vccd1 vccd1
+ _11323_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ curr_PC[15] _11255_/B vssd1 vssd1 vccd1 vccd1 _11254_/X sky130_fd_sc_hd__or2_1
X_10205_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11355__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__B2 _09297_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__A1 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _11185_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11186_/B sky130_fd_sc_hd__xnor2_2
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10137_/C sky130_fd_sc_hd__nor2_1
X_10067_ _10067_/A1 fanout22/X fanout15/X _10490_/A vssd1 vssd1 vccd1 vccd1 _10068_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08523__A1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__B2 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _10968_/A _10968_/B _10968_/C vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08287__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ reg1_val[18] _12767_/B vssd1 vssd1 vccd1 vccd1 _12709_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _12639_/A _12639_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xnor2_4
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09675__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07014__A1 _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09003__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _09851_/B _09851_/A vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__nand2b_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _06993_/A _06994_/B vssd1 vssd1 vccd1 vccd1 _06993_/Y sky130_fd_sc_hd__xnor2_4
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__xor2_1
X_08801_ _08798_/X _12229_/B vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__nand2b_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08543_/A _08672_/B _08543_/B vssd1 vssd1 vccd1 vccd1 _08732_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__09711__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08594_ _12785_/A _08594_/A2 _07043_/Y vssd1 vssd1 vccd1 vccd1 _08595_/D sky130_fd_sc_hd__o21ai_1
X_07614_ _10937_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07618_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07545_ _07665_/A _07665_/B _07524_/X vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13152__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _07475_/A _07518_/A vssd1 vssd1 vccd1 vccd1 _07551_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__B2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09215_ _09199_/X _09214_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ _09146_/A _09858_/A vssd1 vssd1 vccd1 vccd1 _10310_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07089__C _07089_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08986__D1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07253__A1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09100_/A sky130_fd_sc_hd__xnor2_2
X_08028_ _08649_/B fanout83/X fanout79/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08029_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__A1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09979_ _09840_/A _09839_/B _09837_/Y vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12990_ _13144_/A hold238/X vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__and2_1
XANTENNA__12301__A2 _09728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _12085_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _12020_/D sky130_fd_sc_hd__xnor2_2
X_11872_ _11872_/A _11872_/B vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10823_ _10823_/A vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__inv_2
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11371__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__B2 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ _10633_/A _10633_/B _10636_/A vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__A2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10685_ _10654_/Y _10655_/X _10657_/Y _11946_/A _10684_/X vssd1 vssd1 vccd1 vccd1
+ _10685_/X sky130_fd_sc_hd__o221a_1
X_12424_ hold263/A _12387_/X _12347_/B vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_105_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12355_ _09237_/Y _12346_/X _12347_/Y _12351_/Y _12354_/X vssd1 vssd1 vccd1 vccd1
+ _12356_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07244__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ _11306_/A _11306_/B vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08992__A1 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12286_ _12285_/A _12285_/B _12285_/Y _09226_/Y vssd1 vssd1 vccd1 vccd1 _12304_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08992__B2 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ _09252_/B _11236_/Y _11237_/S vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__mux2_1
X_11168_ _11168_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11170_/A sky130_fd_sc_hd__and2_1
X_10119_ _10119_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__xnor2_1
X_11099_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11101_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10303__A1 _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11281__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__A1 _06964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10067__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07330_ _10937_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13005__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ _08823_/A _08823_/B _08820_/A vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07261_ _07171_/X _10712_/A _07182_/Y _07212_/X vssd1 vssd1 vccd1 vccd1 _07262_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12359__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _07192_/A _07192_/B _07192_/C vssd1 vssd1 vccd1 vccd1 _07193_/B sky130_fd_sc_hd__and3_1
XANTENNA__08590__A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ curr_PC[4] _10035_/C vssd1 vssd1 vccd1 vccd1 _09902_/X sky130_fd_sc_hd__or2_1
X_09833_ _09681_/A _09681_/B _09679_/Y vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__a21bo_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11456__A _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ _06975_/A _06967_/A _06967_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _06978_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__10360__A _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _11813_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06761__A3 _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__and2_1
X_09695_ _09695_/A _09695_/B vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08646_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _08712_/A sky130_fd_sc_hd__xnor2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08577_ _08597_/A vssd1 vssd1 vccd1 vccd1 _08577_/Y sky130_fd_sc_hd__inv_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ _07114_/X _07944_/B fanout28/X _07146_/Y vssd1 vssd1 vccd1 vccd1 _07529_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11270__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ _07460_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__and2_1
X_10470_ _10469_/B _10469_/C _10469_/A vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09596__A _11238_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11558__B1 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _09016_/A _09016_/B _09015_/A vssd1 vssd1 vccd1 vccd1 _09139_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__and2_1
XANTENNA__08974__A1 _06973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08974__B2 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12071_ _12138_/B _12071_/B vssd1 vssd1 vccd1 vccd1 _12073_/C sky130_fd_sc_hd__and2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _09557_/X _11021_/X _11237_/S vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__mux2_1
X_12973_ hold240/A _13095_/B2 _13158_/A2 hold207/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__a22o_1
X_11924_ _12007_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11926_/B sky130_fd_sc_hd__and2_1
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07162__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _11685_/X _12016_/A _11853_/Y vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06907__B _06907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11786_ _11700_/B _11702_/B _11700_/A vssd1 vssd1 vccd1 vccd1 _11787_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__11797__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ curr_PC[11] _10926_/C vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11261__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ _10738_/A _10738_/B vssd1 vssd1 vccd1 vccd1 _10862_/B sky130_fd_sc_hd__and2_1
XFILLER_0_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07465__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07465__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12322_/B _12368_/A _12406_/B _12326_/X vssd1 vssd1 vccd1 vccd1 _12407_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _10668_/A vssd1 vssd1 vccd1 vccd1 _10668_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ _06656_/A _12336_/X _12337_/Y vssd1 vssd1 vccd1 vccd1 _12356_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ _12269_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__nand2_1
X_06830_ _06722_/Y _06828_/Y _06829_/X vssd1 vssd1 vccd1 vccd1 _06830_/Y sky130_fd_sc_hd__a21oi_1
X_06761_ _06799_/A _06801_/B1 _12652_/B _06760_/X vssd1 vssd1 vccd1 vccd1 _07264_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10827__A2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06692_ _06706_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _06692_/Y sky130_fd_sc_hd__nor2_1
X_09480_ _09480_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__nor2_1
X_08500_ _07010_/Y _09450_/B1 _07263_/Y _07018_/X vssd1 vssd1 vccd1 vccd1 _08501_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12819__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__S _09180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _08533_/B _09468_/B2 _08591_/B1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08432_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10339__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ fanout50/X _10233_/B2 _10233_/A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 _07314_/B
+ sky130_fd_sc_hd__o22a_1
X_08293_ _08556_/A _08293_/B vssd1 vssd1 vccd1 vccd1 _08338_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07244_ fanout85/X fanout83/X _10466_/A fanout79/X vssd1 vssd1 vccd1 vccd1 _07245_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__A1 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _07175_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07175_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_42_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ _08650_/A _09671_/B _09669_/Y vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__a21oi_2
X_06959_ _06963_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _06959_/Y sky130_fd_sc_hd__nand2_1
X_09747_ hold271/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__xor2_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11914__A _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__B1 _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _11645_/B _09678_/B vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08495__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A _08629_/B _08629_/C vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__or3_2
X_11640_ _11559_/A _07193_/A wire8/X _11639_/Y vssd1 vssd1 vccd1 vccd1 _11641_/B sky130_fd_sc_hd__a31o_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _11571_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10522_ _10522_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _13324_/CLK hold183/X vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13241_ _13375_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_10453_ _11172_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__xnor2_1
X_13172_ hold295/A _13171_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10384_ _10384_/A _10384_/B _10384_/C vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__or3_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08947__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ curr_PC[25] _12186_/C vssd1 vssd1 vccd1 vccd1 _12124_/C sky130_fd_sc_hd__and2_1
XFILLER_0_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _12202_/B fanout9/X fanout4/X fanout67/X vssd1 vssd1 vccd1 vccd1 _12055_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10712__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__B _11808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _10533_/X _11004_/A _11002_/X vssd1 vssd1 vccd1 vccd1 _11005_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12259__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ _12978_/A hold268/X vssd1 vssd1 vccd1 vccd1 _13276_/D sky130_fd_sc_hd__and2_1
X_11907_ _11906_/B _11907_/B vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06637__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12887_ hold165/X _13338_/Q vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08883__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10690__B1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11769_ _12087_/A _11769_/B vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12431__B2 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07749__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12195__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08980_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07931_ _07931_/A _07931_/B vssd1 vssd1 vccd1 vccd1 _07932_/C sky130_fd_sc_hd__nand2_1
X_07862_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__and2_1
X_06813_ _07264_/A reg1_val[6] vssd1 vssd1 vccd1 vccd1 _06813_/Y sky130_fd_sc_hd__nand2b_1
X_09601_ _09552_/Y _09600_/X _12504_/S vssd1 vssd1 vccd1 vccd1 _09601_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07374__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _09533_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__and2_1
X_07793_ _07791_/A _07791_/B _07863_/A vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06744_ reg2_val[9] _06767_/A vssd1 vssd1 vccd1 vccd1 _06744_/X sky130_fd_sc_hd__and2_1
XANTENNA__11473__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_A _06631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ _11711_/S _06675_/B vssd1 vssd1 vccd1 vccd1 _06683_/C sky130_fd_sc_hd__nor2_2
XANTENNA__11453__B wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _09462_/A _09462_/B _09464_/A vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09394_ _09189_/X _09192_/X _09396_/S vssd1 vssd1 vccd1 vccd1 _09394_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07429__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07429__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12973__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ _08336_/A _08336_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07227_ _10468_/A vssd1 vssd1 vccd1 vccd1 _10942_/A sky130_fd_sc_hd__inv_6
XANTENNA__07097__C _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07158_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07601__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12504__S _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ reg1_val[18] reg1_val[19] _07089_/C vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__or3_4
XANTENNA__07394__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07601__B2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout120 _07174_/Y vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__clkbuf_8
Xfanout131 _07078_/X vssd1 vssd1 vccd1 vccd1 _08507_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout164 _11115_/A vssd1 vssd1 vccd1 vccd1 _12178_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout153 _06995_/X vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__clkbuf_8
Xfanout142 _09324_/A vssd1 vssd1 vccd1 vccd1 _08619_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11161__B2 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 _09225_/X vssd1 vssd1 vccd1 vccd1 _12395_/A1 sky130_fd_sc_hd__buf_4
Xfanout175 _07195_/B vssd1 vssd1 vccd1 vccd1 _07299_/B sky130_fd_sc_hd__buf_8
XANTENNA__07904__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _07175_/X _12842_/A2 hold36/X _13144_/A vssd1 vssd1 vccd1 vccd1 hold37/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09657__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12741_/A _12747_/A vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ reg1_val[11] _12673_/B vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__nand2_1
X_11623_ hold295/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11708_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _11554_/A _11554_/B vssd1 vssd1 vccd1 vccd1 _11571_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _11386_/A _11988_/A _11387_/A _11388_/Y vssd1 vssd1 vccd1 vccd1 _11490_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ _10505_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07840__A1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07840__B2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13224_ _12950_/A _13224_/B vssd1 vssd1 vccd1 vccd1 _13224_/Y sky130_fd_sc_hd__nand2b_1
X_10436_ _09223_/Y _10423_/Y _10424_/X _09243_/B _10435_/X vssd1 vssd1 vccd1 vccd1
+ _10436_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06920__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ _13155_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _13156_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10723__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ _10368_/B _10368_/A vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__and2b_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12106_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12106_/Y sky130_fd_sc_hd__xnor2_1
X_13086_ _13109_/A hold266/X vssd1 vssd1 vccd1 vccd1 _13339_/D sky130_fd_sc_hd__and2_1
X_10298_ _10166_/A _10163_/Y _10165_/B vssd1 vssd1 vccd1 vccd1 _10302_/A sky130_fd_sc_hd__o21a_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12037_ hold204/A _12037_/B vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__or2_1
XANTENNA__09008__B _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__S _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12101__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A2 _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ _12857_/B _13202_/B _12855_/X vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08608__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08130_ _09468_/B2 _08274_/B fanout74/X _08591_/B1 vssd1 vssd1 vccd1 vccd1 _08131_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12955__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08061_ _08790_/A _08786_/A vssd1 vssd1 vccd1 vccd1 _08061_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07012_ _06975_/A _06974_/X _06975_/Y _06967_/Y vssd1 vssd1 vccd1 vccd1 _07012_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__B2 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A1 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08963_ _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ _07988_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07914_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12340__B1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ _08894_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _08896_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07845_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _08320_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06727_ _11030_/S _06727_/B vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__nor2_1
X_09515_ _07944_/B _07250_/X _07255_/Y fanout28/X vssd1 vssd1 vccd1 vccd1 _09516_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10654__B1 _10810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ _09766_/A _09446_/B vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__xor2_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _06706_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _06658_/Y sky130_fd_sc_hd__nor2_1
X_06589_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06589_/X sky130_fd_sc_hd__and4bb_1
X_09377_ _09260_/X _09440_/C _09376_/Y vssd1 vssd1 vccd1 vccd1 _09377_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08075__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08259_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ fanout25/X fanout13/X fanout11/X fanout27/X vssd1 vssd1 vccd1 vccd1 _11271_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09575__A1 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11382__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _10221_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11382__B2 _11456_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _10149_/X _10151_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__mux2_1
X_10083_ _11557_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__xnor2_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08948__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10893__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ reg1_val[20] _12767_/B _12720_/A vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ _12654_/A _12651_/Y _12653_/B vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ _12584_/X _12586_/B vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_108_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ _11606_/A _11606_/B vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _11509_/Y _11510_/X _11512_/Y _11946_/A _11536_/X vssd1 vssd1 vccd1 vccd1
+ _11537_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap117 _07178_/Y vssd1 vssd1 vccd1 vccd1 _10327_/B2 sky130_fd_sc_hd__clkbuf_8
X_11468_ _12202_/B fanout44/X _12257_/A fanout46/X vssd1 vssd1 vccd1 vccd1 _11469_/B
+ sky130_fd_sc_hd__o22a_1
Xmax_cap139 _07201_/B vssd1 vssd1 vccd1 vccd1 _07202_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__B _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__xnor2_1
X_13207_ _13207_/A _13207_/B vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10453__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _10417_/Y _10419_/B vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ hold277/X _13186_/A2 _13137_/X _13143_/B2 vssd1 vssd1 vccd1 vccd1 hold278/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ hold89/X _13071_/A2 _13071_/B1 hold12/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold90/A sky130_fd_sc_hd__o221a_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07329__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A _12065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07630_ _09787_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07561_ _10081_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__xnor2_1
X_09300_ _09300_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _09301_/C sky130_fd_sc_hd__or3_1
XANTENNA__12827__B _12841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ _07492_/A _07492_/B vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _12395_/A1 _09230_/X _06876_/Y vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12389__B1 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__A1 _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ reg1_val[5] reg1_val[26] _09180_/S vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11061__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _08624_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _08183_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07002__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09093_ _06875_/A wire8/X _09670_/A vssd1 vssd1 vccd1 vccd1 _09095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _08054_/B _08054_/A vssd1 vssd1 vccd1 vccd1 _08056_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10167__A2 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07032__A2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09309__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11116__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08999_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10810__B _10810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _09930_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _08878_/B sky130_fd_sc_hd__xnor2_2
X_07828_ _07847_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07828_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07759_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07759_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout31_A _07193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _10270_/A _10270_/B _10769_/A _11003_/A vssd1 vssd1 vccd1 vccd1 _10770_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _10315_/A _09670_/A _09428_/Y vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__a21o_1
X_12440_ _12446_/A _12440_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
XFILLER_0_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12371_ _12157_/B _12271_/C _12369_/X _12370_/X vssd1 vssd1 vccd1 vccd1 _12372_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11322_ _11322_/A _11506_/A vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__and2_1
X_11253_ _11253_/A _11253_/B _11253_/C _11252_/X vssd1 vssd1 vccd1 vccd1 _11253_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10158__A2 _10158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _10075_/A _10075_/B _10073_/Y vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07023__A2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _11184_/A _11184_/B vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10135_ _09549_/B _10129_/C _10133_/Y _10650_/A vssd1 vssd1 vccd1 vccd1 _10136_/B
+ sky130_fd_sc_hd__o211a_1
X_10066_ _10066_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08523__A2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10968_ _10968_/A _10968_/B _10968_/C vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__or3_1
XANTENNA__10618__B1 _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09484__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12647__B _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ reg1_val[18] _12767_/B vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10899_ _12025_/S _06824_/Y _10898_/Y vssd1 vssd1 vccd1 vccd1 _10899_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12638_ _12636_/Y _12638_/B vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12569_ _12574_/C _12569_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10183__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A2 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ _08800_/A _08800_/B _12229_/B vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__and3_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _06967_/A _06966_/C _07074_/B vssd1 vssd1 vccd1 vccd1 _06994_/B sky130_fd_sc_hd__a21o_2
XANTENNA__13099__B2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _09653_/B _09656_/B _09653_/A vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__o21ba_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12846__A1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08731_ _08728_/A _08728_/B _08730_/B _08730_/A _10656_/B vssd1 vssd1 vccd1 vccd1
+ _08731_/X sky130_fd_sc_hd__a221o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _08712_/A _08712_/B _08645_/X vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__a21o_1
X_07613_ _07402_/B _07146_/Y _07153_/Y fanout41/X vssd1 vssd1 vccd1 vccd1 _07614_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout166_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ _08601_/A _08601_/B vssd1 vssd1 vccd1 vccd1 _08602_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11742__A _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11821__A2 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07475_ _07475_/A _07475_/B _07474_/X vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__or3b_1
X_09214_ _09206_/X _09213_/X _10148_/S vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _09145_/A _09145_/B vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07253__A2 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _09077_/B vssd1 vssd1 vccd1 vccd1 _09076_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10793__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08027_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11888__A2 _11864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _09978_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__xor2_4
XANTENNA_fanout79_A _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _10937_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08931_/B sky130_fd_sc_hd__xor2_1
X_11940_ _11601_/B _11939_/Y _11938_/X vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__08505__A2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11872_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10822_ _10822_/A _10822_/B vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__xnor2_1
X_10753_ _10753_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _10755_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ _10660_/Y _10661_/X _10671_/X _10683_/X vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08961__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _09252_/X _12421_/Y _12422_/Y vssd1 vssd1 vccd1 vccd1 _12423_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ _09222_/Y _09559_/Y _09574_/X _09155_/S _12353_/X vssd1 vssd1 vccd1 vccd1
+ _12354_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07244__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _11305_/A _11305_/B _11305_/C vssd1 vssd1 vccd1 vccd1 _11306_/B sky130_fd_sc_hd__and3_1
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08992__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12285_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11328__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11236_ _11236_/A vssd1 vssd1 vccd1 vccd1 _11236_/Y sky130_fd_sc_hd__inv_2
X_11167_ _11557_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12828__A1 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10118_ _09986_/A _09986_/B _09984_/Y vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10839__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _11098_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__and2_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10049_ _10736_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10303__A2 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10067__B2 _10490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10067__A1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11803__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07260_ _07611_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07273_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _07192_/A _07192_/B _07192_/C vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__08590__B _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ curr_PC[4] _10035_/C vssd1 vssd1 vccd1 vccd1 _09901_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09832_ _09954_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11456__B _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _10213_/A _07581_/A _07581_/B _07345_/X _10326_/A vssd1 vssd1 vccd1 vccd1
+ _09764_/B sky130_fd_sc_hd__a32o_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ _06975_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _06975_/Y sky130_fd_sc_hd__nor2_1
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08111__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _09694_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08645_ _08646_/B _08646_/A vssd1 vssd1 vccd1 vccd1 _08645_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08576_/A _08588_/A vssd1 vssd1 vccd1 vccd1 _08597_/A sky130_fd_sc_hd__nand2_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06566__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _11361_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__xnor2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08120__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ _09630_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07460_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ _07389_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07396_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11558__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__B2 _07193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ _09128_/A _09128_/B vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_121_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08974__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _09356_/A _09059_/B vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _12070_/A _12070_/B vssd1 vssd1 vccd1 vccd1 _12071_/B sky130_fd_sc_hd__or2_1
X_11021_ _10012_/X _10014_/X _11021_/S vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08187__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ _12978_/A hold241/X vssd1 vssd1 vccd1 vccd1 _13284_/D sky130_fd_sc_hd__and2_1
X_11923_ _11923_/A _11923_/B _11923_/C vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__or3_1
XFILLER_0_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12478__A _12647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__A1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _11854_/A _11937_/A vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11246__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ _09148_/Y _10773_/Y _10774_/X _10804_/X vssd1 vssd1 vccd1 vccd1 _10805_/X
+ sky130_fd_sc_hd__a31o_1
X_11785_ _11785_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11797__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10736_ _10736_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10738_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09787__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07465__A2 _09297_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _09566_/X _09572_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12406_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ _11359_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__xnor2_2
X_13386_ instruction[4] vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
XFILLER_0_121_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12337_ _06656_/A _12336_/X _09226_/Y vssd1 vssd1 vccd1 vccd1 _12337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12268_ _12268_/A vssd1 vssd1 vccd1 vccd1 _12269_/B sky130_fd_sc_hd__inv_2
XFILLER_0_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11557__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _11219_/A _11414_/A vssd1 vssd1 vccd1 vccd1 _11219_/Y sky130_fd_sc_hd__nand2_1
X_12199_ _12199_/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__or2_1
XANTENNA__11721__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ reg2_val[6] _06794_/B vssd1 vssd1 vccd1 vccd1 _06760_/X sky130_fd_sc_hd__and2_1
X_06691_ instruction[28] _06699_/B vssd1 vssd1 vccd1 vccd1 _12632_/B sky130_fd_sc_hd__and2_4
XFILLER_0_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07770__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08459_/B sky130_fd_sc_hd__or2_1
XANTENNA__06900__A1 _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08361_ _08361_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12985__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ _10231_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07372_/A sky130_fd_sc_hd__xnor2_1
X_08292_ _08507_/A2 _08553_/A2 _08551_/B1 _08533_/B vssd1 vssd1 vccd1 vccd1 _08293_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12835__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ _07243_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13012__A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ _07175_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07174_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11356__A1_N _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11712__A1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09815_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__nor2_1
X_06958_ _07243_/A _07251_/A _06958_/C _06958_/D vssd1 vssd1 vccd1 vccd1 _06963_/B
+ sky130_fd_sc_hd__nor4_4
X_09746_ hold322/A hold265/A _13338_/Q _10158_/A2 vssd1 vssd1 vccd1 vccd1 _09747_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__06995__S _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09677_ _09928_/A fanout9/A fanout5/X _09815_/A vssd1 vssd1 vccd1 vccd1 _09678_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06889_ _06927_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09235_/A sky130_fd_sc_hd__or2_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__A1 _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ _08622_/A _08622_/B _08620_/Y vssd1 vssd1 vccd1 vccd1 _08629_/C sky130_fd_sc_hd__o21ba_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08559_ _08559_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _08561_/C sky130_fd_sc_hd__xor2_1
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _10522_/B _10522_/A vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__nand2b_1
X_13240_ _13374_/CLK _13240_/D vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ fanout64/X fanout35/X fanout33/X fanout58/X vssd1 vssd1 vccd1 vccd1 _10453_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13171_ _13171_/A _13171_/B vssd1 vssd1 vccd1 vccd1 _13171_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10383_ _10384_/A _10384_/B _10384_/C vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08947__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ curr_PC[25] _12186_/C vssd1 vssd1 vccd1 vccd1 _12124_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ _12053_/A1 _12050_/X _12052_/Y _12049_/X vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__a31o_4
X_11004_ _11004_/A vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12259__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ hold285/A _13095_/B2 _13158_/A2 hold267/X vssd1 vssd1 vccd1 vccd1 hold268/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06918__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _11907_/B _11906_/B vssd1 vssd1 vccd1 vccd1 _12001_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12886_ hold265/X hold46/X vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08883__B2 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08883__A1 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _11837_/A _11988_/A vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06894__B1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10690__A1 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11768_/A _11939_/A vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12967__B1 _13158_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06934__A _11975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _11359_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10721_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__or2_1
XANTENNA__06653__B _07026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _13375_/CLK _13369_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12195__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11287__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ _07930_/A _07930_/B _07930_/C vssd1 vssd1 vccd1 vccd1 _07931_/B sky130_fd_sc_hd__or3_1
XFILLER_0_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _07861_/A _07931_/A _07861_/C vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__and3_1
X_06812_ _10008_/A _06810_/Y _06811_/Y vssd1 vssd1 vccd1 vccd1 _06812_/X sky130_fd_sc_hd__o21a_1
X_09600_ _12029_/A _09554_/X _09599_/X vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11734__B _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06743_ _06743_/A _10675_/S vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ _09350_/A _09350_/B _09348_/Y vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08323__B1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ reg1_val[20] _06996_/A vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__and2b_1
X_09462_ _09462_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09464_/B sky130_fd_sc_hd__nor2_1
X_09393_ _09186_/X _09188_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09393_/X sky130_fd_sc_hd__mux2_1
X_08413_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout246_A _06893_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08344_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07429__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08320_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _08336_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07226_ reg1_val[13] _07226_/B vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13352_/CLK sky130_fd_sc_hd__clkbuf_8
X_07157_ _09766_/A _07157_/B vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07601__A2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07089_/C sky130_fd_sc_hd__or2_2
Xfanout121 _08320_/A vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__clkbuf_16
Xfanout110 _07213_/Y vssd1 vssd1 vccd1 vccd1 _10067_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout165 _12347_/B vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__buf_4
Xfanout132 _07078_/X vssd1 vssd1 vccd1 vccd1 _10233_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout143 _07129_/Y vssd1 vssd1 vccd1 vccd1 _09324_/A sky130_fd_sc_hd__buf_4
Xfanout154 _08633_/B vssd1 vssd1 vccd1 vccd1 _08619_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07365__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 _12782_/Y vssd1 vssd1 vccd1 vccd1 _12842_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout187 _09149_/X vssd1 vssd1 vccd1 vccd1 _11889_/A1 sky130_fd_sc_hd__buf_4
Xfanout198 _13071_/B1 vssd1 vssd1 vccd1 vccd1 _13053_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__07365__B2 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__B1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout61_A _06999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _09579_/A _09576_/Y _09578_/B vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _12740_/A _12740_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ _12676_/B _12671_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
X_11622_ hold237/A _11529_/B _11705_/B _11621_/Y _12433_/A1 vssd1 vssd1 vccd1 vccd1
+ _11630_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13071__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11554_/A _11554_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _11381_/A _11381_/B _11392_/A vssd1 vssd1 vccd1 vccd1 _11494_/A sky130_fd_sc_hd__a21o_1
X_10504_ _10504_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10505_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07840__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ _13236_/A hold280/X vssd1 vssd1 vccd1 vccd1 _13368_/D sky130_fd_sc_hd__and2_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12491__A _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _10426_/Y _10427_/X _10434_/Y _09196_/S _10433_/X vssd1 vssd1 vccd1 vccd1
+ _10435_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _13187_/A hold298/X vssd1 vssd1 vccd1 vccd1 _13353_/D sky130_fd_sc_hd__and2_1
X_10366_ _10515_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__or2_1
X_12105_ _12103_/Y _12105_/B vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__and2b_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10280_/A _09886_/B _10290_/Y _10291_/X _10296_/X vssd1 vssd1 vccd1 vccd1
+ _10297_/X sky130_fd_sc_hd__o221a_1
X_13085_ hold265/X _13222_/A2 _13084_/X _13095_/B2 vssd1 vssd1 vccd1 vccd1 hold266/A
+ sky130_fd_sc_hd__a22o_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12036_ _10282_/X _12035_/Y _12421_/B vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08553__B1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09305__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ _13197_/A _13198_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ hold311/X hold80/X vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08060_ _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08786_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07011_ _07011_/A _07011_/B vssd1 vssd1 vccd1 vccd1 _07011_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__B2 _12202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07044__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09186__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__and2b_1
X_07913_ _07954_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__xnor2_1
X_08893_ _08894_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout196_A _06925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07844_ _07867_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07898__A2 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07775_ _08521_/A2 _08274_/B fanout74/X _08551_/A2 vssd1 vssd1 vccd1 vccd1 _07776_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10103__B1 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06726_ reg1_val[13] _07255_/A vssd1 vssd1 vccd1 vccd1 _06727_/B sky130_fd_sc_hd__nor2_1
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__nor2_1
X_06657_ instruction[33] _06657_/B vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__and2_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10654__A1 _11863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ _07539_/B _07212_/X _07218_/Y fanout37/X vssd1 vssd1 vccd1 vccd1 _09446_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06588_ _06927_/A _06588_/B vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__nor2_8
X_09376_ _09260_/X _09440_/C _09148_/Y vssd1 vssd1 vccd1 vccd1 _09376_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11603__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ _08624_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _08267_/A _08267_/B _08218_/Y vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__a21o_1
X_07209_ _07210_/A _07210_/B vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__nor2_1
X_10220_ _10221_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__nand2b_1
X_08189_ _08591_/B1 _08274_/B fanout74/X _08619_/B1 vssd1 vssd1 vccd1 vccd1 _08190_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _09432_/X _10150_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _11645_/A fanout27/X fanout25/X fanout51/X vssd1 vssd1 vccd1 vccd1 _10083_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12331__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10984_ _10982_/A _10982_/B _10985_/B vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12723_ _12721_/Y _12723_/B vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ _12610_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__or2_1
XANTENNA__07299__B _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _11776_/A _11604_/B _11604_/C vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11536_ _11516_/Y _11517_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _11536_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__09795__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__nor2_1
X_13206_ _13206_/A _13206_/B vssd1 vssd1 vccd1 vccd1 _13207_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10734__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap118 _07175_/X vssd1 vssd1 vccd1 vccd1 _10222_/A2 sky130_fd_sc_hd__buf_6
X_11398_ _11396_/X _11398_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__and2b_1
X_10418_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ hold305/A _13136_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__mux2_1
X_10349_ _12068_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10351_/B sky130_fd_sc_hd__xor2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _07135_/C _13072_/A2 hold127/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__o21a_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11565__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _12278_/A vssd1 vssd1 vccd1 vccd1 _12019_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08526__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__A1 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__B2 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ _08354_/A2 fanout32/X _10966_/A _08184_/B vssd1 vssd1 vccd1 vccd1 _07561_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11833__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _11612_/A _12431_/A2 _08655_/A vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__a21o_1
X_07491_ _07556_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _07491_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13050__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ reg1_val[4] reg1_val[27] _09180_/S vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11061__B2 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _09301_/A _09092_/B vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08112_ _08649_/B fanout75/X fanout71/X _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08113_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07265__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12843__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08054_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06841__B _06964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_A _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout111_A _07213_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09994_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__and2_1
XANTENNA__09309__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10324__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__A _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _09467_/A _07347_/B fanout15/X _09324_/A vssd1 vssd1 vccd1 vccd1 _08877_/B
+ sky130_fd_sc_hd__o22a_1
X_07827_ _09827_/A _07920_/B _07920_/A vssd1 vssd1 vccd1 vccd1 _07847_/B sky130_fd_sc_hd__mux2_1
X_07758_ _09941_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06709_ reg1_val[16] _07074_/A vssd1 vssd1 vccd1 vccd1 _06711_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07689_ _07689_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__xnor2_2
X_09428_ _10315_/A _09670_/A _08655_/A vssd1 vssd1 vccd1 vccd1 _09428_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout24_A _07215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _09360_/A _09360_/B vssd1 vssd1 vccd1 vccd1 _09359_/Y sky130_fd_sc_hd__nor2_1
X_12370_ _12269_/A _12320_/Y _12369_/X _12272_/Y _12322_/B vssd1 vssd1 vccd1 vccd1
+ _12370_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07256__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _11321_/A _11413_/A vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11252_ _09243_/B _11238_/X _11249_/X _11251_/X vssd1 vssd1 vccd1 vccd1 _11252_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08024__A _08566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11184_/B sky130_fd_sc_hd__xor2_2
X_10203_ _10203_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10134_ _10129_/X _10130_/X _10133_/Y _10650_/A vssd1 vssd1 vccd1 vccd1 _10136_/A
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__08959__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _10212_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__or2_1
XANTENNA__10618__A1 _12202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10967_ _10967_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _10968_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10618__B2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09484__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09484__B2 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10898_ _12025_/S _10898_/B vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13017__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07495__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _12706_/A _12716_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09236__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12637_ reg1_val[4] _12637_/B vssd1 vssd1 vccd1 vccd1 _12638_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13032__A2 _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12568_ _12575_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12569_/B sky130_fd_sc_hd__nand2_2
XANTENNA__06942__A _12378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12499_ _12662_/B _12499_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__or2_1
XANTENNA__06661__B _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11519_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10464__A _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold249/X vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _06991_/A _06991_/B vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__nand2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12846__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08730_ _08730_/A _08730_/B vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__nand2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _08707_/A _08710_/A _08660_/Y _08658_/B vssd1 vssd1 vccd1 vccd1 _08712_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_07612_ _07612_/A _07612_/B vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08592_ _09941_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08601_/B sky130_fd_sc_hd__xnor2_1
X_07543_ _07543_/A _07725_/A vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__or2_1
XANTENNA_fanout159_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _09766_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07474_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ _09209_/X _09212_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09213_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ _09145_/A _09145_/B vssd1 vssd1 vccd1 vccd1 _09371_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10374__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09075_ _10234_/A _09075_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__xnor2_2
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__buf_6
X_08026_ _09941_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__B _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _09975_/Y _09977_/B vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12298__B1 _12393_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _07101_/Y _07402_/B fanout41/X _07114_/X vssd1 vssd1 vccd1 vccd1 _08929_/B
+ sky130_fd_sc_hd__a22o_1
X_08859_ _08605_/A _07593_/Y _08857_/Y _12619_/A vssd1 vssd1 vccd1 vccd1 _08860_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06921__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10821_ _10821_/A _10822_/B vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10752_ _10752_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10753_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08019__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__A1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ _09223_/Y _10669_/X _10682_/Y _09196_/S _10681_/X vssd1 vssd1 vccd1 vccd1
+ _10683_/X sky130_fd_sc_hd__o221a_1
X_12422_ _09252_/X _12421_/Y _09243_/B vssd1 vssd1 vccd1 vccd1 _12422_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _06605_/X _11966_/B _12352_/Y _06607_/B _12396_/A vssd1 vssd1 vccd1 vccd1
+ _12353_/X sky130_fd_sc_hd__a221o_1
X_11304_ _11305_/A _11305_/B _11305_/C vssd1 vssd1 vccd1 vccd1 _11306_/A sky130_fd_sc_hd__a21oi_1
X_12284_ _06868_/Y _12283_/Y _12378_/S vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _10284_/X _10286_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11166_ fanout25/X _12257_/A fanout13/X fanout27/X vssd1 vssd1 vccd1 vccd1 _11167_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07593__A _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13344_/CLK sky130_fd_sc_hd__clkbuf_8
X_10117_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10839__A1 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__A2 _12842_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _10463_/B2 _10466_/B _10466_/C _10228_/A _12202_/B vssd1 vssd1 vccd1 vccd1
+ _10049_/B sky130_fd_sc_hd__o32a_1
XANTENNA__09154__A0 _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10839__B2 _11917_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _12080_/A _11999_/B vssd1 vssd1 vccd1 vccd1 _12001_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10067__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13005__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ reg1_val[20] _07190_/B vssd1 vssd1 vccd1 vccd1 _07192_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_54_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09900_ _09866_/Y _09868_/Y _09873_/X _09899_/X _12504_/S vssd1 vssd1 vccd1 vccd1
+ _09900_/X sky130_fd_sc_hd__o41a_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire8 wire8/A vssd1 vssd1 vccd1 vccd1 wire8/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09831_ _09831_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__or2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11456__C _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ _06967_/A _06967_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__a21o_1
X_09762_ _09674_/A _09674_/B _09672_/Y vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__a21o_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__nor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout276_A _13219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09693_ _09692_/A _09692_/B _09694_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ _08644_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08576_/A _08575_/B _08575_/C vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__nand3_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07171_/X _10326_/A _09450_/B1 _07182_/Y vssd1 vssd1 vccd1 vccd1 _07527_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08120__B2 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _07101_/Y _07944_/B fanout28/X _07114_/X vssd1 vssd1 vccd1 vccd1 _07458_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _07415_/A _07415_/B vssd1 vssd1 vccd1 vccd1 _07388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11558__A2 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ _09125_/Y _09127_/B vssd1 vssd1 vccd1 vccd1 _09128_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ _09058_/A _09058_/B _09058_/C vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _08079_/A _08009_/B vssd1 vssd1 vccd1 vccd1 _08011_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08187__A1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11020_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08187__B2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12971_ hold213/X _13095_/B2 _13158_/A2 hold240/X vssd1 vssd1 vccd1 vccd1 hold241/A
+ sky130_fd_sc_hd__a22o_1
X_11922_ _11923_/A _11923_/B _11923_/C vssd1 vssd1 vccd1 vccd1 _12007_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10297__A2 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ _11682_/X _11766_/A _11765_/A vssd1 vssd1 vccd1 vccd1 _11853_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__07162__A2 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11246__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _12029_/A _10776_/X _10780_/X _10803_/Y vssd1 vssd1 vccd1 vccd1 _10804_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _10735_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10862_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10666_ _10666_/A _10666_/B _10666_/C vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__and3_1
X_13385_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
X_12405_ _12405_/A _12405_/B vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__or2_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ _06993_/Y fanout31/X fanout29/X _11749_/A vssd1 vssd1 vccd1 vccd1 _10598_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12336_ _12335_/A _12334_/X _12335_/Y vssd1 vssd1 vccd1 vccd1 _12336_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _12267_/A _12267_/B _12267_/C vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _11000_/Y _11414_/A _11216_/X vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__a21o_1
X_12198_ _12199_/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__nand2_1
X_11149_ curr_PC[13] curr_PC[14] _11149_/C vssd1 vssd1 vccd1 vccd1 _11255_/B sky130_fd_sc_hd__and3_1
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08866__B _08866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ _11626_/S _06690_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__or2_2
XFILLER_0_78_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08360_ _08624_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07311_ fanout60/X _08590_/B fanout52/X _09648_/A vssd1 vssd1 vccd1 vccd1 _07312_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08338_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07242_ _07243_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07242_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__09189__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07173_ _07113_/A _06954_/B _06958_/C _06956_/X _07299_/B vssd1 vssd1 vccd1 vccd1
+ _07175_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09602__A1 _12053_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09218__A _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09814_ _09814_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09118__B1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ _07255_/A _07175_/A _07179_/A _07213_/A vssd1 vssd1 vccd1 vccd1 _06958_/D
+ sky130_fd_sc_hd__or4_2
X_09745_ hold230/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09745_/X sky130_fd_sc_hd__xor2_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _09240_/A vssd1 vssd1 vccd1 vccd1 _06888_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09676_ _09500_/A _09500_/B _09496_/Y vssd1 vssd1 vccd1 vccd1 _09680_/A sky130_fd_sc_hd__a21oi_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07144__A2 _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ _08632_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _08629_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08580_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08561_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ _07048_/Y _09659_/B2 fanout98/X _09648_/A vssd1 vssd1 vccd1 vccd1 _07510_/B
+ sky130_fd_sc_hd__o22a_1
X_08489_ _08489_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07201__A _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _13170_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13171_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10382_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10384_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _12094_/Y _12095_/X _12098_/Y _12099_/X _12120_/X vssd1 vssd1 vccd1 vccd1
+ _12121_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13153__B2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _12186_/C vssd1 vssd1 vccd1 vccd1 _12052_/Y sky130_fd_sc_hd__inv_2
X_11003_ _11003_/A _11219_/A vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12954_ _12978_/A hold286/X vssd1 vssd1 vccd1 vccd1 _13275_/D sky130_fd_sc_hd__and2_1
XANTENNA__13084__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ _11983_/B _11905_/B vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12885_ hold322/A hold48/X vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08883__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11836_/A _11836_/B vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06894__A1 _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09798__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10690__A2 _10810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A _11854_/A vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10718_ _11917_/B fanout31/X fanout29/X _06993_/Y vssd1 vssd1 vccd1 vccd1 _10719_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12952__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ _10316_/Y _10890_/A _10647_/Y vssd1 vssd1 vccd1 vccd1 _10649_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13368_ _13375_/CLK _13368_/D vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12195__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11568__A _11568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12320_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13299_ _13350_/CLK _13299_/D vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09899__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _07860_/A _07860_/B vssd1 vssd1 vccd1 vccd1 _07861_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08877__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ reg1_val[5] _06811_/B vssd1 vssd1 vccd1 vccd1 _06811_/Y sky130_fd_sc_hd__nand2_1
X_07791_ _07791_/A _07791_/B vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07374__A2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06742_ reg1_val[10] _07213_/A vssd1 vssd1 vccd1 vccd1 _10675_/S sky130_fd_sc_hd__and2_1
X_09530_ _09335_/A _09333_/Y _09332_/X vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__a21bo_1
X_09461_ _09346_/A _09346_/B _09343_/A vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08323__A1 _08619_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B2 _08619_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ _06996_/A reg1_val[20] vssd1 vssd1 vccd1 vccd1 _11711_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09384_/X _09391_/X _11235_/S vssd1 vssd1 vccd1 vccd1 _09392_/X sky130_fd_sc_hd__mux2_1
X_08412_ _08412_/A _08412_/B vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__or2_1
XANTENNA__08087__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06844__B _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10433__A2 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _09403_/S _08274_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ reg1_val[11] reg1_val[12] _07229_/C _07229_/B vssd1 vssd1 vccd1 vccd1 _07226_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07156_ _07146_/Y _07539_/B _07153_/Y fanout37/X vssd1 vssd1 vccd1 vccd1 _07157_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11478__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ _11125_/A _11231_/A _07121_/C vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__or3_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__B1 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout122 _08320_/A vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__buf_12
Xfanout100 _07068_/Y vssd1 vssd1 vccd1 vccd1 _09659_/B2 sky130_fd_sc_hd__buf_6
Xfanout111 _07213_/Y vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__buf_4
Xfanout155 _06991_/Y vssd1 vssd1 vccd1 vccd1 _08633_/B sky130_fd_sc_hd__buf_6
Xfanout144 _07054_/X vssd1 vssd1 vccd1 vccd1 _08572_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout133 _10233_/B2 vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__clkbuf_8
Xfanout199 _13227_/B vssd1 vssd1 vccd1 vccd1 _13071_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _06942_/Y vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__buf_4
Xfanout177 _13072_/A2 vssd1 vssd1 vccd1 vccd1 _13078_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09382__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout188 _07043_/Y vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__buf_12
X_09728_ _09721_/X _09727_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__mux2_2
X_07989_ _07990_/A _07989_/B _07989_/C vssd1 vssd1 vccd1 vccd1 _08154_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout54_A fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09659_ fanout50/X _08184_/B fanout33/X _09659_/B2 vssd1 vssd1 vccd1 vccd1 _09660_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12670_ _12670_/A _12670_/B _12670_/C vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11621_ _11529_/B _11705_/B hold237/A vssd1 vssd1 vccd1 vccd1 _11621_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__B _12756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _12068_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_108_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ _11483_/A _11483_/B vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__xor2_2
X_10503_ _11900_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12772__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ hold279/X _13222_/A2 _13221_/X _12781_/A vssd1 vssd1 vccd1 vccd1 hold280/A
+ sky130_fd_sc_hd__a22o_1
X_10434_ _10288_/S _10287_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10434_/Y sky130_fd_sc_hd__o21ai_2
X_13153_ hold297/X _13186_/A2 _13152_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold298/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12491__B _12492_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ _10365_/A _10365_/B _10365_/C vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__and3_1
X_12104_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__nand2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11137__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10296_ _06757_/Y _12395_/A1 _12394_/A1 _06759_/B _10295_/X vssd1 vssd1 vccd1 vccd1
+ _10296_/X sky130_fd_sc_hd__o221a_1
X_13084_ _13338_/Q _13083_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12035_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08002__B1 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__B1 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08553__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12937_ hold120/X hold314/A vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ hold297/X hold74/X vssd1 vssd1 vccd1 vccd1 _13155_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__06945__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _11733_/A _11733_/B _11732_/A vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12666__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__B _12652_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ hold29/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09805__A1 _09648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__B2 _08590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ _07010_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07010_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__07776__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08241__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _10081_/A _08961_/B vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__xnor2_1
X_07912_ _07908_/A _07908_/B _07957_/A vssd1 vssd1 vccd1 vccd1 _07988_/A sky130_fd_sc_hd__o21bai_1
X_08892_ _09020_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__nor2_1
X_07843_ _08320_/A _07843_/B vssd1 vssd1 vccd1 vccd1 _07867_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06839__B _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A _07043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07016__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__A1 _07111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06725_ reg1_val[13] _07255_/A vssd1 vssd1 vccd1 vccd1 _11030_/S sky130_fd_sc_hd__and2_1
X_09513_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__nor2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06656_ _06656_/A _12285_/A _06656_/C _06655_/X vssd1 vssd1 vccd1 vccd1 _06656_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__10654__A2 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _09930_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__xnor2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06587_ instruction[3] _06588_/B vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__nor2_8
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _09996_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09440_/C sky130_fd_sc_hd__xnor2_2
X_08326_ _08649_/B _10585_/B2 _10067_/A1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 _08327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _08269_/A _08269_/B _08247_/Y vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07208_ reg1_val[18] _07208_/B vssd1 vssd1 vccd1 vccd1 _07210_/B sky130_fd_sc_hd__xnor2_2
X_08188_ _08445_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__xnor2_2
X_07139_ _07138_/B _12132_/A _12193_/A vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08232__B1 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__B2 _13108_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _09568_/X _09571_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10840__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _10081_/A _10081_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10893__A2 _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _10859_/A _11296_/B _10860_/A _10863_/A vssd1 vssd1 vccd1 vccd1 _10985_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ reg1_val[21] _12773_/A vssd1 vssd1 vccd1 vccd1 _12723_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _12651_/Y _12653_/B vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__nand2b_2
X_12584_ _12616_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ _11776_/A _11604_/B _11604_/C vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__or3_1
XFILLER_0_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11535_ _12107_/B1 _11523_/X _11527_/Y _11534_/X vssd1 vssd1 vccd1 vccd1 _11535_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11467_/B sky130_fd_sc_hd__nor2_1
X_13205_ _13226_/A hold292/X vssd1 vssd1 vccd1 vccd1 _13364_/D sky130_fd_sc_hd__and2_1
XANTENNA__11358__B1 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11397_ _11397_/A _11397_/B _11395_/Y vssd1 vssd1 vccd1 vccd1 _11398_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10417_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08223__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _13136_/A _13136_/B vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__xnor2_1
X_10348_ _07402_/B _07250_/X _07255_/Y fanout40/X vssd1 vssd1 vccd1 vccd1 _10349_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ hold126/X _13071_/A2 _13071_/B1 hold89/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold127/A sky130_fd_sc_hd__o221a_1
X_10279_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__or2_1
XANTENNA__12441__S _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _12154_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08526__A1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08526__B2 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11833__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07490_ _07490_/A _07490_/B vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11833__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10197__A _11361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _09156_/X _09159_/X _09722_/S vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11061__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12794__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _08633_/B _10466_/B _10466_/C _09300_/A fanout55/X vssd1 vssd1 vccd1 vccd1
+ _09092_/B sky130_fd_sc_hd__o32a_1
X_08111_ _08566_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08183_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07265__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__A1 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _08012_/X _08040_/B _08041_/Y vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11349__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09962__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09993_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10324__B2 _10490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _12785_/A fanout9/A vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__nor2_2
X_07826_ _07826_/A _07869_/A vssd1 vssd1 vccd1 vccd1 _07920_/B sky130_fd_sc_hd__nand2_1
X_07757_ _08619_/B2 _09659_/B2 fanout98/X _08619_/A2 vssd1 vssd1 vccd1 vccd1 _07758_/B
+ sky130_fd_sc_hd__o22a_1
X_06708_ _07074_/A reg1_val[16] vssd1 vssd1 vccd1 vccd1 _06711_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11824__B2 _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ _07788_/A _07788_/B _07677_/X vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__a21o_1
X_06639_ _06637_/Y _06707_/B1 _06712_/B reg2_val[24] vssd1 vssd1 vccd1 vccd1 _06641_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_09427_ _09427_/A _09427_/B _09415_/X vssd1 vssd1 vccd1 vccd1 _09427_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09358_ _09124_/A _09124_/B _09122_/X vssd1 vssd1 vccd1 vccd1 _09360_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout17_A _08985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07256__B2 fanout71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08309_ _08346_/A _08346_/B _08270_/Y vssd1 vssd1 vccd1 vccd1 _08682_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10835__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11320_ _11108_/A _11213_/Y _11215_/B vssd1 vssd1 vccd1 vccd1 _11320_/X sky130_fd_sc_hd__o21a_1
X_09289_ _10230_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ _09155_/S _11339_/B _11237_/X _09223_/Y vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11182_ _11900_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__xnor2_2
X_10202_ _11169_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__xnor2_1
X_10133_ _10133_/A _10133_/B vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06782__A3 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08975__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ _10966_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10618__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09484__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _10779_/A _10777_/X _10794_/S vssd1 vssd1 vccd1 vccd1 _10898_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07495__A1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__B2 _09114_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ reg1_val[17] _12767_/B vssd1 vssd1 vccd1 vccd1 _12716_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12636_ reg1_val[4] _12637_/B vssd1 vssd1 vccd1 vccd1 _12636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09236__A2 _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08444__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _12575_/C _12567_/B vssd1 vssd1 vccd1 vccd1 _12574_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12498_ _12662_/B _12499_/B vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__nand2_1
X_11518_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__nand2_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _11447_/Y _11539_/B _12053_/A1 vssd1 vssd1 vccd1 vccd1 _11449_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__12960__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__B1 _10466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ _13236_/A hold284/X vssd1 vssd1 vccd1 vccd1 _13346_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _09671_/A _06990_/B vssd1 vssd1 vccd1 vccd1 _06991_/B sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08660_/A vssd1 vssd1 vccd1 vccd1 _08660_/Y sky130_fd_sc_hd__inv_2
X_07611_ _07611_/A _07611_/B vssd1 vssd1 vccd1 vccd1 _07612_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07183__B1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__B1 _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ _08619_/A2 _08619_/B1 _08591_/B1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 _08592_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07542_ _07543_/A _07542_/B _07542_/C _07542_/D vssd1 vssd1 vccd1 vccd1 _07725_/A
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07473_ _07128_/Y _07539_/B fanout37/X _08476_/A vssd1 vssd1 vccd1 vccd1 _07474_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09210_/X _09211_/X _09402_/S vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07238__A1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _09145_/A _09145_/B vssd1 vssd1 vccd1 vccd1 _09143_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06852__B _07029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08986__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09074_ fanout58/X _10233_/B2 _10233_/A1 fanout56/X vssd1 vssd1 vccd1 vccd1 _09075_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout2 fanout3/X vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_4
X_08025_ _08619_/B2 fanout75/X fanout71/X _08619_/A2 vssd1 vssd1 vccd1 vccd1 _08026_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11917__C _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__nand2_1
X_08927_ _09827_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08931_/A sky130_fd_sc_hd__xnor2_1
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08858_/Y sky130_fd_sc_hd__xnor2_2
X_07809_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08789_ _08789_/A _08789_/B _08789_/C vssd1 vssd1 vccd1 vccd1 _08790_/B sky130_fd_sc_hd__and3_1
X_10820_ _10942_/A _07236_/B fanout6/X _10819_/Y vssd1 vssd1 vccd1 vccd1 _10822_/B
+ sky130_fd_sc_hd__o31ai_2
X_10751_ _10752_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10751_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11273__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12421_ reg1_val[30] _12421_/B _12421_/C vssd1 vssd1 vccd1 vccd1 _12421_/Y sky130_fd_sc_hd__nand3_1
X_10682_ _10288_/S _10015_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10682_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12352_ _06605_/X _12431_/A2 _12395_/A1 vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10233__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _11066_/A _11066_/B _11184_/B _11185_/B _11185_/A vssd1 vssd1 vccd1 vccd1
+ _11305_/C sky130_fd_sc_hd__a32oi_2
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12283_ _06858_/A _12162_/A _12160_/X _12282_/X vssd1 vssd1 vccd1 vccd1 _12283_/Y
+ sky130_fd_sc_hd__o31ai_1
X_11234_ _11234_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11165_ _11305_/B _11165_/B vssd1 vssd1 vccd1 vccd1 _11186_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07593__B _07593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__xor2_1
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10839__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ _10942_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__xnor2_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ _11998_/A _11998_/B _11998_/C vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__or3_1
XFILLER_0_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10949_ fanout56/X fanout46/X fanout44/X _11837_/A vssd1 vssd1 vccd1 vccd1 _10950_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12619_ _12619_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06979__B1 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11724__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09830_ _09831_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__nand2_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09761_ _09697_/A _09697_/B _09698_/Y vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__o21ai_4
X_06973_ _06973_/A _12621_/A vssd1 vssd1 vccd1 vccd1 _06973_/Y sky130_fd_sc_hd__nand2_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08713_/B sky130_fd_sc_hd__xor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09692_ _09692_/A _09692_/B vssd1 vssd1 vccd1 vccd1 _09694_/B sky130_fd_sc_hd__nor2_2
XANTENNA__07156__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_A _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08574_ _08600_/A _08600_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08575_/C sky130_fd_sc_hd__a21o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07525_ _07525_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07541_/A sky130_fd_sc_hd__xor2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07024__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08120__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07456_ _11361_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06582__B _06922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07387_ _07387_/A _07387_/B vssd1 vssd1 vccd1 vccd1 _07415_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _09126_/A _09126_/B vssd1 vssd1 vccd1 vccd1 _09127_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__A1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ _09058_/A _09058_/B _09058_/C vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09908__B1 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__S _09385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__B2 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _08079_/A _08009_/B vssd1 vssd1 vccd1 vccd1 _08008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08187__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__and2_1
X_12970_ _12978_/A hold214/X vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__and2_1
X_11921_ _11921_/A _11921_/B vssd1 vssd1 vccd1 vccd1 _11923_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06757__B _07202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _11852_/A _11852_/B vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__nand2_2
X_10803_ _09243_/B _10790_/X _10802_/X vssd1 vssd1 vccd1 vccd1 _10803_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08647__B1 _07153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__nand2_1
X_10734_ _11169_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10736_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _10666_/A _10666_/B _10666_/C vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__a21oi_1
X_13384_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12404_ wire8/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10596_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__xor2_2
X_12335_ _12335_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12335_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12266_ _12267_/A _12267_/B _12267_/C vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11217_ _11217_/A _11321_/A vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__nor2_1
X_12197_ _12197_/A vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__inv_2
X_11148_ _07251_/A _06940_/B _06941_/X _11147_/X vssd1 vssd1 vccd1 vccd1 _11148_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11079_ _11296_/A fanout9/A fanout5/X _11188_/A vssd1 vssd1 vccd1 vccd1 _11080_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06948__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A2 _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__A _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__B _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12434__A1 _11946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07328_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08290_ _08573_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__xnor2_2
X_07241_ _07251_/A _06954_/X _06958_/C _06958_/D _07299_/B vssd1 vssd1 vccd1 vccd1
+ _07243_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07172_ _07169_/Y _07172_/B vssd1 vssd1 vccd1 vccd1 _07172_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_5_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10933__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09813_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09814_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10920__A1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__A1 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__B2 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06956_ _07179_/A _07213_/A vssd1 vssd1 vccd1 vccd1 _06956_/X sky130_fd_sc_hd__or2_1
X_09744_ hold325/A hold285/A hold321/A _10427_/A2 vssd1 vssd1 vccd1 vccd1 _09745_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06887_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09240_/A sky130_fd_sc_hd__nand2_2
X_09675_ _09675_/A _11155_/A vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nor2_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07144__A3 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _08648_/A _08626_/B vssd1 vssd1 vccd1 vccd1 _08632_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13190__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08557_ _08586_/A _08563_/B _08550_/X vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07508_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07718_/B sky130_fd_sc_hd__or2_1
X_08488_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08736_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07439_ _10233_/B2 fanout98/X _10233_/A1 fanout83/X vssd1 vssd1 vccd1 vccd1 _07440_/B
+ sky130_fd_sc_hd__o22a_1
X_10450_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _09109_/A _09109_/B vssd1 vssd1 vccd1 vccd1 _09110_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10381_ _11557_/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__xnor2_2
X_12120_ _12100_/Y _12101_/X _12108_/Y _12119_/X vssd1 vssd1 vccd1 vccd1 _12120_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09409__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ curr_PC[23] curr_PC[24] _12051_/C vssd1 vssd1 vccd1 vccd1 _12186_/C sky130_fd_sc_hd__and3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _10766_/Y _11219_/A _11000_/Y vssd1 vssd1 vccd1 vccd1 _11002_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10911__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ hold321/A _13095_/B2 _13158_/A2 hold285/X vssd1 vssd1 vccd1 vccd1 hold286/A
+ sky130_fd_sc_hd__a22o_1
X_11904_ _11903_/B _11904_/B vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10675__A0 _09886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12884_ _12882_/X _12884_/B vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07540__B1 _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11836_/A _11836_/B vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12416__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11766_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11937_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10427__B1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12967__A2 _13095_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ _11172_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _06683_/C _11695_/X _11696_/Y vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10648_ _10650_/C _10767_/A vssd1 vssd1 vccd1 vccd1 _10890_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _13375_/CLK _13367_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
X_10579_ fanout42/X _07237_/Y _07243_/X fanout41/X vssd1 vssd1 vccd1 vccd1 _10580_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06950__B _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__B _11917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ _13350_/CLK hold206/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dfxtp_1
X_12318_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ _12029_/A _12228_/X _12229_/X _12248_/X vssd1 vssd1 vccd1 vccd1 _12249_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12352__B1 _12395_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _09886_/A _06808_/Y _06809_/X vssd1 vssd1 vccd1 vccd1 _06810_/Y sky130_fd_sc_hd__a21oi_1
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__xnor2_1
X_06741_ reg1_val[10] _07213_/A vssd1 vssd1 vccd1 vccd1 _06743_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08859__B1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _09318_/A _09318_/B _09315_/A vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08323__A2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06672_ reg2_val[20] _06712_/B _06707_/B1 _06671_/Y vssd1 vssd1 vccd1 vccd1 _06996_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08411_ _08412_/A _08412_/B vssd1 vssd1 vccd1 vccd1 _08411_/X sky130_fd_sc_hd__or2_1
XANTENNA__11523__S _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09391_ _09387_/X _09390_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _08351_/B _08351_/A vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08087__B2 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07302__A _10466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08273_ _10468_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _08336_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07224_ _07224_/A _07224_/B vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07155_ _07155_/A vssd1 vssd1 vccd1 vccd1 _07155_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07086_ reg1_val[11] reg1_val[12] reg1_val[13] _07229_/C vssd1 vssd1 vccd1 vccd1
+ _07121_/C sky130_fd_sc_hd__or4_4
XANTENNA__08133__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout101 _07068_/Y vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__buf_4
XANTENNA__12343__B1 _12421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13185__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout134 _07072_/Y vssd1 vssd1 vccd1 vccd1 _10233_/B2 sky130_fd_sc_hd__buf_8
Xfanout123 _07167_/Y vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__clkbuf_16
Xfanout145 _07054_/X vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__buf_6
Xfanout156 _12280_/A vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__buf_4
Xfanout178 _12782_/Y vssd1 vssd1 vccd1 vccd1 _13072_/A2 sky130_fd_sc_hd__buf_4
Xfanout189 _07043_/Y vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__buf_12
Xfanout167 _09196_/S vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__clkbuf_8
X_07988_ _07988_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07989_/C sky130_fd_sc_hd__xnor2_1
X_06939_ _11781_/S _09233_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _06939_/X sky130_fd_sc_hd__or3_2
X_09727_ _09723_/X _09726_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _09727_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout47_A _07111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _10613_/A _09658_/B vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__xnor2_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10838__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _06793_/Y _09587_/X _09588_/Y vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__o21ai_1
X_08609_ _09671_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08610_/C sky130_fd_sc_hd__xnor2_1
X_11620_ hold255/A _11620_/B vssd1 vssd1 vccd1 vccd1 _11705_/B sky130_fd_sc_hd__or2_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _06978_/X fanout42/X fanout40/X _07012_/Y vssd1 vssd1 vccd1 vccd1 _11552_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07212__A _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ fanout51/X fanout46/X fanout44/X _11456_/A vssd1 vssd1 vccd1 vccd1 _10503_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11483_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ hold287/A _13220_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10433_ _06754_/B _12394_/A1 _10428_/Y _06752_/Y _10432_/X vssd1 vssd1 vccd1 vccd1
+ _10433_/X sky130_fd_sc_hd__o221a_1
X_13152_ hold311/A _13151_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13152_/X sky130_fd_sc_hd__mux2_1
X_10364_ _10365_/A _10365_/B _10365_/C vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12103_/Y sky130_fd_sc_hd__nor2_1
X_10295_ _07202_/A _06940_/B _10293_/Y _10294_/X vssd1 vssd1 vccd1 vccd1 _10295_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11137__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ _13083_/A _13083_/B vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__xor2_1
XANTENNA__09573__S _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12034_ _12032_/Y _12034_/B vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08002__A1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08553__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ _13193_/A _12935_/B _12859_/X vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__a21o_1
X_12867_ hold320/A hold50/X vssd1 vssd1 vccd1 vccd1 _13160_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11818_ _11910_/A _11818_/B vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13124__A _13134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13062__A1 _11900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _07263_/Y _13078_/B2 hold42/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13248_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09805__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _11749_/A _11917_/C vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06961__A _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10483__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08241__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08960_ _08184_/B _11188_/A _11083_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _08961_/B
+ sky130_fd_sc_hd__o22a_1
X_07911_ _07956_/B _07911_/B vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__and2b_1
X_08891_ _08891_/A _08891_/B _08891_/C vssd1 vssd1 vccd1 vccd1 _08892_/B sky130_fd_sc_hd__and3_1
XANTENNA__09741__A1 _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _08551_/A2 _08274_/B fanout74/X _08551_/B1 vssd1 vssd1 vccd1 vccd1 _07843_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12203__A _12404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__B1 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__B _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__and2_1
X_07773_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06724_ _06799_/A _06801_/B1 _12691_/B _06723_/X vssd1 vssd1 vccd1 vccd1 _07255_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10103__A2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__B1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06655_ _12098_/A _06655_/B _12417_/A _12162_/A vssd1 vssd1 vccd1 vccd1 _06655_/X
+ sky130_fd_sc_hd__and4_1
X_09443_ _07264_/X _07347_/B fanout15/X _09928_/A vssd1 vssd1 vccd1 vccd1 _09444_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09374_ _09374_/A _09374_/B vssd1 vssd1 vccd1 vccd1 _09375_/B sky130_fd_sc_hd__or2_2
XFILLER_0_19_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06586_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06588_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08325_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12800__A1 _10213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ _08256_/A _08256_/B vssd1 vssd1 vccd1 vccd1 _08269_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08187_ _08551_/B1 _10227_/B1 _10463_/A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 _08188_/B
+ sky130_fd_sc_hd__o22a_1
X_07207_ _07207_/A _07207_/B vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__nor2_2
X_07138_ _12193_/A _07138_/B vssd1 vssd1 vccd1 vccd1 _07138_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08232__A1 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A2 _13222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__B2 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ reg1_val[8] _07069_/B vssd1 vssd1 vccd1 vccd1 _07071_/B sky130_fd_sc_hd__xor2_2
X_10080_ _11837_/A fanout35/X fanout32/X fanout60/X vssd1 vssd1 vccd1 vccd1 _10081_/B
+ sky130_fd_sc_hd__o22a_1
X_10982_ _10982_/A _10982_/B vssd1 vssd1 vccd1 vccd1 _10985_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ reg1_val[21] _12773_/A vssd1 vssd1 vccd1 vccd1 _12721_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12652_ reg1_val[7] _12652_/B vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ _12178_/A2 _11542_/X _11809_/D _11889_/A1 vssd1 vssd1 vccd1 vccd1 _11603_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__A1 _07248_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12583_ reg1_val[22] curr_PC[22] _12615_/S vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11534_ _09237_/Y _11529_/Y _11530_/X _11533_/X vssd1 vssd1 vccd1 vccd1 _11534_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__and2_1
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11358__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ hold291/X _13209_/A2 _13203_/X _13204_/B2 vssd1 vssd1 vccd1 vccd1 hold292/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11358__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap109 _10490_/A vssd1 vssd1 vccd1 vccd1 _09114_/B1 sky130_fd_sc_hd__buf_4
X_10416_ _10302_/A _10299_/Y _10301_/B vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08223__A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _11397_/A _11397_/B _11395_/Y vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10030__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08223__B2 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ _13135_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13136_/B sky130_fd_sc_hd__nand2_1
X_10347_ _11900_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12307__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _12065_/A _13072_/A2 _13065_/X vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__o21a_1
X_10278_ _06814_/Y _10277_/Y _12025_/S vssd1 vssd1 vccd1 vccd1 _10280_/B sky130_fd_sc_hd__mux2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08501__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _11689_/B _12271_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__08526__A2 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12958__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__A _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ hold50/X hold320/A vssd1 vssd1 vccd1 vccd1 _13160_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11833__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _09671_/A _09090_/B vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__xor2_1
X_08110_ _06875_/A fanout83/X fanout79/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08111_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07265__A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08041_ _08072_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08041_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08943_ _08944_/B _08944_/A vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10324__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _08874_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08874_/Y sky130_fd_sc_hd__nand2_1
X_07825_ _07826_/A _07825_/B _07825_/C vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07756_ _08566_/A _07756_/B vssd1 vssd1 vccd1 vccd1 _07761_/A sky130_fd_sc_hd__xnor2_2
X_06707_ reg2_val[16] _06712_/B _06707_/B1 _06706_/Y vssd1 vssd1 vccd1 vccd1 _07074_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__11824__A2 wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _09226_/Y _09417_/Y _09418_/X _09419_/Y _09425_/X vssd1 vssd1 vccd1 vccd1
+ _09427_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07788_/B sky130_fd_sc_hd__xnor2_1
X_06638_ reg2_val[24] _06712_/B _06707_/B1 _06637_/Y vssd1 vssd1 vccd1 vccd1 _06975_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13026__A1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ _12415_/A vssd1 vssd1 vccd1 vccd1 _06569_/Y sky130_fd_sc_hd__inv_2
X_09357_ _09110_/A _09110_/B _09108_/Y vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ fanout56/X _10463_/B2 _10228_/A fanout62/X vssd1 vssd1 vccd1 vccd1 _09289_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07256__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _08308_/A _08308_/B vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07697__A _10468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ _08573_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11250_ _11131_/A _09215_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11181_ _12059_/A fanout46/X fanout44/X _11980_/A vssd1 vssd1 vccd1 vccd1 _11182_/B
+ sky130_fd_sc_hd__o22a_1
X_10201_ _12059_/A fanout77/X fanout73/X _11980_/A vssd1 vssd1 vccd1 vccd1 _10202_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06831__A_N _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _09541_/X _09703_/X _09704_/X _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1
+ _10133_/B sky130_fd_sc_hd__a2111oi_1
XANTENNA__07964__B1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__and2_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10965_ _10965_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ reg1_val[16] _12767_/B _12716_/A vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _11776_/A _10896_/B _08731_/X vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__or3b_1
XANTENNA__07495__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12635_ _12634_/A _12631_/Y _12633_/B vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__o21a_2
X_12566_ _12610_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08444__A1 _08619_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _06877_/B _11513_/X _11515_/Y _11612_/A vssd1 vssd1 vccd1 vccd1 _11517_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08444__B2 _09403_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ reg1_val[9] curr_PC[9] _12525_/S vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ curr_PC[16] curr_PC[17] _11448_/C vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _11379_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09944__A1 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ hold283/X _12780_/B _13117_/X _12781_/A vssd1 vssd1 vccd1 vccd1 hold284/A
+ sky130_fd_sc_hd__a22o_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold106/X _13055_/A2 _13053_/B1 hold26/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold107/A sky130_fd_sc_hd__o221a_1
XANTENNA__07707__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08590_ _12785_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08601_/A sky130_fd_sc_hd__nor2_1
X_07610_ _07611_/A _07611_/B vssd1 vssd1 vccd1 vccd1 _07610_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06686__A _06706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07541_ _07541_/A _07541_/B _07541_/C vssd1 vssd1 vccd1 vccd1 _07542_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08132__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07472_ _07666_/A _07666_/B _07471_/C vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__a21oi_1
X_09211_ reg1_val[8] reg1_val[23] _09560_/A vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _09142_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06997__A1 _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__A2 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09073_ _09073_/A _09073_/B vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout3 fanout3/A vssd1 vssd1 vccd1 vccd1 fanout3/X sky130_fd_sc_hd__buf_4
X_08024_ _08566_/A _08024_/B vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__nor2_1
X_08926_ fanout45/X _07197_/Y _08926_/B1 _07814_/B vssd1 vssd1 vccd1 vccd1 _08927_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _08971_/C _08858_/B vssd1 vssd1 vccd1 vccd1 _08857_/Y sky130_fd_sc_hd__xnor2_4
X_07808_ _07808_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08788_ _08767_/B _08767_/C _08776_/X _08787_/B vssd1 vssd1 vccd1 vccd1 _08789_/C
+ sky130_fd_sc_hd__a211o_1
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07850_/B sky130_fd_sc_hd__xnor2_4
X_10750_ _10606_/A _10694_/A _10609_/A vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _10673_/Y _10674_/X _10676_/X _10680_/X vssd1 vssd1 vccd1 vccd1 _10681_/X
+ sky130_fd_sc_hd__o211a_1
X_09409_ _12621_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09409_/X sky130_fd_sc_hd__and2_1
XFILLER_0_118_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ _12420_/A _12420_/B _12420_/C vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__and3_1
XANTENNA__10233__A1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ hold287/A _12349_/X _12350_/Y vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10233__B2 _10233_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11302_ _11189_/A _11189_/B _11192_/A vssd1 vssd1 vccd1 vccd1 _11307_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _06628_/B _06652_/Y _06626_/X vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11233_ _11126_/B _11128_/B _11126_/A vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11165_/B sky130_fd_sc_hd__nand2_1
X_11095_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11095_/Y sky130_fd_sc_hd__nand2_1
X_10115_ _10113_/A _10113_/B _10116_/B vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__o21ba_1
X_10046_ _12202_/A fanout85/X _10466_/A _12059_/A vssd1 vssd1 vccd1 vccd1 _10047_/B
+ sky130_fd_sc_hd__o22a_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11997_ _11998_/A _11998_/B _11998_/C vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__o21ai_1
X_10948_ _10948_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__or2_1
XANTENNA__12997__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10879_ _10880_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12618_ _12619_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ _12549_/A _12549_/B _12549_/C vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11421__B1 _11889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06979__A1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 curr_PC[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__B2 fanout64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12690__B _12691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__B2 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A1 _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06972_ _06973_/A _12621_/A vssd1 vssd1 vccd1 vccd1 _08605_/A sky130_fd_sc_hd__and2_4
X_09760_ _09702_/A _09702_/B _09700_/X vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__a21oi_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _09714_/B _09714_/C vssd1 vssd1 vccd1 vccd1 _08713_/A sky130_fd_sc_hd__nand2_1
X_09691_ _09506_/A _09506_/B _09504_/Y vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__a21o_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ _08650_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07156__A1 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__B2 _06564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout164_A _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08573_ _08573_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__xor2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07524_ _07514_/A _07719_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07524_/X sky130_fd_sc_hd__a21o_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10463__A1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__B2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07455_ _07182_/Y _10326_/A _07218_/Y _07171_/X vssd1 vssd1 vccd1 vccd1 _07456_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06863__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07386_ _07386_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07387_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _09126_/A _09126_/B vssd1 vssd1 vccd1 vccd1 _09125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07975__A _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07631__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _09056_/A _09056_/B vssd1 vssd1 vccd1 vccd1 _09058_/C sky130_fd_sc_hd__or2_1
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09908__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _08007_/A _08007_/B vssd1 vssd1 vccd1 vccd1 _08009_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09908__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout77_A _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__xnor2_2
X_09889_ hold317/A _10158_/A2 _10156_/C _09240_/X vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__a31o_1
X_11920_ _11921_/A _11921_/B vssd1 vssd1 vccd1 vccd1 _11998_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07698__A2 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ _11851_/A vssd1 vssd1 vccd1 vccd1 _11852_/B sky130_fd_sc_hd__inv_2
XFILLER_0_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07162__A4 _07121_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__B1 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _11782_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _11782_/Y sky130_fd_sc_hd__xnor2_1
X_10802_ _09223_/Y _10789_/X _10801_/Y _09153_/Y _10800_/X vssd1 vssd1 vccd1 vccd1
+ _10802_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ fanout74/X _07302_/X fanout13/X _08274_/B vssd1 vssd1 vccd1 vccd1 _10734_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08647__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__A _10933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ _10550_/A _10547_/Y _10549_/B vssd1 vssd1 vccd1 vccd1 _10666_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13383_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__and2_1
X_12403_ _12373_/Y _12374_/X _06943_/Y vssd1 vssd1 vccd1 vccd1 _12403_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _06615_/B _12283_/Y _06613_/X vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13098__S fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ _12320_/B _12265_/B vssd1 vssd1 vccd1 vccd1 _12267_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11216_ _10999_/A _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__o21ba_1
X_12196_ _12310_/A _12196_/B vssd1 vssd1 vccd1 vccd1 _12197_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10914__C1 _12433_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _11889_/A1 _11115_/X _11116_/Y _11146_/X vssd1 vssd1 vccd1 vccd1 _11147_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11078_ _11078_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06948__B _07127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09324__B _11155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12966__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06964__A _06996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09340__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07240_ _06954_/X _06958_/C _06958_/D _07299_/B vssd1 vssd1 vccd1 vccd1 _07251_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07171_ _07169_/Y _07172_/B vssd1 vssd1 vccd1 vccd1 _07171_/X sky130_fd_sc_hd__and2b_2
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__A2 _07146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06585__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__A2 _07944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout281_A _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ _07217_/A _07195_/A vssd1 vssd1 vccd1 vccd1 _06958_/C sky130_fd_sc_hd__or2_4
X_09743_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08326__B1 _10067_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__A1_N _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ instruction[6] _06884_/X _06885_/Y vssd1 vssd1 vccd1 vccd1 _06886_/X sky130_fd_sc_hd__o21a_1
X_09674_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__xnor2_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _12619_/A _08605_/B _08605_/C _07146_/Y _08605_/A vssd1 vssd1 vccd1 vccd1
+ _08626_/B sky130_fd_sc_hd__a32o_1
XANTENNA__07035__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08563_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09826__B1 _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A _10902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _08556_/A _07507_/B vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11633__B1 _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__B2 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08487_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08746_/B sky130_fd_sc_hd__or2_1
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _07448_/B _07516_/A _07448_/A vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _07369_/A _07369_/B vssd1 vssd1 vccd1 vccd1 _07453_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07065__B1 _07093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ _09109_/A _09109_/B vssd1 vssd1 vccd1 vccd1 _09108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ fanout62/X fanout27/X fanout25/X fanout61/X vssd1 vssd1 vccd1 vccd1 _10381_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09039_ _08805_/B _08805_/C _09544_/A _08918_/X _09706_/A vssd1 vssd1 vccd1 vccd1
+ _09042_/A sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12050_ curr_PC[24] _12050_/B vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__or2_1
X_11001_ _11001_/A _11110_/A vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12361__A1 _08857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12952_ _12978_/A _12952_/B vssd1 vssd1 vccd1 vccd1 _13274_/D sky130_fd_sc_hd__and2_1
XANTENNA__09144__B _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _11904_/B _11903_/B vssd1 vssd1 vccd1 vccd1 _11983_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10675__A1 _12394_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12883_ hold271/X hold104/X vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07540__A1 _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _12404_/B _11834_/B vssd1 vssd1 vccd1 vccd1 _11836_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09817__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11765_/A vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__inv_2
XFILLER_0_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _12202_/B fanout35/X fanout33/X _12202_/A vssd1 vssd1 vccd1 vccd1 _10717_/B
+ sky130_fd_sc_hd__o22a_1
X_11696_ _06683_/C _11695_/X _09226_/Y vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _10403_/X _10527_/X _10528_/X vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ _13375_/CLK _13366_/D vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__dfxtp_1
X_10578_ _10578_/A _10578_/B vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06950__C _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13297_ _13297_/CLK hold201/X vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__dfxtp_1
X_12317_ _07301_/Y _11917_/C _12258_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _12319_/B
+ sky130_fd_sc_hd__a31o_1
X_12248_ _06924_/Y _12235_/X _12242_/Y _12247_/X vssd1 vssd1 vccd1 vccd1 _12248_/X
+ sky130_fd_sc_hd__a211o_1
X_12179_ _12431_/A2 _09235_/X _12179_/S vssd1 vssd1 vccd1 vccd1 _12179_/X sky130_fd_sc_hd__mux2_1
X_06740_ _06799_/A _06801_/B1 _12673_/B _06739_/X vssd1 vssd1 vccd1 vccd1 _07213_/A
+ sky130_fd_sc_hd__a31o_4
X_06671_ _06706_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08859__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _08410_/A _08410_/B vssd1 vssd1 vccd1 vccd1 _08412_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13065__C1 _13016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09390_ _09388_/X _09389_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12812__C1 _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13080__A2 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ _08341_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08087__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07302__B _10466_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _08591_/B1 _08400_/B fanout82/X _08619_/B1 vssd1 vssd1 vccd1 vccd1 _08273_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07223_ _07084_/A _07084_/B _07224_/B vssd1 vssd1 vccd1 vccd1 _07223_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11918__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A _11169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ _07150_/A _07150_/B _12065_/A vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07085_ reg1_val[8] reg1_val[9] reg1_val[10] _07085_/D vssd1 vssd1 vccd1 vccd1 _07229_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__A2 _11188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout113 _07201_/X vssd1 vssd1 vccd1 vccd1 _08551_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout135 _08445_/A vssd1 vssd1 vccd1 vccd1 _10230_/A sky130_fd_sc_hd__clkbuf_16
Xfanout124 _07210_/A vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__clkbuf_16
Xfanout146 _08590_/B vssd1 vssd1 vccd1 vccd1 _08594_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout179 _12839_/B vssd1 vssd1 vccd1 vccd1 _12841_/B sky130_fd_sc_hd__buf_4
Xfanout168 _09153_/Y vssd1 vssd1 vccd1 vccd1 _09196_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__09245__A _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _12280_/A vssd1 vssd1 vccd1 vccd1 _11776_/A sky130_fd_sc_hd__buf_4
X_07987_ _07986_/A _07986_/B _07986_/C vssd1 vssd1 vccd1 vccd1 _07989_/B sky130_fd_sc_hd__a21oi_1
X_06938_ _11781_/S _09233_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__nor3_2
X_09726_ _09724_/X _09725_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06869_ _12285_/A _06868_/Y _06851_/Y vssd1 vssd1 vccd1 vccd1 _12335_/B sky130_fd_sc_hd__o21ai_1
X_09657_ fanout57/X fanout85/X _10466_/A fanout62/X vssd1 vssd1 vccd1 vccd1 _09658_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _06793_/Y _09587_/X _11612_/A vssd1 vssd1 vccd1 vccd1 _09588_/Y sky130_fd_sc_hd__a21oi_1
X_08608_ _07010_/Y _07146_/Y _07153_/Y _07018_/X vssd1 vssd1 vccd1 vccd1 _08609_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08559_/B _08559_/A vssd1 vssd1 vccd1 vccd1 _08542_/C sky130_fd_sc_hd__and2b_1
X_11550_ _11663_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__nand2_1
X_10501_ _10501_/A _10501_/B vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout6_A fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _11481_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__nand2_1
X_13220_ _13220_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ _07195_/A _06940_/B _10430_/Y _10431_/X vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08324__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13151_/A _13151_/B vssd1 vssd1 vccd1 vccd1 _13151_/Y sky130_fd_sc_hd__xnor2_1
X_10363_ _10491_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10365_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10042__C1 _11645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10593__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _12035_/A _12032_/Y _12034_/B vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__o21a_1
X_13082_ _13109_/A hold274/X vssd1 vssd1 vccd1 vccd1 _13338_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10294_ hold313/A _12349_/A _10558_/C _12393_/B1 vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__a31o_1
X_12033_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09735__C1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _12859_/X _12935_/B vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ hold281/X hold139/X vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__nand2b_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11817_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11818_/B sky130_fd_sc_hd__or2_1
XANTENNA__06945__C _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07403__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13062__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ hold41/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__or2_1
XFILLER_0_56_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09266__B2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11748_ _11748_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _11679_/A _11679_/B _11679_/C vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10820__A1 _10942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__S _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12022__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13349_ _13363_/CLK _13349_/D vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08241__A2 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10336__B1 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07910_ _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__xnor2_1
X_08890_ _08891_/A _08891_/B _08891_/C vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07284__S _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _10468_/A _07841_/B vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07752__A1 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__B2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _11361_/A _07772_/B vssd1 vssd1 vccd1 vccd1 _07774_/B sky130_fd_sc_hd__xnor2_1
X_06723_ reg2_val[13] _06794_/B vssd1 vssd1 vccd1 vccd1 _06723_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09511_ _09827_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07504__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06654_ _12179_/S _06654_/B vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__or2_2
X_09442_ _09363_/A _09363_/B _09364_/Y vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__o21ai_4
X_06585_ instruction[15] _06575_/X _06584_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__o211a_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _09371_/B _09034_/Y _09371_/D _09372_/X _09143_/Y vssd1 vssd1 vccd1 vccd1
+ _09374_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout244_A _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ _09941_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08328_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11603__A3 _11809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__A2 _13072_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ _08249_/A _08249_/B _08251_/B _08313_/A vssd1 vssd1 vccd1 vccd1 _08269_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08186_/X sky130_fd_sc_hd__and2b_1
X_07206_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07207_/B sky130_fd_sc_hd__nor2_1
X_07137_ _07138_/B _12132_/A vssd1 vssd1 vccd1 vccd1 _07137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__A2 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _07068_/A _07068_/B vssd1 vssd1 vccd1 vccd1 _07068_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10981_ _10824_/A _10824_/B _10825_/Y vssd1 vssd1 vccd1 vccd1 _10987_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09703__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _09037_/B _09706_/X _09707_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _09710_/B
+ sky130_fd_sc_hd__o211a_2
X_12720_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
XFILLER_0_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ reg1_val[7] _12652_/B vssd1 vssd1 vccd1 vccd1 _12651_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08319__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ _12178_/A2 _11542_/X _11809_/D vssd1 vssd1 vccd1 vccd1 _11602_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12783__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ _12588_/B _12582_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12252__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11533_ _09155_/S _11022_/X _11034_/X _09222_/Y _11532_/Y vssd1 vssd1 vccd1 vccd1
+ _11533_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10802__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ _11740_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11358__A2 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13203_ hold269/X _13202_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _10414_/A _10414_/B _10414_/Y _11612_/A vssd1 vssd1 vccd1 vccd1 _10415_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11395_ _11282_/Y _11285_/B _11290_/A vssd1 vssd1 vccd1 vccd1 _11395_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08223__A2 _08274_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13134_ _13134_/A hold306/X vssd1 vssd1 vccd1 vccd1 _13349_/D sky130_fd_sc_hd__and2_1
X_10346_ _11456_/A fanout46/X fanout44/X _11386_/A vssd1 vssd1 vccd1 vccd1 _10347_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12307__A1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07431__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__B2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ hold92/X _13071_/A2 _13071_/B1 hold126/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ _13065_/X sky130_fd_sc_hd__o221a_1
X_10277_ _06763_/A _10141_/Y _06765_/B vssd1 vssd1 vccd1 vccd1 _10277_/Y sky130_fd_sc_hd__a21oi_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12016_ _12016_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12271_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13287_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12918_ _13155_/A _13156_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__B _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ hold68/X hold287/A vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11046__A1 _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__A _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06972__A _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__B _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12794__A1 _07114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10557__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08942_ _08842_/A _08841_/Y _08837_/Y vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08873_ _08874_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08873_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout194_A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _09671_/A _07824_/B vssd1 vssd1 vccd1 vccd1 _07825_/C sky130_fd_sc_hd__xor2_1
X_07755_ _06875_/A fanout62/X fanout60/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _07756_/B
+ sky130_fd_sc_hd__o22a_1
X_06706_ _06706_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _06706_/Y sky130_fd_sc_hd__nor2_1
X_07686_ _07768_/A _07768_/B _07682_/X vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06637_ _06706_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _06637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _09586_/A _09595_/B _09412_/X _12171_/A _09424_/X vssd1 vssd1 vccd1 vccd1
+ _09425_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06568_ reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__inv_6
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _09356_/A _09356_/B vssd1 vssd1 vccd1 vccd1 _09361_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07978__A _09630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09287_ _10231_/A _09287_/B vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08989__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ _08305_/A _08305_/B _08306_/X vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _08572_/A2 _08521_/A2 _08926_/B1 _08594_/A2 vssd1 vssd1 vccd1 vccd1 _08239_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__or2_1
X_08169_ _08071_/A _08070_/B _08070_/C vssd1 vssd1 vccd1 vccd1 _08170_/B sky130_fd_sc_hd__o21a_1
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12124__A _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _09855_/X _09993_/X _09994_/X vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07964__A1 _08533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__B2 _08507_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _07053_/X fanout7/X _10061_/Y _09938_/A vssd1 vssd1 vccd1 vccd1 _10064_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10964_ _10964_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__and2_1
XFILLER_0_97_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12703_/A _12703_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xor2_4
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ _11863_/A _08731_/X _10896_/B vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__a21bo_1
X_12634_ _12634_/A _12634_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ _12610_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _12575_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08444__A2 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ _11513_/X _11515_/Y _06877_/B vssd1 vssd1 vccd1 vccd1 _11516_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12496_ _12502_/B _12496_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XFILLER_0_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11447_ curr_PC[16] _11448_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11378_ _12065_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09944__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13117_ hold313/A _13116_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_10329_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10458_/A sky130_fd_sc_hd__or2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07128__A _09725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _07180_/C _13052_/A2 hold171/X vssd1 vssd1 vccd1 vccd1 _13322_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__07707__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__B2 _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06915__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__A2 _10222_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__A2 _09243_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06686__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _08476_/A _07539_/B _09766_/A vssd1 vssd1 vccd1 vccd1 _07542_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08132__B2 _08553_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__A1 _08553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07471_ _07666_/A _07666_/B _07471_/C vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__and3_1
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ reg1_val[9] reg1_val[22] _09560_/A vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ _09141_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ _09073_/A _09073_/B vssd1 vssd1 vccd1 vccd1 _09072_/Y sky130_fd_sc_hd__nor2_1
X_08023_ _06875_/A _09659_/B2 fanout98/X _08551_/B2 vssd1 vssd1 vccd1 vccd1 _08024_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10952__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout4 fanout5/X vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__buf_6
XANTENNA_fanout207_A _08476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08941_/B _08853_/B _08866_/B _08867_/B _08867_/A vssd1 vssd1 vccd1 vccd1
+ _08938_/B sky130_fd_sc_hd__a32o_1
X_08856_ _06850_/B _06851_/B _07300_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _08858_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08787_ _08787_/A _08787_/B vssd1 vssd1 vccd1 vccd1 _08789_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07738_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07850_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__A1 _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ _08594_/A2 fanout98/X fanout83/X _08572_/A2 vssd1 vssd1 vccd1 vccd1 _07670_/B
+ sky130_fd_sc_hd__o22a_2
X_10680_ _07213_/A _06940_/B _10678_/Y _10679_/X vssd1 vssd1 vccd1 vccd1 _10680_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout22_A _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _09408_/A vssd1 vssd1 vccd1 vccd1 _09408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07882__B1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ fanout27/X _11188_/A _11083_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _09340_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ hold287/A _12349_/X _09239_/Y vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10233__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ _11186_/A _11186_/B _11193_/Y vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11958__A _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ _12280_/A _12280_/C _12280_/B vssd1 vssd1 vccd1 vccd1 _12281_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _11230_/X _11232_/B vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11305_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _09974_/A _09974_/B _09972_/Y vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__a21oi_4
X_11094_ _10967_/A _10967_/B _10965_/A vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__a21o_1
X_10045_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
X_11996_ _12073_/B _11996_/B vssd1 vssd1 vccd1 vccd1 _11998_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09311__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ _10948_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12617_/A _12617_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
X_10878_ _10878_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12029__A _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ _12549_/A _12549_/B _12549_/C vssd1 vssd1 vccd1 vccd1 _12559_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12479_ _12488_/A _12479_/B vssd1 vssd1 vccd1 vccd1 _12481_/C sky130_fd_sc_hd__nand2_1
XANTENNA_2 curr_PC[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06979__A2 fanout67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11724__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08242__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10932__B1 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _07026_/B _06971_/B vssd1 vssd1 vccd1 vccd1 _06971_/Y sky130_fd_sc_hd__xnor2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _09714_/C sky130_fd_sc_hd__xor2_1
X_09690_ _09456_/A _09456_/B _09459_/A vssd1 vssd1 vccd1 vccd1 _09695_/A sky130_fd_sc_hd__o21ai_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _09403_/S _08641_/A2 _09324_/A _08649_/B vssd1 vssd1 vccd1 vccd1 _08642_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07156__A2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A0 _09219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ _09403_/S _08572_/A2 _08619_/B1 _08590_/B vssd1 vssd1 vccd1 vccd1 _08573_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _07522_/B _07522_/C _07522_/A vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10463__A2 fanout11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06821__A_N _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ _07454_/A _07454_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07385_ _07385_/A _07385_/B _07420_/A vssd1 vssd1 vccd1 vccd1 _07386_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09124_ _09124_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _09126_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09054_/B _09055_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09908__A2 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A _10286_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08006_ _08078_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__or2_1
XANTENNA__11176__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09959_/B sky130_fd_sc_hd__xnor2_1
X_08908_ _08909_/B _08909_/A vssd1 vssd1 vccd1 vccd1 _08908_/Y sky130_fd_sc_hd__nand2b_1
X_09888_ _10158_/A2 _10156_/C hold317/A vssd1 vssd1 vccd1 vccd1 _09888_/Y sky130_fd_sc_hd__a21oi_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ fanout62/X _10233_/B2 _10233_/A1 fanout60/X vssd1 vssd1 vccd1 vccd1 _08840_/B
+ sky130_fd_sc_hd__o22a_1
X_11850_ _11850_/A _11850_/B _11850_/C vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__and3_1
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ _11779_/X _11780_/X _11781_/S vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ _11131_/A _09880_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__08647__A2 _07128_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _10942_/A _10732_/B vssd1 vssd1 vccd1 vccd1 _10738_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07231__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10666_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ _11557_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__xnor2_2
X_13382_ instruction[6] vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
X_12402_ _08971_/C _11446_/B _12401_/X _12504_/S vssd1 vssd1 vccd1 vccd1 dest_val[30]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12791__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__A _11052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _12333_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12320_/A _12263_/C _12263_/A vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11215_ _11213_/Y _11215_/B vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__nand2b_2
X_12195_ fanout14/X fanout12/X fanout6/X fanout22/X vssd1 vssd1 vccd1 vccd1 _12196_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08032__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11117_/Y _11118_/X _11123_/X _11145_/X vssd1 vssd1 vccd1 vccd1 _11146_/X
+ sky130_fd_sc_hd__o211a_1
X_11077_ _11077_/A _11077_/B vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__xnor2_1
X_10028_ _10026_/Y _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11890__A1 _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08099__A0 _09795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06964__B _06964_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ _07150_/A _11978_/Y _11977_/X vssd1 vssd1 vccd1 vccd1 _12056_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08237__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12982__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07170_ _11168_/A _07180_/C vssd1 vssd1 vccd1 vccd1 _07172_/B sky130_fd_sc_hd__nand2_2
XANTENNA__06980__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08023__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09742_/X sky130_fd_sc_hd__or2_1
X_06954_ _07113_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06954_/X sky130_fd_sc_hd__or2_1
XANTENNA__08326__B2 _08641_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__A1 _08649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06885_ instruction[6] _06943_/B _09233_/A vssd1 vssd1 vccd1 vccd1 _06885_/Y sky130_fd_sc_hd__a21oi_1
X_09673_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__xor2_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08632_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_119_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09826__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A1 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _08533_/B fanout83/X fanout79/X _08507_/A2 vssd1 vssd1 vccd1 vccd1 _07507_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08486_ _08678_/B vssd1 vssd1 vccd1 vccd1 _08486_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13374_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07437_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ _09787_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13199__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09107_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09109_/B sky130_fd_sc_hd__xnor2_2
X_07299_ _08971_/B _07299_/B vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ _09038_/A _09038_/B _12383_/A _12420_/C vssd1 vssd1 vccd1 vccd1 _10310_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08014__B1 _10463_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _10763_/X _10884_/X _10886_/B vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08565__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ hold321/X _13158_/A2 fanout3/X _13108_/B2 vssd1 vssd1 vccd1 vccd1 _12952_/B
+ sky130_fd_sc_hd__a22o_1
X_11902_ _12065_/A _11902_/B vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__xnor2_1
X_12882_ hold104/X hold271/X vssd1 vssd1 vccd1 vccd1 _12882_/X sky130_fd_sc_hd__and2b_1
X_11833_ _11980_/A fanout9/X fanout4/X fanout57/X vssd1 vssd1 vccd1 vccd1 _11834_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07540__A2 _07539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06784__B _07145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__B2 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__A1 _07264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__and3_1
XFILLER_0_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10726_/A sky130_fd_sc_hd__xnor2_1
X_11695_ _06840_/Y _11694_/Y _11781_/S vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10646_ _10646_/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__nand2_4
XANTENNA__09587__S _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ _13375_/CLK _13365_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
X_10577_ _10577_/A vssd1 vssd1 vccd1 vccd1 _10578_/B sky130_fd_sc_hd__inv_2
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13350_/CLK _13296_/D vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__dfxtp_1
X_12316_ _12366_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12319_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06950__D _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12247_ _09237_/Y _12237_/X _12238_/Y _12246_/X vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _13300_/Q _12178_/A2 _12236_/B _12177_/Y _11242_/A vssd1 vssd1 vccd1 vccd1
+ _12183_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ _11958_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__A2 _07593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ instruction[30] _06699_/B vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__and2_4
XFILLER_0_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12696__B _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__A1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07819__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _08337_/A _08337_/B _08339_/Y vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ _08271_/A _08271_/B vssd1 vssd1 vccd1 vccd1 _08305_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07224_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11918__A2 _11988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07153_ _10286_/S _07153_/B vssd1 vssd1 vccd1 vccd1 _07153_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ _07084_/A _07084_/B vssd1 vssd1 vccd1 vccd1 _07224_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 _10463_/A1 vssd1 vssd1 vccd1 vccd1 _10228_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11551__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _10736_/A vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__buf_12
Xfanout147 _07048_/Y vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__buf_6
Xfanout125 _07163_/X vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__buf_12
Xfanout114 _07197_/Y vssd1 vssd1 vccd1 vccd1 _08521_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout158 _06943_/Y vssd1 vssd1 vccd1 vccd1 _12280_/A sky130_fd_sc_hd__buf_4
Xfanout169 _09155_/S vssd1 vssd1 vccd1 vccd1 _09180_/S sky130_fd_sc_hd__clkbuf_8
X_07986_ _07986_/A _07986_/B _07986_/C vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__and3_1
X_06937_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09229_/B sky130_fd_sc_hd__nand2b_4
XANTENNA__07046__A _09668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _09393_/X _09403_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ _09656_/A _09656_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__xnor2_2
X_06868_ _06858_/A _06867_/X _06852_/Y vssd1 vssd1 vccd1 vccd1 _06868_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _08648_/A _08607_/B _08607_/C vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__or3_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _06799_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _06799_/X sky130_fd_sc_hd__and2_1
X_09587_ _06804_/X _09586_/Y _12025_/S vssd1 vssd1 vccd1 vccd1 _09587_/X sky130_fd_sc_hd__mux2_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08469_ _08594_/A2 _08553_/B1 _09468_/B2 _08572_/A2 vssd1 vssd1 vccd1 vccd1 _08470_/B
+ sky130_fd_sc_hd__o22a_1
X_10500_ _10500_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10501_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ _11479_/B _11480_/B vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09200__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10431_ hold283/A _12349_/A _10429_/X _12393_/B1 vssd1 vssd1 vccd1 vccd1 _10431_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ _13150_/A _13150_/B vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10593__A1 _11980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ _11169_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10042__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ _12349_/A _10558_/C hold313/A vssd1 vssd1 vccd1 vccd1 _10293_/Y sky130_fd_sc_hd__a21oi_1
X_13081_ _13108_/B2 _13079_/Y _13080_/X _13222_/A2 _13338_/Q vssd1 vssd1 vccd1 vccd1
+ hold274/A sky130_fd_sc_hd__a32o_1
X_12101_ _12339_/A1 _08792_/A _08792_/B _11946_/A vssd1 vssd1 vccd1 vccd1 _12101_/X
+ sky130_fd_sc_hd__a31o_1
X_12032_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06779__B _07097_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ hold289/X hold108/X vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ hold139/X hold281/X vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11816_ _11817_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__nand2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12796_ _07101_/Y _13078_/B2 hold22/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13247_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__A2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ _11661_/A _11661_/B _11649_/A vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__o21a_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11678_ _11679_/A _11679_/B _11679_/C vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06961__C _11446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ _10509_/A _10509_/C _10509_/B vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12022__A1 _12280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08226__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ _13372_/CLK _13348_/D vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _13287_/CLK hold224/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06689__B _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A1 _10228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__B2 _10463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _08926_/B1 _08400_/B fanout82/X _08521_/A2 vssd1 vssd1 vccd1 vccd1 _07841_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07752__A2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _08553_/A2 fanout32/X _08551_/B1 _08184_/B vssd1 vssd1 vccd1 vccd1 _07772_/B
+ sky130_fd_sc_hd__o22a_1
X_06722_ _06879_/B vssd1 vssd1 vccd1 vccd1 _06722_/Y sky130_fd_sc_hd__inv_2
X_09510_ _07814_/B _10859_/A _10327_/B2 fanout45/X vssd1 vssd1 vccd1 vccd1 _09511_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07504__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06653_ reg1_val[26] _07026_/B vssd1 vssd1 vccd1 vccd1 _06654_/B sky130_fd_sc_hd__and2b_1
X_09441_ _09368_/A _09368_/B _09366_/X vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__a21oi_4
X_06584_ instruction[22] _06922_/B vssd1 vssd1 vccd1 vccd1 _06584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09257__A2 _12525_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09372_ _09145_/B _09145_/A _09033_/B _09033_/A vssd1 vssd1 vccd1 vccd1 _09372_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08323_ _08619_/A2 _08521_/A2 _08926_/B1 _08619_/B2 vssd1 vssd1 vccd1 vccd1 _08324_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout237_A _06973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08313_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08185_ _10081_/A _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__mux2_1
X_07205_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07207_/A sky130_fd_sc_hd__and2_1
X_07136_ _07135_/A _07135_/B _07135_/C vssd1 vssd1 vccd1 vccd1 _12132_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__B2 _07077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A1 _07968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _07067_/A _07068_/B vssd1 vssd1 vccd1 vccd1 _07067_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__A1 _10859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B2 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _09996_/A _10128_/A _09372_/X _09143_/Y vssd1 vssd1 vccd1 vccd1 _09708_/X
+ sky130_fd_sc_hd__or4bb_1
X_07969_ _07970_/B _07970_/C _08566_/A vssd1 vssd1 vccd1 vccd1 _07973_/A sky130_fd_sc_hd__a21oi_1
X_10980_ _10874_/A _10874_/B _10872_/Y vssd1 vssd1 vccd1 vccd1 _10989_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout52_A _07052_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _09480_/B _09483_/B _09480_/A vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__o21bai_2
X_12650_ _12649_/A _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__o21ba_2
X_11601_ _11767_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11809_/D sky130_fd_sc_hd__xor2_4
XANTENNA__12252__A1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12788__C1 _13109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12588_/A _12577_/Y _12573_/A vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12252__B2 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _12395_/A1 _11531_/X _06698_/B vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ fanout29/X _07593_/Y _08857_/Y fanout31/X vssd1 vssd1 vccd1 vccd1 _11464_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13202_/Y sky130_fd_sc_hd__xnor2_1
X_10414_ _10414_/A _10414_/B vssd1 vssd1 vccd1 vccd1 _10414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ _11295_/A _11295_/B _11298_/A vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__o21ai_2
X_13133_ hold305/X _13209_/A2 _13132_/X _13143_/B2 vssd1 vssd1 vccd1 vccd1 hold306/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10566__B2 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07431__A1 _10327_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12307__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07431__B2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13064_ _07148_/C _13072_/A2 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o21a_1
X_10276_ _10315_/A _10276_/B _10276_/C vssd1 vssd1 vccd1 vccd1 _10276_/X sky130_fd_sc_hd__or3_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _11853_/Y _12016_/B _12013_/X vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__a21bo_1
X_12917_ hold74/X hold297/X vssd1 vssd1 vccd1 vccd1 _13155_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07498__A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__B2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12848_ wire8/A _13072_/A2 hold63/X _13236_/A vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__o211a_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12779_ _12782_/A hold198/X vssd1 vssd1 vccd1 vccd1 _12780_/C sky130_fd_sc_hd__nor2_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06972__B _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12794__A2 _13078_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12990__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09990_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06776__A3 _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _08847_/X _08941_/B vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _12310_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08874_/B sky130_fd_sc_hd__nand2_1
X_07823_ _09297_/B2 fanout50/X _09659_/B2 _09297_/A1 vssd1 vssd1 vccd1 vccd1 _07824_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _07765_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07754_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06705_ instruction[0] instruction[1] instruction[2] instruction[26] pred_val vssd1
+ vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__o311a_4
X_07685_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__xnor2_2
X_06636_ instruction[34] _06657_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__and2_4
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09424_ reg1_val[1] _07129_/A _11966_/B _09423_/X vssd1 vssd1 vccd1 vccd1 _09424_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06567_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06567_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _09128_/A _09127_/B _09125_/Y vssd1 vssd1 vccd1 vccd1 _09365_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ fanout55/X _08590_/B _09648_/A fanout67/X vssd1 vssd1 vccd1 vccd1 _09287_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08989__B2 _12785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__A1 _09324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _08314_/B _08314_/A vssd1 vssd1 vccd1 vccd1 _08306_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _08445_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08168_ _08776_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _08168_/X sky130_fd_sc_hd__or2_1
X_08099_ _09795_/A _08144_/B _08144_/A vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__mux2_2
X_07119_ _09827_/A _07119_/B vssd1 vssd1 vccd1 vccd1 _07142_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ _09546_/X _09547_/X _10129_/C vssd1 vssd1 vccd1 vccd1 _10130_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07964__A2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _10061_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10061_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07177__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _10964_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10965_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07234__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12702_ _12703_/A _12703_/B vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _10812_/X _11041_/B _10893_/Y vssd1 vssd1 vccd1 vccd1 _10894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12225__A1 _12415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06792__B _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12633_ _12631_/Y _12633_/B vssd1 vssd1 vccd1 vccd1 _12634_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_108_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ reg1_val[19] curr_PC[19] _12615_/S vssd1 vssd1 vccd1 vccd1 _12566_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _11781_/S _11515_/B vssd1 vssd1 vccd1 vccd1 _11515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ _12495_/A _12495_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09929__B1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ _11446_/A _11446_/B vssd1 vssd1 vccd1 vccd1 _11446_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _06978_/X _07151_/A _07155_/A _07012_/Y vssd1 vssd1 vccd1 vccd1 _11378_/B
+ sky130_fd_sc_hd__a22o_1
X_13116_ _13116_/A _13116_/B vssd1 vssd1 vccd1 vccd1 _13116_/Y sky130_fd_sc_hd__xnor2_1
X_10328_ _12131_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10330_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ hold170/X _13055_/A2 _13053_/B1 hold106/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold171/A sky130_fd_sc_hd__o221a_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10261_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07707__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08132__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _09827_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _07471_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10227__B1 _10227_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09093__B1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ _09141_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__and2_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09071_ _10230_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09073_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ _08020_/A _08020_/B _08066_/A vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout5 fanout5/A vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07319__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08924_ _08907_/A _08907_/B _08908_/Y vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__o21ai_4
X_08855_ _09671_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08865_/A sky130_fd_sc_hd__xnor2_2
X_07806_ _07806_/A _07806_/B vssd1 vssd1 vccd1 vccd1 _07856_/A sky130_fd_sc_hd__xnor2_4
X_08786_ _08786_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _08787_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08659__A0 _08650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07737_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07668_ _08445_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07331__B1 _08551_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06619_ _06617_/Y _06707_/B1 _06712_/B reg2_val[30] vssd1 vssd1 vccd1 vccd1 _08971_/C
+ sky130_fd_sc_hd__a2bb2o_4
X_09407_ _09392_/X _09406_/X _11131_/A vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__mux2_2
XANTENNA__07882__B2 _09467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__A1 _09675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07600_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10218__B1 _07250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _09827_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09084__B1 fanout73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _11300_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ _09268_/B _09269_/B vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _12280_/A _12280_/B _12280_/C vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__or3_1
X_11231_ _11231_/A curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _12310_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__xnor2_1
X_10113_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__or2_2
X_11093_ _10948_/A _10948_/B _10968_/A vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12789__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ _10042_/X _10044_/B vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09444__A _09930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ _11995_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _11996_/B sky130_fd_sc_hd__and2_1
XANTENNA__09311__A1 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ _10946_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10948_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12997__A2 _13204_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07899__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__B2 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10877_ _10878_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10877_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12616_ _12616_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _12610_/A _12547_/B vssd1 vssd1 vccd1 vccd1 _12549_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11421__A2 _11451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ _12647_/B _12478_/B vssd1 vssd1 vccd1 vccd1 _12479_/B sky130_fd_sc_hd__or2_1
XANTENNA_3 dest_pred_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ _11338_/A _11335_/Y _11337_/B vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__B2 _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A1 _11749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06970_ _07026_/B _06971_/B vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__xor2_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08640_ _08648_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10160__A2 _06940_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _08600_/A _08600_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand3_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10448__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__B1 _10233_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _07522_/A _07522_/B _07522_/C vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07602__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__and2_1
XANTENNA__11124__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11948__B1 _12025_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ _07385_/B _07420_/A _07385_/A vssd1 vssd1 vccd1 vccd1 _07386_/A sky130_fd_sc_hd__o21a_1
X_09123_ _09123_/A _09123_/B vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _09055_/B _09054_/B vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08005_ _08556_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08078_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11176__B2 _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__A1 _07031_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10923__A1 _09223_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__B2 _09196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09956_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__and2_1
X_09887_ hold271/A hold322/A hold265/A _13338_/Q vssd1 vssd1 vccd1 vccd1 _10156_/C
+ sky130_fd_sc_hd__or4_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__xor2_2
X_08769_ _08769_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__nand2_2
X_11780_ _06683_/C _11694_/Y _11711_/S vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__a21o_1
X_10800_ _10800_/A _10800_/B _10800_/C vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__and3_1
XFILLER_0_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ fanout82/X fanout12/X fanout6/X _08400_/B vssd1 vssd1 vccd1 vccd1 _10732_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09203__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _12375_/Y _12376_/X _12379_/X _12380_/Y _12400_/X vssd1 vssd1 vccd1 vccd1
+ _12401_/X sky130_fd_sc_hd__a221o_1
X_10662_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10593_ _11980_/A fanout27/X fanout25/X fanout56/X vssd1 vssd1 vccd1 vccd1 _10594_/B
+ sky130_fd_sc_hd__o22a_1
X_13381_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ _06943_/Y _12374_/C _12330_/Y _09148_/Y vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__o31a_1
X_12263_ _12263_/A _12320_/A _12263_/C vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__nor3_1
X_11214_ _11214_/A _11214_/B _11214_/C vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__nand3_1
X_12194_ _12255_/A _12194_/B vssd1 vssd1 vccd1 vccd1 _12199_/A sky130_fd_sc_hd__and2_1
XANTENNA__08032__A1 _09468_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__B2 _08591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _09223_/Y _11132_/Y _11133_/X _11144_/X vssd1 vssd1 vccd1 vccd1 _11145_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06798__A _12621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11077_/B _11077_/A vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__and2b_1
X_10027_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__nand2_1
XANTENNA_max_cap115_A _07179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11890__A2 _11446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11978_ _12065_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _11978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _10812_/B _11041_/B _11776_/A vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13276__CLK _13297_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09220__B1 _11958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09771__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A1 _07402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__B1 _12107_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06953_ _07113_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06963_/A sky130_fd_sc_hd__nor2_4
X_09741_ _12025_/S _09595_/A _09740_/X _09739_/X vssd1 vssd1 vccd1 vccd1 _09743_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08326__A2 _10585_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06884_ _06656_/X _06884_/B _06884_/C _06884_/D vssd1 vssd1 vccd1 vccd1 _06884_/X
+ sky130_fd_sc_hd__and4b_1
X_09672_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09672_/Y sky130_fd_sc_hd__nor2_1
X_08623_ _07018_/X _07128_/Y _07153_/Y _07010_/Y vssd1 vssd1 vccd1 vccd1 _08624_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout267_A _06591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08554_ _08624_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09826__A2 _11083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _09668_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07332__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ _08459_/B _08459_/C _08459_/A vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07436_ _07436_/A _07436_/B vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10693__A _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ fanout85/X fanout75/X fanout71/X _10466_/A vssd1 vssd1 vccd1 vccd1 _07368_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09106_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09107_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13138__A2 _13186_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ _07299_/B _08971_/D _08971_/B vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__a21oi_4
X_09037_ _09371_/B _09037_/B vssd1 vssd1 vccd1 vccd1 _12420_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08014__A1 _08926_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__B2 _08521_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08565__A2 _07101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07507__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__B wire8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _10233_/A1 _12257_/A fanout13/X _07072_/Y vssd1 vssd1 vccd1 vccd1 _09940_/B
+ sky130_fd_sc_hd__o22a_2
X_12950_ _12950_/A _13224_/B vssd1 vssd1 vccd1 vccd1 fanout3/A sky130_fd_sc_hd__or2_1
X_11901_ _07155_/Y fanout11/X fanout6/X _07151_/Y vssd1 vssd1 vccd1 vccd1 _11902_/B
+ sky130_fd_sc_hd__o22a_1
X_12881_ _12879_/X _12881_/B vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__nand2b_1
X_11832_ _11740_/A _11740_/B _11745_/A vssd1 vssd1 vccd1 vccd1 _11836_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13074__A1 _12310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07242__A _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10715_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ _11611_/A _11609_/B _11626_/S vssd1 vssd1 vccd1 vccd1 _11694_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10645_ _10645_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__nand2_1
X_13364_ _13364_/CLK _13364_/D vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10576_ _10933_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__xor2_1
X_12315_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__or2_1
XANTENNA__09450__B1 _09450_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _13352_/CLK _13295_/D vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12337__B1 _09226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12246_ _09222_/Y _09875_/Y _09881_/X _09155_/S _12245_/Y vssd1 vssd1 vccd1 vccd1
+ _12246_/X sky130_fd_sc_hd__a221o_1
X_12177_ _12347_/B _12236_/B _13300_/Q vssd1 vssd1 vccd1 vccd1 _12177_/Y sky130_fd_sc_hd__a21oi_1
X_11128_ _11128_/A _11128_/B vssd1 vssd1 vccd1 vccd1 _11129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11059_ _11359_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11060_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12469__S _12504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07152__A _07152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__A1 _07255_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07819__A1 _08633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__B2 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08270_ _08308_/A _08308_/B vssd1 vssd1 vccd1 vccd1 _08270_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _07221_/A _07221_/B vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__xnor2_4
X_07152_ _07152_/A _07153_/B vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09079__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07083_ _07428_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _07084_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout104 _07283_/X vssd1 vssd1 vccd1 vccd1 _10463_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11551__B2 _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__A1 _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _10468_/A vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__clkbuf_16
Xfanout126 _07163_/X vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07755__B1 fanout60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 _06942_/Y vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__clkbuf_8
Xfanout148 _07017_/X vssd1 vssd1 vccd1 vccd1 _08641_/A2 sky130_fd_sc_hd__clkbuf_8
X_07985_ _07985_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _07986_/C sky130_fd_sc_hd__xor2_1
X_06936_ _11975_/A _06936_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
X_09724_ _09400_/X _09402_/X _09724_/S vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__mux2_1
X_06867_ _12162_/A _06866_/X _06853_/X vssd1 vssd1 vccd1 vccd1 _06867_/X sky130_fd_sc_hd__a21o_1
X_09655_ _10234_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09542__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _08607_/B _08607_/C _08648_/A vssd1 vssd1 vccd1 vccd1 _08610_/A sky130_fd_sc_hd__o21ai_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__nand2_1
X_06798_ _12621_/A _07129_/A vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07062__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08546_/A _08546_/B _08530_/Y vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _08472_/A _08472_/B vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07419_ _07419_/A _07419_/B vssd1 vssd1 vccd1 vccd1 _07420_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10430_ _12349_/A _10429_/X hold283/A vssd1 vssd1 vccd1 vccd1 _10430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _08445_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _12202_/A _08274_/B fanout74/X _12059_/A vssd1 vssd1 vccd1 vccd1 _10362_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10593__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10292_ hold309/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10558_/C sky130_fd_sc_hd__or2_1
XANTENNA__11966__B _11966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ hold3/X fanout3/X hold273/X vssd1 vssd1 vccd1 vccd1 _13080_/X sky130_fd_sc_hd__a21o_1
X_12100_ _12339_/A1 _08792_/B _08792_/A vssd1 vssd1 vccd1 vccd1 _12100_/Y sky130_fd_sc_hd__a21oi_1
X_12031_ _11955_/B _11957_/B _11953_/X vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09735__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12143__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _13188_/A _13189_/A _13188_/B vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12797__B _12797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ hold295/X hold59/X vssd1 vssd1 vccd1 vccd1 _13170_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11058__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _12068_/A _11815_/B vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__xnor2_1
X_12795_ hold21/X _12797_/B vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__or2_1
XFILLER_0_126_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11760_/A sky130_fd_sc_hd__xor2_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11677_ _11677_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _11679_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10820__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10628_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06961__D _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08226__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__B2 _08551_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ _13372_/CLK _13347_/D vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__dfxtp_1
X_10559_ _12349_/A _10677_/B hold303/A vssd1 vssd1 vccd1 vccd1 _10559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ _13297_/CLK _13278_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _12280_/A _12229_/B _08798_/X vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__or3b_1
XANTENNA__11533__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A1 _09155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _10468_/A _07770_/B vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__xnor2_1
X_06721_ _06721_/A _11137_/S vssd1 vssd1 vccd1 vccd1 _06879_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09440_ _10310_/A _10310_/B _09440_/C vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__or3_2
X_06652_ _12179_/S vssd1 vssd1 vccd1 vccd1 _06652_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13038__A1 _10735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06583_ instruction[12] _06575_/X _06582_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ _09371_/A _09371_/B _09371_/C _09371_/D vssd1 vssd1 vccd1 vccd1 _09374_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08322_ _08648_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08312_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout132_A _07078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07204_ _09630_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07206_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _09403_/S _08184_/B vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07135_ _07135_/A _07135_/B _07135_/C vssd1 vssd1 vccd1 vccd1 _07138_/B sky130_fd_sc_hd__and3_1
XANTENNA__10575__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ reg1_val[9] _07066_/B vssd1 vssd1 vccd1 vccd1 _07066_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__A2 _07347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _08605_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _07970_/C sky130_fd_sc_hd__nand2_1
X_06919_ instruction[20] _06575_/X _06918_/X _06699_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09707_ _09369_/X _09541_/X _09542_/X vssd1 vssd1 vccd1 vccd1 _09707_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09272__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ _09671_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _07899_/Y sky130_fd_sc_hd__xnor2_1
X_09638_ _09493_/A _09493_/B _09490_/A vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _09431_/X _09568_/X _10286_/S vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__mux2_1
X_12580_ _12610_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _10772_/B _11219_/Y _11598_/Y _11599_/Y _11596_/Y vssd1 vssd1 vccd1 vccd1
+ _11601_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12252__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _09886_/B _12394_/A1 _11531_/S vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09211__S _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__A _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11462_ _12065_/A _11462_/B vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__xor2_1
X_11393_ _11291_/A _11291_/B _11299_/X vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__o21ba_1
X_13201_ _13226_/A hold270/X vssd1 vssd1 vccd1 vccd1 _13363_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _06816_/X _10412_/X _12025_/S vssd1 vssd1 vccd1 vccd1 _10414_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ hold308/A _13131_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_1
X_10344_ _10344_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10345_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07967__B1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07431__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13063_ hold123/A _13071_/A2 _13071_/B1 hold92/X _13016_/A vssd1 vssd1 vccd1 vccd1
+ hold93/A sky130_fd_sc_hd__o221a_1
X_10275_ _10315_/A _10276_/B _10276_/C vssd1 vssd1 vccd1 vccd1 _10275_/Y sky130_fd_sc_hd__o21ai_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _12014_/A _12085_/A vssd1 vssd1 vccd1 vccd1 _12016_/B sky130_fd_sc_hd__nor2_1
X_12916_ _13150_/A _13151_/A _13150_/B vssd1 vssd1 vccd1 vccd1 _13156_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07498__A2 _08400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ hold62/X _12847_/B vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12778_ hold1/X _12778_/B vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__nand2_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07430__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _12068_/A _11729_/B vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12951__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ _08940_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__nor2_2
X_08871_ _12310_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08874_/A sky130_fd_sc_hd__or2_2
X_07822_ _07821_/A _07821_/B _07821_/C vssd1 vssd1 vccd1 vccd1 _07825_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09092__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _09827_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07765_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06704_ _06704_/A _06704_/B vssd1 vssd1 vccd1 vccd1 _11428_/A sky130_fd_sc_hd__nand2_1
X_07684_ _08624_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__xnor2_2
X_06635_ _12115_/S _06635_/B vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__or2_2
XFILLER_0_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09423_ _09422_/X _09421_/Y _12396_/A _07129_/A vssd1 vssd1 vccd1 vccd1 _09423_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10966__A _10966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _08305_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08314_/B sky130_fd_sc_hd__xnor2_2
X_06566_ _12619_/A vssd1 vssd1 vccd1 vccd1 _06566_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08989__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09285_ _09285_/A _09285_/B vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ _08553_/A2 _10227_/B1 _10463_/A1 _08553_/B1 vssd1 vssd1 vccd1 vccd1 _08237_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08786_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09267__A _09766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _09928_/A _07814_/B _08553_/B1 fanout45/X vssd1 vssd1 vccd1 vccd1 _07119_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _10081_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _06949_/Y _06967_/A _06996_/A vssd1 vssd1 vccd1 vccd1 _07891_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ _10234_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07177__A1 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _11155_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10964_/B sky130_fd_sc_hd__xnor2_1
X_12701_ reg1_val[15] _12696_/B _12699_/A vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__a21o_2
X_10893_ _10812_/X _11041_/B _09148_/Y vssd1 vssd1 vccd1 vccd1 _10893_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07250__A _07251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ reg1_val[3] _12632_/B vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__nand2_1
X_12563_ _12568_/B _12563_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XFILLER_0_93_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _12495_/A _12495_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__a21o_1
X_11514_ _06704_/B _11426_/B _06704_/A vssd1 vssd1 vccd1 vccd1 _11515_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09929__A1 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _11422_/Y _11444_/X _06941_/X vssd1 vssd1 vccd1 vccd1 _11445_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11376_ _11376_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11379_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ _13115_/A _13115_/B vssd1 vssd1 vccd1 vccd1 _13116_/B sky130_fd_sc_hd__nand2_1
X_10327_ _10859_/A _07347_/B fanout14/X _10327_/B2 vssd1 vssd1 vccd1 vccd1 _10328_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06612__B1 _06767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10258_/A _10258_/B vssd1 vssd1 vccd1 vccd1 _10259_/B sky130_fd_sc_hd__xnor2_4
X_13046_ _11169_/A _13052_/A2 hold173/X vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__a21boi_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ _10189_/A _10189_/B vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09865__B1 _09148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10227__A1 _07593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09093__A1 _06875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11424__B1 _12029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ fanout62/X _10463_/B2 _10228_/A fanout60/X vssd1 vssd1 vccd1 vccd1 _09071_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__or2_1
XFILLER_0_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12506__A _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout6 fanout7/X vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09815__A _09815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _08910_/A _08910_/B _08911_/Y vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08356__B1 _08551_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08854_ _09297_/A1 fanout55/X _12257_/A _09297_/B2 vssd1 vssd1 vccd1 vccd1 _08855_/B
+ sky130_fd_sc_hd__o22a_1
X_08785_ _08060_/A _08060_/B _08784_/X vssd1 vssd1 vccd1 vccd1 _08789_/A sky130_fd_sc_hd__o21ai_1
X_07805_ _07858_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__nand2_1
X_07736_ _07736_/A _07736_/B vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ fanout71/X _10227_/B1 _10463_/A1 _08354_/A2 vssd1 vssd1 vccd1 vccd1 _07668_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__07331__B2 _07814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 _09928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06618_ reg2_val[30] _06767_/A _06707_/B1 _06617_/Y vssd1 vssd1 vccd1 vccd1 _08858_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_09406_ _09398_/X _09405_/X _10902_/A vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07882__A2 _08096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07598_/X sky130_fd_sc_hd__or2_1
XANTENNA__10218__B2 _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07070__A _09938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09337_ _07814_/B _10327_/B2 _10589_/A fanout45/X vssd1 vssd1 vccd1 vccd1 _09338_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09084__A1 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _09269_/B _09268_/B vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09084__B2 _11386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08219_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ _09191_/X _09198_/X _10284_/S vssd1 vssd1 vccd1 vccd1 _09199_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11230_ _11231_/A curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ fanout51/X _07347_/B fanout15/X _11456_/A vssd1 vssd1 vccd1 vccd1 _11162_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _09919_/A _09919_/B _09922_/A vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__a21o_2
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__or2_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ _07263_/Y _11645_/B _09950_/Y _09952_/Y vssd1 vssd1 vccd1 vccd1 _10044_/B
+ sky130_fd_sc_hd__a211o_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07245__A _09787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11990__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ _11995_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _12073_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09311__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ _10946_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07322__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _10876_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08076__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10209__A1 _07218_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10209__B2 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ reg1_val[27] curr_PC[27] _12615_/S vssd1 vssd1 vccd1 vccd1 _12616_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ reg1_val[16] curr_PC[16] _12615_/S vssd1 vssd1 vccd1 vccd1 _12547_/B sky130_fd_sc_hd__mux2_2
X_12477_ _12647_/B _12478_/B vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 instruction[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11230__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10932__A2 _07151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ hold176/X _13055_/A2 _13053_/B1 hold186/X _13057_/C1 vssd1 vssd1 vccd1 vccd1
+ hold187/A sky130_fd_sc_hd__o221a_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07155__A _07155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12996__A _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ _09301_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08571_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10448__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06994__A _06994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A _09370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _07518_/A _07518_/C _07518_/B vssd1 vssd1 vccd1 vccd1 _07522_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10448__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__B2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ _07451_/A _07451_/B _07480_/A vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07383_ _07419_/A _07419_/B vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _09123_/B _09123_/A vssd1 vssd1 vccd1 vccd1 _09122_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout212_A _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09053_ _10937_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09054_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08004_ _08533_/B _10067_/A1 _08926_/B1 _08507_/A2 vssd1 vssd1 vccd1 vccd1 _08005_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11176__A2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap240 _09669_/A vssd1 vssd1 vccd1 vccd1 _08648_/A sky130_fd_sc_hd__buf_6
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12125__A1 _06908_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _09955_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__xor2_1
X_09886_ _09886_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__nor2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08906_ _07651_/A _07651_/B _07649_/X vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__11884__B1 _09595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08837_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07001__B1 _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08768_ _08767_/B _08767_/C _08776_/B vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__a21o_1
X_08699_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__xor2_2
X_07719_ _07719_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10730_ _10587_/A _10587_/B _10589_/X vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__o21ai_1
X_10661_ _10660_/A _10660_/B _11612_/A vssd1 vssd1 vccd1 vccd1 _10661_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _12383_/Y _12384_/X _12399_/Y vssd1 vssd1 vccd1 vccd1 _12400_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ instruction[15] vssd1 vssd1 vccd1 vccd1 loadstore_dest[4] sky130_fd_sc_hd__buf_12
XFILLER_0_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ _11052_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08624__A _08624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12280_/A _12330_/Y _12374_/C vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12262_ _12262_/A _12315_/A vssd1 vssd1 vccd1 vccd1 _12263_/C sky130_fd_sc_hd__and2_1
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _11214_/A _11214_/B _11214_/C vssd1 vssd1 vccd1 vccd1 _11213_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06579__C1 _06699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12194_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10914__A2 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__A2 _08184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__B1 _07299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _09196_/S _11143_/Y _11142_/X _11138_/X vssd1 vssd1 vccd1 vccd1 _11144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _11191_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11077_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06798__B _07129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12824__C1 _13144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _11900_/A _07148_/C fanout6/X _12065_/A vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07703__A _08320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928_ _11149_/C _10927_/Y _12490_/S _10925_/X vssd1 vssd1 vccd1 vccd1 dest_val[12]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ _10859_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08534__A _08556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ _12530_/A _12530_/B _12530_/C vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12355__A1 _09237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A2 _09659_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__A1 _12171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A2 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06952_ _07202_/A _07264_/A _06952_/C _07097_/C vssd1 vssd1 vccd1 vccd1 _06954_/B
+ sky130_fd_sc_hd__or4_4
X_09740_ _09586_/A _09586_/B _06793_/A vssd1 vssd1 vccd1 vccd1 _09740_/X sky130_fd_sc_hd__a21bo_1
.ends

