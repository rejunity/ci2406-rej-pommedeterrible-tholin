// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    int_return,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_dest,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output int_return;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [4:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [4:0] loadstore_dest;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [4:0] reg1_idx;
 input [31:0] reg1_val;
 output [4:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(curr_PC[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(reg2_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(reg2_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(reg2_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(reg2_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(curr_PC[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(reg2_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(reg2_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg2_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg2_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg2_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg2_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg2_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(dest_pred_val));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg2_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg2_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(instruction[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(reg1_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(reg1_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg1_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg2_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg2_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg2_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg1_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(reg1_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(reg1_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06569__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A2 (.DIODE(_04670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__B (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__B (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__B (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__A2_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__B (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A_N (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__A (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06646__A (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06646__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__B (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06650__A2_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__A_N (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__B (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__B (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__A2_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A_N (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__B (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__A_N (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__B (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__B (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__A_N (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__B (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__B (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__B (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A_N (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A_N (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__B (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A2 (.DIODE(_04670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A3 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__B (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A2 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A3 (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__B (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__B (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__A3 (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__B (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__B (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__A3 (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__B (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__B (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A2 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A3 (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A3 (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__B (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__B (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A3 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__A2 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__A3 (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__B (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__B (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A3 (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__B (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A3 (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__C1 (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__C_N (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A3 (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A3 (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A3 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A3 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__B (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__B (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A3 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A3 (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__A3 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__A3 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__B (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__B (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__B (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A_N (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A_N (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__A_N (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__A_N (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__A_N (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A_N (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A_N (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__A_N (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__B (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__B (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__B (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__B (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__B (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__B (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__B (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A1 (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A (.DIODE(_04383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__B (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__B (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B (.DIODE(_06441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__C (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__C (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__B (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__C (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__D (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__D (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__B (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__B (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__C (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__D (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__B (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__C (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__D (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A1 (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__C1 (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A1 (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__S (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__A1 (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__B1 (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__B (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B1 (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__C_N (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__B1 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A (.DIODE(_00154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__B (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A (.DIODE(_00154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A1 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__S (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__C (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__C (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A3 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A4 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A3 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__A (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__A2 (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__C (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__D (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A3 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__B (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__A (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A3 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A4 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__C1 (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A3 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B1 (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__C1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A3 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A4 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A2 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__A (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A3 (.DIODE(_00183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A4 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__C (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A1 (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A1 (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__S (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A2 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A3 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__A (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A1 (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A1 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A1 (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__A (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B (.DIODE(_00343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B (.DIODE(_00343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A1 (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__B2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A1 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A1 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__C (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A2 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A1 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B2 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B2 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A2 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__B2 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B2 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__B2 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A2 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A1 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A1 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__B1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A3 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__B (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__B1 (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B1 (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__B (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__B (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__B1 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A2 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__B1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B2 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B2 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__B2 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__B2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A1 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__B2 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A1 (.DIODE(_00154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A2 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A1 (.DIODE(_00154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A2 (.DIODE(_00155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__B1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A (.DIODE(_01419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A (.DIODE(_01419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__A (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A (.DIODE(_01573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A2 (.DIODE(_01573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08500__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08500__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A (.DIODE(_01573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A2 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A2 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__B1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__B1 (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__A2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A2 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__B1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A0 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A2 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__B1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A2 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__B1 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A1 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__B2 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__B (.DIODE(_01926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__B (.DIODE(_01926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A2 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08836__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A2 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__B1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B (.DIODE(_01962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__D (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A4 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__A1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A3 (.DIODE(_01962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A2 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__B2 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__B1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__B1 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__B1 (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__D1 (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A1 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__B2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__B2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__B2 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09069__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A2 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A3 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A1 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__B (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__S (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__S (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09165__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__S (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A2 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A2 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__B1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A1 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A1 (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A2 (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__B (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__C (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__B1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A1 (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__B (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A1_N (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__S (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__S (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A2 (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A3 (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A3 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A3 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A2 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A2 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__A1_N (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__B1 (.DIODE(_02532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A2 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__A2 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__B1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__B2 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A2 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__B (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A1 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__B2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__B1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A2 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B1 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__A (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A1 (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A2 (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__B (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__C (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__A (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__S (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A2 (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__C1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A1 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A2 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B1 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__B1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A2 (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A2 (.DIODE(_02847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A1 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__B2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A2 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A3 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__B1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__B1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__B1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__A3 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B1 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__B1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__B1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A1 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__B2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__B2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__B2 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A2 (.DIODE(_03125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10041__A1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__C1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A2 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__A3 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__B2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__B2 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A2 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B2 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A1 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__B1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__B1 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__A1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__B2 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A1 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A2 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B1 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A1 (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A2 (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__C (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A2 (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A2 (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__S (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__S (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A1_N (.DIODE(_06285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A2_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B1_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A2 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__B1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A2 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A3 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A1 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B2 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__B (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__B (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A (.DIODE(_03410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__C1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A1_N (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A2_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__A (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A1 (.DIODE(_00687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A2 (.DIODE(_00688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__B (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__C (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__B1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A2 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__B1 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__A1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B2 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__S (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__C1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B2 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__B2 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A1 (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__B (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__B (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A2 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B1 (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A2 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A3 (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__S (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A1_N (.DIODE(_06148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A2_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__B2 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A2 (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B2 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__A1 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__B2 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A1 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__B2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__A (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__A (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A2 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__B1 (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__B (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__B (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__C1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__S (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A1_N (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A2_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__A (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__B (.DIODE(_03858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A_N (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__B1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__A1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B2 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A1 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__B2 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A2 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A3 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10838__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10840__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A1 (.DIODE(_03410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__A2 (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A2 (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__C1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A1 (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__A2 (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B2 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__A1 (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A2 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__C1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__S (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__C (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__B (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A1 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__B2 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B2 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A1 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B2 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11083__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11083__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A1 (.DIODE(_03739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__C (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__B1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A1_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A2_N (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A1_N (.DIODE(_05965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A2_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B2 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A1 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A2 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A2 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__C1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__S (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A1 (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A1_N (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__B (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__B (.DIODE(_04355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__B (.DIODE(_04355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A1 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__B2 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A1 (.DIODE(_03410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__B1 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__A3 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A2_N (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B2 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A1_N (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__A1_N (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__A3 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__B1 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__B2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__A1 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__B2 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A2 (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A2 (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__A (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__B (.DIODE(_04516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__B1 (.DIODE(_04550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__C (.DIODE(_04550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A1 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__B2 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A2 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__B1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A1 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B2 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__B1 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__A3 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11532__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__B2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B1 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B2 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B1 (.DIODE(_05766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A2 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A (.DIODE(_04550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A (.DIODE(_04550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A (.DIODE(_04694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__A (.DIODE(_04694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__B1 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A3 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11618__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__C1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__B1 (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__B2 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A1 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A3 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__B1 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A1 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A2 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__B2 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__C1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__B1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__B2 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A1 (.DIODE(_05550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A3 (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__B1 (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__B (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A1 (.DIODE(_04694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B1 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A0 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__B2 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A1 (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__B (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__D (.DIODE(_04706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A2 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__B1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B1 (.DIODE(_04980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A1 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A2 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__B2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A2 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A1 (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__B1 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__B (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__C (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__A1 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11948__A2 (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11948__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__C1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__C1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__11966__B (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__A1 (.DIODE(_05410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__B (.DIODE(_05081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A2 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A1 (.DIODE(_04980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__C1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A0 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__A1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__B1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__C1 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B1 (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A2 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__C1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__A2 (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B2 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__C1 (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__C1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(_05312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A1 (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__C (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__A1 (.DIODE(_05040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__C1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__B2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B2 (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__B1 (.DIODE(_00668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__C1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A2 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__C1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A2 (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__C1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A2 (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12350__B1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A2 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12354__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__C1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A2 (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__B1 (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__C1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12415__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A2 (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__B1 (.DIODE(_02321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A1 (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A2 (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__B2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__B1 (.DIODE(_05603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A1 (.DIODE(_05258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__A (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__A (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__A (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__A (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__B (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__B (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__A (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__B (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__B (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__B (.DIODE(_05676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B (.DIODE(_05676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__A (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__B (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__B (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__B (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__B (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__B (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__B (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__B (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__B (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__B (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__B (.DIODE(_05528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__B (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__B (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__B (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__B (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__B (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__B (.DIODE(_05388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__B (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__B (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__B (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__B (.DIODE(_05019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__B (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__B (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__B (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__B (.DIODE(_04779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__B (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A2 (.DIODE(_04942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A2_N (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__B (.DIODE(_00186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__B (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A (.DIODE(_04383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(_04383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A1 (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A1 (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A1 (.DIODE(_00243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A1 (.DIODE(_00211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A1 (.DIODE(_00198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A1 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A1 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A1 (.DIODE(_00315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A2 (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__C1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__B (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A1 (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__C1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A1 (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__C1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__C1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__A1 (.DIODE(_00347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A1 (.DIODE(_00334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A2 (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A1 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A2 (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__C1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A1 (.DIODE(_00148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A1 (.DIODE(_06522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A1 (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A2 (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A1 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__C1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__B (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__B (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A1 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__B (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A1 (.DIODE(_00690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A1 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__B (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A1 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A1 (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A1 (.DIODE(_00328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__A1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A1 (.DIODE(_00343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A1 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__A2 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__C (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__A2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__B (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13228__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__13274__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13297__CLK (.DIODE(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(_00165_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_00165_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(_00242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(_06464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(_05931_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(_02082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(_05930_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(_02082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(_00140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(_06449_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(_02082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_02081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(_00312_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(_04383_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(_00312_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_04670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(_04670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(_00269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(_00156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(_00156_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(_00149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(_00149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(_06535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_06535_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap102_A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap109_A (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap112_A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap115_A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap118_A (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(_02069_));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06561_ (.A(net300),
    .Y(_04350_));
 sky130_fd_sc_hd__inv_2 _06562_ (.A(net318),
    .Y(_04361_));
 sky130_fd_sc_hd__inv_2 _06563_ (.A(net338),
    .Y(_04372_));
 sky130_fd_sc_hd__inv_2 _06564_ (.A(net261),
    .Y(_04383_));
 sky130_fd_sc_hd__inv_2 _06565_ (.A(instruction[3]),
    .Y(_04394_));
 sky130_fd_sc_hd__inv_2 _06566_ (.A(net292),
    .Y(_04405_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(instruction[41]),
    .Y(_04416_));
 sky130_fd_sc_hd__inv_6 _06568_ (.A(reg1_val[31]),
    .Y(_04427_));
 sky130_fd_sc_hd__inv_2 _06569_ (.A(net294),
    .Y(_04438_));
 sky130_fd_sc_hd__inv_2 _06570_ (.A(rst),
    .Y(_04448_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(instruction[0]),
    .B(pred_val),
    .Y(_04459_));
 sky130_fd_sc_hd__and2_1 _06572_ (.A(pred_val),
    .B(instruction[1]),
    .X(_04470_));
 sky130_fd_sc_hd__o31a_1 _06573_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(pred_val),
    .X(_04481_));
 sky130_fd_sc_hd__and4b_4 _06574_ (.A_N(instruction[1]),
    .B(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04492_));
 sky130_fd_sc_hd__or3b_4 _06575_ (.A(_04470_),
    .B(_04459_),
    .C_N(instruction[2]),
    .X(_04503_));
 sky130_fd_sc_hd__or2_1 _06576_ (.A(instruction[20]),
    .B(_04492_),
    .X(_04514_));
 sky130_fd_sc_hd__o211a_4 _06577_ (.A1(instruction[13]),
    .A2(_04503_),
    .B1(_04514_),
    .C1(net273),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__or2_1 _06578_ (.A(instruction[21]),
    .B(_04492_),
    .X(_04535_));
 sky130_fd_sc_hd__o211a_4 _06579_ (.A1(instruction[14]),
    .A2(_04503_),
    .B1(_04535_),
    .C1(net273),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__or2_1 _06580_ (.A(instruction[18]),
    .B(_04492_),
    .X(_04555_));
 sky130_fd_sc_hd__o211a_4 _06581_ (.A1(instruction[11]),
    .A2(_04503_),
    .B1(_04555_),
    .C1(net273),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__or2_1 _06582_ (.A(instruction[19]),
    .B(_04492_),
    .X(_04576_));
 sky130_fd_sc_hd__o211a_4 _06583_ (.A1(instruction[12]),
    .A2(_04503_),
    .B1(_04576_),
    .C1(net273),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__or2_1 _06584_ (.A(instruction[22]),
    .B(_04492_),
    .X(_04597_));
 sky130_fd_sc_hd__o211a_4 _06585_ (.A1(instruction[15]),
    .A2(_04503_),
    .B1(_04597_),
    .C1(net273),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__or4bb_4 _06586_ (.A(instruction[0]),
    .B(instruction[1]),
    .C_N(instruction[2]),
    .D_N(pred_val),
    .X(_04618_));
 sky130_fd_sc_hd__nor2_8 _06587_ (.A(instruction[3]),
    .B(_04618_),
    .Y(is_load));
 sky130_fd_sc_hd__nor2_8 _06588_ (.A(_04394_),
    .B(_04618_),
    .Y(is_store));
 sky130_fd_sc_hd__and4bb_1 _06589_ (.A_N(instruction[0]),
    .B_N(instruction[2]),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04648_));
 sky130_fd_sc_hd__or4bb_1 _06590_ (.A(instruction[0]),
    .B(instruction[2]),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04659_));
 sky130_fd_sc_hd__o311a_4 _06591_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04670_));
 sky130_fd_sc_hd__and4bb_2 _06592_ (.A_N(instruction[1]),
    .B_N(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04681_));
 sky130_fd_sc_hd__or4bb_4 _06593_ (.A(instruction[1]),
    .B(instruction[2]),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04692_));
 sky130_fd_sc_hd__and2_4 _06594_ (.A(instruction[25]),
    .B(net273),
    .X(_04703_));
 sky130_fd_sc_hd__o211a_1 _06595_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04714_));
 sky130_fd_sc_hd__o211ai_1 _06596_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04725_));
 sky130_fd_sc_hd__a21o_1 _06597_ (.A1(instruction[41]),
    .A2(_04681_),
    .B1(_04714_),
    .X(_04736_));
 sky130_fd_sc_hd__a21oi_4 _06598_ (.A1(instruction[41]),
    .A2(_04681_),
    .B1(_04714_),
    .Y(_04746_));
 sky130_fd_sc_hd__a221o_2 _06599_ (.A1(instruction[24]),
    .A2(_04670_),
    .B1(_04681_),
    .B2(instruction[41]),
    .C1(_04714_),
    .X(_04757_));
 sky130_fd_sc_hd__nand2_4 _06600_ (.A(net272),
    .B(_04757_),
    .Y(_04768_));
 sky130_fd_sc_hd__and2_4 _06601_ (.A(instruction[39]),
    .B(net274),
    .X(_04779_));
 sky130_fd_sc_hd__nor2_1 _06602_ (.A(net253),
    .B(_04779_),
    .Y(_04790_));
 sky130_fd_sc_hd__o2bb2a_1 _06603_ (.A1_N(reg2_val[29]),
    .A2_N(net268),
    .B1(net225),
    .B2(_04790_),
    .X(_04801_));
 sky130_fd_sc_hd__a2bb2o_2 _06604_ (.A1_N(_04790_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[29]),
    .X(_04812_));
 sky130_fd_sc_hd__and2_1 _06605_ (.A(reg1_val[29]),
    .B(_04812_),
    .X(_04823_));
 sky130_fd_sc_hd__or2_1 _06606_ (.A(reg1_val[29]),
    .B(_04812_),
    .X(_04834_));
 sky130_fd_sc_hd__and2b_1 _06607_ (.A_N(_04823_),
    .B(_04834_),
    .X(_04844_));
 sky130_fd_sc_hd__inv_2 _06608_ (.A(_04844_),
    .Y(_04855_));
 sky130_fd_sc_hd__and2_4 _06609_ (.A(instruction[38]),
    .B(net274),
    .X(_04866_));
 sky130_fd_sc_hd__nor2_1 _06610_ (.A(net253),
    .B(_04866_),
    .Y(_04877_));
 sky130_fd_sc_hd__o2bb2a_1 _06611_ (.A1_N(reg2_val[28]),
    .A2_N(net268),
    .B1(net225),
    .B2(_04877_),
    .X(_04888_));
 sky130_fd_sc_hd__a2bb2o_4 _06612_ (.A1_N(_04877_),
    .A2_N(net225),
    .B1(net270),
    .B2(reg2_val[28]),
    .X(_04899_));
 sky130_fd_sc_hd__and2_1 _06613_ (.A(reg1_val[28]),
    .B(_04899_),
    .X(_04910_));
 sky130_fd_sc_hd__or2_1 _06614_ (.A(reg1_val[28]),
    .B(_04899_),
    .X(_04921_));
 sky130_fd_sc_hd__and2b_1 _06615_ (.A_N(_04910_),
    .B(_04921_),
    .X(_04931_));
 sky130_fd_sc_hd__and2_4 _06616_ (.A(instruction[40]),
    .B(net274),
    .X(_04942_));
 sky130_fd_sc_hd__nor2_1 _06617_ (.A(net253),
    .B(_04942_),
    .Y(_04953_));
 sky130_fd_sc_hd__o2bb2a_1 _06618_ (.A1_N(reg2_val[30]),
    .A2_N(net270),
    .B1(net225),
    .B2(_04953_),
    .X(_04964_));
 sky130_fd_sc_hd__a2bb2o_4 _06619_ (.A1_N(_04953_),
    .A2_N(net225),
    .B1(net269),
    .B2(reg2_val[30]),
    .X(_04975_));
 sky130_fd_sc_hd__and2_1 _06620_ (.A(reg1_val[30]),
    .B(_04975_),
    .X(_04986_));
 sky130_fd_sc_hd__nor2_1 _06621_ (.A(reg1_val[30]),
    .B(_04975_),
    .Y(_04997_));
 sky130_fd_sc_hd__or2_2 _06622_ (.A(_04986_),
    .B(_04997_),
    .X(_05008_));
 sky130_fd_sc_hd__and2_4 _06623_ (.A(instruction[37]),
    .B(net274),
    .X(_05019_));
 sky130_fd_sc_hd__nor2_1 _06624_ (.A(net253),
    .B(_05019_),
    .Y(_05029_));
 sky130_fd_sc_hd__o2bb2a_2 _06625_ (.A1_N(reg2_val[27]),
    .A2_N(net269),
    .B1(_04768_),
    .B2(_05029_),
    .X(_05040_));
 sky130_fd_sc_hd__and2b_1 _06626_ (.A_N(reg1_val[27]),
    .B(_05040_),
    .X(_05051_));
 sky130_fd_sc_hd__nand2b_1 _06627_ (.A_N(_05040_),
    .B(reg1_val[27]),
    .Y(_05062_));
 sky130_fd_sc_hd__nand2b_2 _06628_ (.A_N(_05051_),
    .B(_05062_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _06629_ (.A(_05008_),
    .B(_05073_),
    .Y(_05084_));
 sky130_fd_sc_hd__and2_4 _06630_ (.A(instruction[35]),
    .B(net274),
    .X(_05095_));
 sky130_fd_sc_hd__nor2_1 _06631_ (.A(_04746_),
    .B(_05095_),
    .Y(_05106_));
 sky130_fd_sc_hd__o2bb2a_4 _06632_ (.A1_N(reg2_val[25]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05106_),
    .X(_05116_));
 sky130_fd_sc_hd__and2b_1 _06633_ (.A_N(_05116_),
    .B(reg1_val[25]),
    .X(_05127_));
 sky130_fd_sc_hd__and2b_1 _06634_ (.A_N(reg1_val[25]),
    .B(_05116_),
    .X(_05138_));
 sky130_fd_sc_hd__or2_2 _06635_ (.A(_05127_),
    .B(_05138_),
    .X(_05149_));
 sky130_fd_sc_hd__and2_4 _06636_ (.A(instruction[34]),
    .B(net274),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_1 _06637_ (.A(net253),
    .B(_05160_),
    .Y(_05171_));
 sky130_fd_sc_hd__o2bb2a_2 _06638_ (.A1_N(reg2_val[24]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05171_),
    .X(_05182_));
 sky130_fd_sc_hd__a2bb2o_1 _06639_ (.A1_N(_05171_),
    .A2_N(net225),
    .B1(net269),
    .B2(reg2_val[24]),
    .X(_05193_));
 sky130_fd_sc_hd__nand2_1 _06640_ (.A(reg1_val[24]),
    .B(_05193_),
    .Y(_05203_));
 sky130_fd_sc_hd__or2_1 _06641_ (.A(reg1_val[24]),
    .B(_05193_),
    .X(_05214_));
 sky130_fd_sc_hd__nand2_2 _06642_ (.A(_05203_),
    .B(_05214_),
    .Y(_05225_));
 sky130_fd_sc_hd__and2_1 _06643_ (.A(reg2_val[31]),
    .B(net269),
    .X(_05236_));
 sky130_fd_sc_hd__o21ba_2 _06644_ (.A1(_04416_),
    .A2(_04768_),
    .B1_N(_05236_),
    .X(_05247_));
 sky130_fd_sc_hd__a31o_4 _06645_ (.A1(instruction[41]),
    .A2(net272),
    .A3(_04757_),
    .B1(_05236_),
    .X(_05258_));
 sky130_fd_sc_hd__xnor2_2 _06646_ (.A(_04427_),
    .B(_05258_),
    .Y(_05269_));
 sky130_fd_sc_hd__xnor2_4 _06647_ (.A(reg1_val[31]),
    .B(_05258_),
    .Y(_05279_));
 sky130_fd_sc_hd__and2_4 _06648_ (.A(instruction[36]),
    .B(net274),
    .X(_05290_));
 sky130_fd_sc_hd__nor2_1 _06649_ (.A(net253),
    .B(_05290_),
    .Y(_05301_));
 sky130_fd_sc_hd__o2bb2a_4 _06650_ (.A1_N(reg2_val[26]),
    .A2_N(net270),
    .B1(_04768_),
    .B2(_05301_),
    .X(_05312_));
 sky130_fd_sc_hd__and2b_1 _06651_ (.A_N(_05312_),
    .B(reg1_val[26]),
    .X(_05323_));
 sky130_fd_sc_hd__inv_2 _06652_ (.A(_05323_),
    .Y(_05334_));
 sky130_fd_sc_hd__and2b_1 _06653_ (.A_N(reg1_val[26]),
    .B(_05312_),
    .X(_05344_));
 sky130_fd_sc_hd__or2_2 _06654_ (.A(_05323_),
    .B(_05344_),
    .X(_05355_));
 sky130_fd_sc_hd__and4_1 _06655_ (.A(_05149_),
    .B(_05225_),
    .C(_05279_),
    .D(_05355_),
    .X(_05366_));
 sky130_fd_sc_hd__or4b_1 _06656_ (.A(_04844_),
    .B(_04931_),
    .C(_05084_),
    .D_N(_05366_),
    .X(_05377_));
 sky130_fd_sc_hd__and2_4 _06657_ (.A(instruction[33]),
    .B(net274),
    .X(_05388_));
 sky130_fd_sc_hd__nor2_1 _06658_ (.A(net253),
    .B(_05388_),
    .Y(_05399_));
 sky130_fd_sc_hd__o2bb2a_4 _06659_ (.A1_N(reg2_val[23]),
    .A2_N(net270),
    .B1(_04768_),
    .B2(_05399_),
    .X(_05410_));
 sky130_fd_sc_hd__and2b_1 _06660_ (.A_N(_05410_),
    .B(reg1_val[23]),
    .X(_05420_));
 sky130_fd_sc_hd__and2b_1 _06661_ (.A_N(reg1_val[23]),
    .B(_05410_),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_2 _06662_ (.A(_05420_),
    .B(_05431_),
    .Y(_05442_));
 sky130_fd_sc_hd__and2_4 _06663_ (.A(instruction[32]),
    .B(net273),
    .X(_05453_));
 sky130_fd_sc_hd__nor2_1 _06664_ (.A(net253),
    .B(_05453_),
    .Y(_05464_));
 sky130_fd_sc_hd__o2bb2a_4 _06665_ (.A1_N(reg2_val[22]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05464_),
    .X(_05474_));
 sky130_fd_sc_hd__a2bb2o_4 _06666_ (.A1_N(_05464_),
    .A2_N(_04768_),
    .B1(net269),
    .B2(reg2_val[22]),
    .X(_05485_));
 sky130_fd_sc_hd__and2_1 _06667_ (.A(reg1_val[22]),
    .B(_05485_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _06668_ (.A(reg1_val[22]),
    .B(_05485_),
    .Y(_05507_));
 sky130_fd_sc_hd__nor2_2 _06669_ (.A(_05496_),
    .B(_05507_),
    .Y(_05518_));
 sky130_fd_sc_hd__and2_4 _06670_ (.A(instruction[30]),
    .B(net273),
    .X(_05528_));
 sky130_fd_sc_hd__nor2_1 _06671_ (.A(net253),
    .B(_05528_),
    .Y(_05539_));
 sky130_fd_sc_hd__o2bb2a_4 _06672_ (.A1_N(reg2_val[20]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05539_),
    .X(_05550_));
 sky130_fd_sc_hd__and2b_1 _06673_ (.A_N(_05550_),
    .B(reg1_val[20]),
    .X(_05561_));
 sky130_fd_sc_hd__and2b_1 _06674_ (.A_N(reg1_val[20]),
    .B(_05550_),
    .X(_05572_));
 sky130_fd_sc_hd__nor2_2 _06675_ (.A(_05561_),
    .B(_05572_),
    .Y(_05582_));
 sky130_fd_sc_hd__o311a_4 _06676_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05593_));
 sky130_fd_sc_hd__nor2_1 _06677_ (.A(net253),
    .B(_05593_),
    .Y(_05604_));
 sky130_fd_sc_hd__o2bb2a_2 _06678_ (.A1_N(reg2_val[21]),
    .A2_N(net269),
    .B1(_04768_),
    .B2(_05604_),
    .X(_05614_));
 sky130_fd_sc_hd__inv_2 _06679_ (.A(_05614_),
    .Y(_05623_));
 sky130_fd_sc_hd__and2_1 _06680_ (.A(reg1_val[21]),
    .B(_05623_),
    .X(_05633_));
 sky130_fd_sc_hd__nor2_1 _06681_ (.A(reg1_val[21]),
    .B(_05623_),
    .Y(_05642_));
 sky130_fd_sc_hd__nor2_2 _06682_ (.A(_05633_),
    .B(_05642_),
    .Y(_05652_));
 sky130_fd_sc_hd__nor4_1 _06683_ (.A(_05442_),
    .B(_05518_),
    .C(_05582_),
    .D(_05652_),
    .Y(_05662_));
 sky130_fd_sc_hd__inv_2 _06684_ (.A(_05662_),
    .Y(_05671_));
 sky130_fd_sc_hd__and2_4 _06685_ (.A(instruction[29]),
    .B(net273),
    .X(_05681_));
 sky130_fd_sc_hd__nor2_1 _06686_ (.A(net253),
    .B(_05681_),
    .Y(_05690_));
 sky130_fd_sc_hd__o2bb2a_4 _06687_ (.A1_N(reg2_val[19]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05690_),
    .X(_05700_));
 sky130_fd_sc_hd__and2b_1 _06688_ (.A_N(_05700_),
    .B(reg1_val[19]),
    .X(_05709_));
 sky130_fd_sc_hd__and2b_1 _06689_ (.A_N(reg1_val[19]),
    .B(_05700_),
    .X(_05719_));
 sky130_fd_sc_hd__or2_2 _06690_ (.A(_05709_),
    .B(_05719_),
    .X(_05728_));
 sky130_fd_sc_hd__and2_4 _06691_ (.A(instruction[28]),
    .B(net273),
    .X(_05738_));
 sky130_fd_sc_hd__nor2_1 _06692_ (.A(net253),
    .B(_05738_),
    .Y(_05747_));
 sky130_fd_sc_hd__o2bb2a_2 _06693_ (.A1_N(reg2_val[18]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05747_),
    .X(_05757_));
 sky130_fd_sc_hd__a2bb2o_4 _06694_ (.A1_N(_05747_),
    .A2_N(net225),
    .B1(net269),
    .B2(reg2_val[18]),
    .X(_05766_));
 sky130_fd_sc_hd__and2_1 _06695_ (.A(reg1_val[18]),
    .B(_05766_),
    .X(_05775_));
 sky130_fd_sc_hd__nor2_1 _06696_ (.A(reg1_val[18]),
    .B(_05766_),
    .Y(_05784_));
 sky130_fd_sc_hd__nor2_1 _06697_ (.A(_05775_),
    .B(_05784_),
    .Y(_05793_));
 sky130_fd_sc_hd__or2_1 _06698_ (.A(_05775_),
    .B(_05784_),
    .X(_05802_));
 sky130_fd_sc_hd__and2_4 _06699_ (.A(instruction[27]),
    .B(net273),
    .X(_05811_));
 sky130_fd_sc_hd__nor2_1 _06700_ (.A(net253),
    .B(_05811_),
    .Y(_05820_));
 sky130_fd_sc_hd__o2bb2a_4 _06701_ (.A1_N(reg2_val[17]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05820_),
    .X(_05829_));
 sky130_fd_sc_hd__nand2b_1 _06702_ (.A_N(_05829_),
    .B(reg1_val[17]),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2b_1 _06703_ (.A_N(reg1_val[17]),
    .B(_05829_),
    .Y(_05848_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(_05838_),
    .B(_05848_),
    .Y(_05857_));
 sky130_fd_sc_hd__o311a_4 _06705_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[26]),
    .C1(pred_val),
    .X(_05865_));
 sky130_fd_sc_hd__nor2_1 _06706_ (.A(net253),
    .B(_05865_),
    .Y(_05874_));
 sky130_fd_sc_hd__o2bb2a_4 _06707_ (.A1_N(reg2_val[16]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05874_),
    .X(_05883_));
 sky130_fd_sc_hd__and2b_1 _06708_ (.A_N(_05883_),
    .B(reg1_val[16]),
    .X(_05892_));
 sky130_fd_sc_hd__and2b_1 _06709_ (.A_N(reg1_val[16]),
    .B(_05883_),
    .X(_05901_));
 sky130_fd_sc_hd__inv_2 _06710_ (.A(_05901_),
    .Y(_05910_));
 sky130_fd_sc_hd__or2_1 _06711_ (.A(_05892_),
    .B(_05901_),
    .X(_05919_));
 sky130_fd_sc_hd__and2_1 _06712_ (.A(reg2_val[15]),
    .B(net269),
    .X(_05928_));
 sky130_fd_sc_hd__a31o_4 _06713_ (.A1(net272),
    .A2(_04670_),
    .A3(net253),
    .B1(_05928_),
    .X(_05935_));
 sky130_fd_sc_hd__and2_1 _06714_ (.A(net290),
    .B(_05935_),
    .X(_05941_));
 sky130_fd_sc_hd__nor2_1 _06715_ (.A(net290),
    .B(_05935_),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _06716_ (.A(_05941_),
    .B(_05947_),
    .Y(_05953_));
 sky130_fd_sc_hd__and2_1 _06717_ (.A(reg2_val[14]),
    .B(net270),
    .X(_05959_));
 sky130_fd_sc_hd__a31o_4 _06718_ (.A1(net271),
    .A2(_04746_),
    .A3(_04942_),
    .B1(_05959_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_1 _06719_ (.A(net291),
    .B(_05965_),
    .Y(_05971_));
 sky130_fd_sc_hd__and2_1 _06720_ (.A(net291),
    .B(_05965_),
    .X(_05982_));
 sky130_fd_sc_hd__nor2_2 _06721_ (.A(_05971_),
    .B(_05982_),
    .Y(_05993_));
 sky130_fd_sc_hd__inv_2 _06722_ (.A(_05993_),
    .Y(_06004_));
 sky130_fd_sc_hd__and2_1 _06723_ (.A(reg2_val[13]),
    .B(net268),
    .X(_06015_));
 sky130_fd_sc_hd__a31o_4 _06724_ (.A1(net271),
    .A2(net252),
    .A3(_04779_),
    .B1(_06015_),
    .X(_06026_));
 sky130_fd_sc_hd__and2_1 _06725_ (.A(reg1_val[13]),
    .B(_06026_),
    .X(_06037_));
 sky130_fd_sc_hd__nor2_1 _06726_ (.A(reg1_val[13]),
    .B(_06026_),
    .Y(_06048_));
 sky130_fd_sc_hd__nor2_1 _06727_ (.A(_06037_),
    .B(_06048_),
    .Y(_06059_));
 sky130_fd_sc_hd__and2_1 _06728_ (.A(reg2_val[12]),
    .B(net270),
    .X(_06070_));
 sky130_fd_sc_hd__a31o_4 _06729_ (.A1(net272),
    .A2(net252),
    .A3(_04866_),
    .B1(_06070_),
    .X(_06081_));
 sky130_fd_sc_hd__and2_1 _06730_ (.A(reg1_val[12]),
    .B(_06081_),
    .X(_06088_));
 sky130_fd_sc_hd__nor2_1 _06731_ (.A(reg1_val[12]),
    .B(_06081_),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_2 _06732_ (.A(_06088_),
    .B(_06094_),
    .Y(_06100_));
 sky130_fd_sc_hd__inv_2 _06733_ (.A(_06100_),
    .Y(_06106_));
 sky130_fd_sc_hd__and2_1 _06734_ (.A(reg2_val[11]),
    .B(net268),
    .X(_06112_));
 sky130_fd_sc_hd__a31o_4 _06735_ (.A1(net272),
    .A2(_04746_),
    .A3(_05019_),
    .B1(_06112_),
    .X(_06118_));
 sky130_fd_sc_hd__and2_1 _06736_ (.A(reg1_val[11]),
    .B(_06118_),
    .X(_06124_));
 sky130_fd_sc_hd__nor2_1 _06737_ (.A(reg1_val[11]),
    .B(_06118_),
    .Y(_06130_));
 sky130_fd_sc_hd__nor2_1 _06738_ (.A(_06124_),
    .B(_06130_),
    .Y(_06136_));
 sky130_fd_sc_hd__and2_1 _06739_ (.A(reg2_val[10]),
    .B(net270),
    .X(_06142_));
 sky130_fd_sc_hd__a31o_4 _06740_ (.A1(net271),
    .A2(net252),
    .A3(_05290_),
    .B1(_06142_),
    .X(_06148_));
 sky130_fd_sc_hd__nor2_1 _06741_ (.A(reg1_val[10]),
    .B(_06148_),
    .Y(_06154_));
 sky130_fd_sc_hd__and2_1 _06742_ (.A(reg1_val[10]),
    .B(_06148_),
    .X(_06160_));
 sky130_fd_sc_hd__nor2_1 _06743_ (.A(_06154_),
    .B(_06160_),
    .Y(_06169_));
 sky130_fd_sc_hd__and2_1 _06744_ (.A(reg2_val[9]),
    .B(net270),
    .X(_06178_));
 sky130_fd_sc_hd__a31o_4 _06745_ (.A1(net271),
    .A2(net252),
    .A3(_05095_),
    .B1(_06178_),
    .X(_06187_));
 sky130_fd_sc_hd__inv_2 _06746_ (.A(_06187_),
    .Y(_06196_));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(reg1_val[9]),
    .B(_06187_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand2_1 _06748_ (.A(reg1_val[9]),
    .B(_06187_),
    .Y(_06214_));
 sky130_fd_sc_hd__nand2b_1 _06749_ (.A_N(_06205_),
    .B(_06214_),
    .Y(_06223_));
 sky130_fd_sc_hd__and2_1 _06750_ (.A(reg2_val[8]),
    .B(net268),
    .X(_06232_));
 sky130_fd_sc_hd__a31o_4 _06751_ (.A1(net271),
    .A2(_04746_),
    .A3(_05160_),
    .B1(_06232_),
    .X(_06241_));
 sky130_fd_sc_hd__nor2_1 _06752_ (.A(reg1_val[8]),
    .B(_06241_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand2_1 _06753_ (.A(reg1_val[8]),
    .B(_06241_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand2b_1 _06754_ (.A_N(_06249_),
    .B(_06258_),
    .Y(_06267_));
 sky130_fd_sc_hd__and2_1 _06755_ (.A(reg2_val[7]),
    .B(net268),
    .X(_06276_));
 sky130_fd_sc_hd__a31o_4 _06756_ (.A1(net271),
    .A2(net252),
    .A3(_05388_),
    .B1(_06276_),
    .X(_06285_));
 sky130_fd_sc_hd__nor2_1 _06757_ (.A(reg1_val[7]),
    .B(_06285_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _06758_ (.A(reg1_val[7]),
    .B(_06285_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2b_2 _06759_ (.A_N(_06292_),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__and2_1 _06760_ (.A(reg2_val[6]),
    .B(net268),
    .X(_06301_));
 sky130_fd_sc_hd__a31o_4 _06761_ (.A1(net271),
    .A2(net252),
    .A3(_05453_),
    .B1(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__or2_1 _06762_ (.A(reg1_val[6]),
    .B(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__inv_2 _06763_ (.A(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__and2_1 _06764_ (.A(reg1_val[6]),
    .B(_06302_),
    .X(_06305_));
 sky130_fd_sc_hd__nor2_1 _06765_ (.A(_06304_),
    .B(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__o2111a_1 _06766_ (.A1(_04416_),
    .A2(_04692_),
    .B1(_04725_),
    .C1(_05593_),
    .D1(net272),
    .X(_06307_));
 sky130_fd_sc_hd__or3b_2 _06767_ (.A(net270),
    .B(_04736_),
    .C_N(_05593_),
    .X(_06308_));
 sky130_fd_sc_hd__a21oi_4 _06768_ (.A1(reg2_val[5]),
    .A2(net268),
    .B1(net251),
    .Y(_06309_));
 sky130_fd_sc_hd__a21o_2 _06769_ (.A1(reg2_val[5]),
    .A2(net268),
    .B1(net251),
    .X(_06310_));
 sky130_fd_sc_hd__nor2_1 _06770_ (.A(reg1_val[5]),
    .B(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__and2_1 _06771_ (.A(reg1_val[5]),
    .B(_06310_),
    .X(_06312_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(reg1_val[5]),
    .B(_06310_),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_1 _06773_ (.A(_06311_),
    .B(_06312_),
    .Y(_06314_));
 sky130_fd_sc_hd__or2_1 _06774_ (.A(_06311_),
    .B(_06312_),
    .X(_06315_));
 sky130_fd_sc_hd__and2_1 _06775_ (.A(reg2_val[4]),
    .B(net268),
    .X(_06316_));
 sky130_fd_sc_hd__a31o_1 _06776_ (.A1(net271),
    .A2(net252),
    .A3(_05528_),
    .B1(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__a31oi_4 _06777_ (.A1(net271),
    .A2(net252),
    .A3(_05528_),
    .B1(_06316_),
    .Y(_06318_));
 sky130_fd_sc_hd__or2_1 _06778_ (.A(reg1_val[4]),
    .B(net222),
    .X(_06319_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(reg1_val[4]),
    .B(net222),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_2 _06780_ (.A(_06319_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__and2_1 _06781_ (.A(reg2_val[3]),
    .B(net268),
    .X(_06322_));
 sky130_fd_sc_hd__a31oi_4 _06782_ (.A1(net271),
    .A2(net252),
    .A3(_05681_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__a31o_4 _06783_ (.A1(net271),
    .A2(net252),
    .A3(_05681_),
    .B1(_06322_),
    .X(_06324_));
 sky130_fd_sc_hd__nor2_1 _06784_ (.A(reg1_val[3]),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__or2_1 _06785_ (.A(reg1_val[3]),
    .B(_06324_),
    .X(_06326_));
 sky130_fd_sc_hd__and2_1 _06786_ (.A(reg1_val[3]),
    .B(_06324_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_1 _06787_ (.A(_06325_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__and2_1 _06788_ (.A(reg2_val[2]),
    .B(net268),
    .X(_06329_));
 sky130_fd_sc_hd__a31oi_4 _06789_ (.A1(net271),
    .A2(net252),
    .A3(_05738_),
    .B1(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a31o_1 _06790_ (.A1(net271),
    .A2(net252),
    .A3(_05738_),
    .B1(_06329_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(reg1_val[2]),
    .B(net216),
    .Y(_06332_));
 sky130_fd_sc_hd__or2_2 _06792_ (.A(reg1_val[2]),
    .B(net216),
    .X(_06333_));
 sky130_fd_sc_hd__nand2_2 _06793_ (.A(_06332_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__and2_1 _06794_ (.A(reg2_val[1]),
    .B(net268),
    .X(_06335_));
 sky130_fd_sc_hd__a31oi_4 _06795_ (.A1(net271),
    .A2(net252),
    .A3(_05811_),
    .B1(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__a31o_1 _06796_ (.A1(net271),
    .A2(net252),
    .A3(_05811_),
    .B1(_06335_),
    .X(_06337_));
 sky130_fd_sc_hd__or2_1 _06797_ (.A(net289),
    .B(net212),
    .X(_06338_));
 sky130_fd_sc_hd__xnor2_2 _06798_ (.A(net289),
    .B(net213),
    .Y(_06339_));
 sky130_fd_sc_hd__and2_1 _06799_ (.A(net271),
    .B(_05865_),
    .X(_06340_));
 sky130_fd_sc_hd__a22oi_4 _06800_ (.A1(reg2_val[0]),
    .A2(net268),
    .B1(net252),
    .B2(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__a22o_1 _06801_ (.A1(reg2_val[0]),
    .A2(net268),
    .B1(net252),
    .B2(_06340_),
    .X(_06342_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(net287),
    .B(net206),
    .Y(_06343_));
 sky130_fd_sc_hd__and2_1 _06803_ (.A(net289),
    .B(_06336_),
    .X(_06344_));
 sky130_fd_sc_hd__a21o_1 _06804_ (.A1(_06339_),
    .A2(_06343_),
    .B1(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__and2_1 _06805_ (.A(reg1_val[2]),
    .B(_06330_),
    .X(_06346_));
 sky130_fd_sc_hd__a21oi_1 _06806_ (.A1(_06334_),
    .A2(_06345_),
    .B1(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(reg1_val[3]),
    .B(net219),
    .Y(_06348_));
 sky130_fd_sc_hd__o21ai_1 _06808_ (.A1(_06328_),
    .A2(_06347_),
    .B1(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__and2_1 _06809_ (.A(reg1_val[4]),
    .B(_06318_),
    .X(_06350_));
 sky130_fd_sc_hd__a21oi_1 _06810_ (.A1(_06321_),
    .A2(_06349_),
    .B1(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(reg1_val[5]),
    .B(_06309_),
    .Y(_06352_));
 sky130_fd_sc_hd__o21a_1 _06812_ (.A1(_06314_),
    .A2(_06351_),
    .B1(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nand2b_1 _06813_ (.A_N(_06302_),
    .B(reg1_val[6]),
    .Y(_06354_));
 sky130_fd_sc_hd__o21ai_1 _06814_ (.A1(_06306_),
    .A2(_06353_),
    .B1(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__and2b_1 _06815_ (.A_N(_06285_),
    .B(reg1_val[7]),
    .X(_06356_));
 sky130_fd_sc_hd__a21o_1 _06816_ (.A1(_06300_),
    .A2(_06355_),
    .B1(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__and2b_1 _06817_ (.A_N(_06241_),
    .B(reg1_val[8]),
    .X(_06358_));
 sky130_fd_sc_hd__a21o_1 _06818_ (.A1(_06267_),
    .A2(_06357_),
    .B1(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__and2_1 _06819_ (.A(reg1_val[9]),
    .B(_06196_),
    .X(_06360_));
 sky130_fd_sc_hd__a21oi_1 _06820_ (.A1(_06223_),
    .A2(_06359_),
    .B1(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__and2b_1 _06821_ (.A_N(_06148_),
    .B(reg1_val[10]),
    .X(_06362_));
 sky130_fd_sc_hd__o21ba_1 _06822_ (.A1(_06169_),
    .A2(_06361_),
    .B1_N(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__and2b_1 _06823_ (.A_N(_06118_),
    .B(reg1_val[11]),
    .X(_06364_));
 sky130_fd_sc_hd__o21bai_1 _06824_ (.A1(_06136_),
    .A2(_06363_),
    .B1_N(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__and2b_1 _06825_ (.A_N(_06081_),
    .B(reg1_val[12]),
    .X(_06366_));
 sky130_fd_sc_hd__a21oi_1 _06826_ (.A1(_06106_),
    .A2(_06365_),
    .B1(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__and2b_1 _06827_ (.A_N(_06026_),
    .B(reg1_val[13]),
    .X(_06368_));
 sky130_fd_sc_hd__o21bai_1 _06828_ (.A1(_06059_),
    .A2(_06367_),
    .B1_N(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__and2b_1 _06829_ (.A_N(_05965_),
    .B(net291),
    .X(_06370_));
 sky130_fd_sc_hd__a21oi_1 _06830_ (.A1(_06004_),
    .A2(_06369_),
    .B1(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__and2b_1 _06831_ (.A_N(_05935_),
    .B(net290),
    .X(_06372_));
 sky130_fd_sc_hd__o21bai_1 _06832_ (.A1(_05953_),
    .A2(_06371_),
    .B1_N(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__and2_1 _06833_ (.A(reg1_val[16]),
    .B(_05883_),
    .X(_06374_));
 sky130_fd_sc_hd__a21o_1 _06834_ (.A1(_05919_),
    .A2(_06373_),
    .B1(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__and2_1 _06835_ (.A(reg1_val[17]),
    .B(_05829_),
    .X(_06376_));
 sky130_fd_sc_hd__a21o_1 _06836_ (.A1(_05857_),
    .A2(_06375_),
    .B1(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__and2_1 _06837_ (.A(reg1_val[18]),
    .B(_05757_),
    .X(_06378_));
 sky130_fd_sc_hd__a21o_1 _06838_ (.A1(_05802_),
    .A2(_06377_),
    .B1(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__and2_1 _06839_ (.A(reg1_val[19]),
    .B(_05700_),
    .X(_06380_));
 sky130_fd_sc_hd__a21oi_2 _06840_ (.A1(_05728_),
    .A2(_06379_),
    .B1(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(reg1_val[21]),
    .B(_05614_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _06842_ (.A(reg1_val[20]),
    .B(_05550_),
    .Y(_06383_));
 sky130_fd_sc_hd__o21a_1 _06843_ (.A1(_05652_),
    .A2(_06383_),
    .B1(_06382_),
    .X(_06384_));
 sky130_fd_sc_hd__nand2_1 _06844_ (.A(reg1_val[22]),
    .B(_05474_),
    .Y(_06385_));
 sky130_fd_sc_hd__o21a_1 _06845_ (.A1(_05518_),
    .A2(_06384_),
    .B1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__nand2_1 _06846_ (.A(reg1_val[23]),
    .B(_05410_),
    .Y(_06387_));
 sky130_fd_sc_hd__o221ai_4 _06847_ (.A1(_05671_),
    .A2(_06381_),
    .B1(_06386_),
    .B2(_05442_),
    .C1(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__and2b_1 _06848_ (.A_N(_05377_),
    .B(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(reg1_val[30]),
    .B(_04964_),
    .Y(_06390_));
 sky130_fd_sc_hd__and2_1 _06850_ (.A(reg1_val[29]),
    .B(_04801_),
    .X(_06391_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(reg1_val[28]),
    .B(_04888_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(reg1_val[27]),
    .B(_05040_),
    .Y(_06393_));
 sky130_fd_sc_hd__and2_1 _06853_ (.A(reg1_val[26]),
    .B(_05312_),
    .X(_06394_));
 sky130_fd_sc_hd__and2_1 _06854_ (.A(reg1_val[25]),
    .B(_05116_),
    .X(_06395_));
 sky130_fd_sc_hd__and2_1 _06855_ (.A(reg1_val[24]),
    .B(_05182_),
    .X(_06396_));
 sky130_fd_sc_hd__a21o_1 _06856_ (.A1(_05149_),
    .A2(_06396_),
    .B1(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__a21o_1 _06857_ (.A1(_05355_),
    .A2(_06397_),
    .B1(_06394_),
    .X(_06398_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(_05073_),
    .B(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__a21o_1 _06859_ (.A1(_06393_),
    .A2(_06399_),
    .B1(_04931_),
    .X(_06400_));
 sky130_fd_sc_hd__a21oi_1 _06860_ (.A1(_06392_),
    .A2(_06400_),
    .B1(_04844_),
    .Y(_06401_));
 sky130_fd_sc_hd__o21ai_1 _06861_ (.A1(_06391_),
    .A2(_06401_),
    .B1(_05008_),
    .Y(_06402_));
 sky130_fd_sc_hd__a21oi_1 _06862_ (.A1(_06390_),
    .A2(_06402_),
    .B1(_05269_),
    .Y(_06403_));
 sky130_fd_sc_hd__or2_1 _06863_ (.A(_04427_),
    .B(_05258_),
    .X(_06404_));
 sky130_fd_sc_hd__or4b_1 _06864_ (.A(instruction[6]),
    .B(_06389_),
    .C(_06403_),
    .D_N(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__a21o_1 _06865_ (.A1(_05225_),
    .A2(_06388_),
    .B1(_06396_),
    .X(_06406_));
 sky130_fd_sc_hd__a21o_1 _06866_ (.A1(_05149_),
    .A2(_06406_),
    .B1(_06395_),
    .X(_06407_));
 sky130_fd_sc_hd__a21o_1 _06867_ (.A1(_05355_),
    .A2(_06407_),
    .B1(_06394_),
    .X(_06408_));
 sky130_fd_sc_hd__a21boi_1 _06868_ (.A1(_05073_),
    .A2(_06408_),
    .B1_N(_06393_),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ai_1 _06869_ (.A1(_04931_),
    .A2(_06409_),
    .B1(_06392_),
    .Y(_06410_));
 sky130_fd_sc_hd__a21o_1 _06870_ (.A1(_04855_),
    .A2(_06410_),
    .B1(_06391_),
    .X(_06411_));
 sky130_fd_sc_hd__a21bo_1 _06871_ (.A1(_05008_),
    .A2(_06411_),
    .B1_N(_06390_),
    .X(_06412_));
 sky130_fd_sc_hd__o21ai_1 _06872_ (.A1(_05269_),
    .A2(_06412_),
    .B1(_06404_),
    .Y(_06413_));
 sky130_fd_sc_hd__a21bo_1 _06873_ (.A1(instruction[6]),
    .A2(_06413_),
    .B1_N(_06405_),
    .X(_06414_));
 sky130_fd_sc_hd__or2_4 _06874_ (.A(instruction[3]),
    .B(instruction[4]),
    .X(_06415_));
 sky130_fd_sc_hd__nor2_2 _06875_ (.A(net287),
    .B(net209),
    .Y(_06416_));
 sky130_fd_sc_hd__nor2_1 _06876_ (.A(net293),
    .B(net206),
    .Y(_06417_));
 sky130_fd_sc_hd__and4_1 _06877_ (.A(_05728_),
    .B(_05802_),
    .C(_05857_),
    .D(_05919_),
    .X(_06418_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(_06223_),
    .B(_06300_),
    .Y(_06419_));
 sky130_fd_sc_hd__or4_1 _06879_ (.A(_05953_),
    .B(_05993_),
    .C(_06059_),
    .D(_06100_),
    .X(_06420_));
 sky130_fd_sc_hd__or4_1 _06880_ (.A(_06136_),
    .B(_06169_),
    .C(_06419_),
    .D(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__o211a_1 _06881_ (.A1(_06304_),
    .A2(_06305_),
    .B1(_06315_),
    .C1(_06321_),
    .X(_06422_));
 sky130_fd_sc_hd__o2111a_1 _06882_ (.A1(_06416_),
    .A2(_06417_),
    .B1(_06267_),
    .C1(_06334_),
    .D1(_06339_),
    .X(_06423_));
 sky130_fd_sc_hd__and4bb_1 _06883_ (.A_N(_06328_),
    .B_N(_06421_),
    .C(_06422_),
    .D(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__and4b_1 _06884_ (.A_N(_05377_),
    .B(_05662_),
    .C(_06418_),
    .D(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__a21oi_1 _06885_ (.A1(instruction[6]),
    .A2(_05269_),
    .B1(_06415_),
    .Y(_06426_));
 sky130_fd_sc_hd__o21a_1 _06886_ (.A1(instruction[6]),
    .A2(_06425_),
    .B1(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__nand2_2 _06887_ (.A(instruction[3]),
    .B(instruction[4]),
    .Y(_06428_));
 sky130_fd_sc_hd__inv_2 _06888_ (.A(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__or2_2 _06889_ (.A(_04394_),
    .B(instruction[4]),
    .X(_06430_));
 sky130_fd_sc_hd__a221o_2 _06890_ (.A1(instruction[3]),
    .A2(_06414_),
    .B1(_06425_),
    .B2(_06429_),
    .C1(_06427_),
    .X(_06431_));
 sky130_fd_sc_hd__xor2_4 _06891_ (.A(instruction[5]),
    .B(_06431_),
    .X(dest_pred_val));
 sky130_fd_sc_hd__and3_1 _06892_ (.A(instruction[2]),
    .B(_04459_),
    .C(_04470_),
    .X(_06432_));
 sky130_fd_sc_hd__nand3_4 _06893_ (.A(instruction[2]),
    .B(_04459_),
    .C(_04470_),
    .Y(_06433_));
 sky130_fd_sc_hd__a21o_4 _06894_ (.A1(_04492_),
    .A2(dest_pred_val),
    .B1(net249),
    .X(take_branch));
 sky130_fd_sc_hd__and4_1 _06895_ (.A(reg1_idx[3]),
    .B(reg1_idx[0]),
    .C(reg1_idx[1]),
    .D(reg1_idx[4]),
    .X(_06434_));
 sky130_fd_sc_hd__and3_4 _06896_ (.A(reg1_idx[2]),
    .B(net249),
    .C(_06434_),
    .X(int_return));
 sky130_fd_sc_hd__a21oi_2 _06897_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(instruction[4]),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2b_4 _06898_ (.A_N(instruction[5]),
    .B(instruction[6]),
    .Y(_06436_));
 sky130_fd_sc_hd__a221oi_4 _06899_ (.A1(net270),
    .A2(_04692_),
    .B1(_06436_),
    .B2(instruction[4]),
    .C1(_06435_),
    .Y(_06437_));
 sky130_fd_sc_hd__a221o_1 _06900_ (.A1(net270),
    .A2(_04692_),
    .B1(_06436_),
    .B2(instruction[4]),
    .C1(_06435_),
    .X(_06438_));
 sky130_fd_sc_hd__nor2_2 _06901_ (.A(net260),
    .B(_06437_),
    .Y(_06439_));
 sky130_fd_sc_hd__nand2_2 _06902_ (.A(_04383_),
    .B(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_8 _06903_ (.A(div_complete),
    .B(net204),
    .Y(busy));
 sky130_fd_sc_hd__and4b_4 _06904_ (.A_N(instruction[2]),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06441_));
 sky130_fd_sc_hd__and2_4 _06905_ (.A(instruction[11]),
    .B(_06441_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _06906_ (.A(instruction[12]),
    .B(_06441_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _06907_ (.A(instruction[13]),
    .B(_06441_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or3_2 _06908_ (.A(net272),
    .B(_04681_),
    .C(net249),
    .X(_06442_));
 sky130_fd_sc_hd__and2_4 _06909_ (.A(instruction[11]),
    .B(_06442_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _06910_ (.A(instruction[12]),
    .B(_06442_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _06911_ (.A(instruction[13]),
    .B(_06442_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _06912_ (.A(instruction[14]),
    .B(_06442_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _06913_ (.A(instruction[15]),
    .B(_06442_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__or2_1 _06914_ (.A(instruction[25]),
    .B(_04492_),
    .X(_06443_));
 sky130_fd_sc_hd__o211a_4 _06915_ (.A1(instruction[18]),
    .A2(_04503_),
    .B1(_06443_),
    .C1(net273),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__or2_1 _06916_ (.A(instruction[26]),
    .B(_04492_),
    .X(_06444_));
 sky130_fd_sc_hd__o211a_4 _06917_ (.A1(instruction[19]),
    .A2(_04503_),
    .B1(_06444_),
    .C1(net273),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__or2_1 _06918_ (.A(instruction[27]),
    .B(_04492_),
    .X(_06445_));
 sky130_fd_sc_hd__o211a_4 _06919_ (.A1(instruction[20]),
    .A2(_04503_),
    .B1(_06445_),
    .C1(net273),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__or2_1 _06920_ (.A(instruction[28]),
    .B(_04492_),
    .X(_06446_));
 sky130_fd_sc_hd__o211a_4 _06921_ (.A1(instruction[21]),
    .A2(_04503_),
    .B1(_06446_),
    .C1(net273),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__or2_1 _06922_ (.A(instruction[29]),
    .B(_04492_),
    .X(_06447_));
 sky130_fd_sc_hd__o211a_4 _06923_ (.A1(instruction[22]),
    .A2(_04503_),
    .B1(_06447_),
    .C1(net273),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__nor3_2 _06924_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06430_),
    .Y(_06448_));
 sky130_fd_sc_hd__or3_4 _06925_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06430_),
    .X(_06449_));
 sky130_fd_sc_hd__or2_4 _06926_ (.A(instruction[6]),
    .B(instruction[5]),
    .X(_06450_));
 sky130_fd_sc_hd__nand2_4 _06927_ (.A(_04394_),
    .B(instruction[4]),
    .Y(_06451_));
 sky130_fd_sc_hd__nor2_2 _06928_ (.A(_06450_),
    .B(_06451_),
    .Y(_06452_));
 sky130_fd_sc_hd__or2_2 _06929_ (.A(_06450_),
    .B(_06451_),
    .X(_06453_));
 sky130_fd_sc_hd__a31o_1 _06930_ (.A1(instruction[17]),
    .A2(net196),
    .A3(_06453_),
    .B1(net270),
    .X(_06454_));
 sky130_fd_sc_hd__nor2_1 _06931_ (.A(instruction[6]),
    .B(is_load),
    .Y(_06455_));
 sky130_fd_sc_hd__o211a_1 _06932_ (.A1(instruction[40]),
    .A2(_04692_),
    .B1(_06454_),
    .C1(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__a32o_2 _06933_ (.A1(instruction[24]),
    .A2(instruction[7]),
    .A3(is_load),
    .B1(_04736_),
    .B2(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__nand2_8 _06934_ (.A(net247),
    .B(_06457_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a22o_2 _06935_ (.A1(instruction[7]),
    .A2(is_load),
    .B1(net253),
    .B2(_06456_),
    .X(_06458_));
 sky130_fd_sc_hd__nand2_8 _06936_ (.A(net247),
    .B(_06458_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__nand2b_4 _06937_ (.A_N(instruction[6]),
    .B(instruction[5]),
    .Y(_06459_));
 sky130_fd_sc_hd__nor3_2 _06938_ (.A(net284),
    .B(_06415_),
    .C(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__or3_2 _06939_ (.A(net284),
    .B(_06415_),
    .C(_06459_),
    .X(_06461_));
 sky130_fd_sc_hd__nand2_1 _06940_ (.A(net206),
    .B(net242),
    .Y(_06462_));
 sky130_fd_sc_hd__a21o_2 _06941_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(net242),
    .X(_06463_));
 sky130_fd_sc_hd__nor2_4 _06942_ (.A(net286),
    .B(_05279_),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_2 _06943_ (.A(net294),
    .B(_05269_),
    .Y(_06465_));
 sky130_fd_sc_hd__and2_1 _06944_ (.A(reg1_val[31]),
    .B(net295),
    .X(_06466_));
 sky130_fd_sc_hd__and3_4 _06945_ (.A(net292),
    .B(reg1_val[31]),
    .C(net294),
    .X(_06467_));
 sky130_fd_sc_hd__xor2_4 _06946_ (.A(net289),
    .B(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__xnor2_4 _06947_ (.A(net289),
    .B(_06467_),
    .Y(_06469_));
 sky130_fd_sc_hd__and2_2 _06948_ (.A(net295),
    .B(_05258_),
    .X(_06470_));
 sky130_fd_sc_hd__nand2_2 _06949_ (.A(net295),
    .B(_05258_),
    .Y(_06471_));
 sky130_fd_sc_hd__and4_1 _06950_ (.A(_06323_),
    .B(_06330_),
    .C(_06336_),
    .D(net210),
    .X(_06472_));
 sky130_fd_sc_hd__or4_4 _06951_ (.A(_06324_),
    .B(net216),
    .C(net213),
    .D(net208),
    .X(_06473_));
 sky130_fd_sc_hd__or4_4 _06952_ (.A(_06285_),
    .B(_06302_),
    .C(_06310_),
    .D(net222),
    .X(_06474_));
 sky130_fd_sc_hd__nor2_4 _06953_ (.A(_06473_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__or2_1 _06954_ (.A(_06473_),
    .B(_06474_),
    .X(_06476_));
 sky130_fd_sc_hd__or2_4 _06955_ (.A(_06187_),
    .B(_06241_),
    .X(_06477_));
 sky130_fd_sc_hd__or2_1 _06956_ (.A(_06118_),
    .B(_06148_),
    .X(_06478_));
 sky130_fd_sc_hd__or4_2 _06957_ (.A(_06026_),
    .B(_06081_),
    .C(_06118_),
    .D(_06148_),
    .X(_06479_));
 sky130_fd_sc_hd__nor4_4 _06958_ (.A(_05935_),
    .B(_05965_),
    .C(_06477_),
    .D(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_1 _06959_ (.A(_06475_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__and2_1 _06960_ (.A(_05829_),
    .B(_05883_),
    .X(_06482_));
 sky130_fd_sc_hd__and4_1 _06961_ (.A(_05700_),
    .B(_05757_),
    .C(_05829_),
    .D(_05883_),
    .X(_06483_));
 sky130_fd_sc_hd__and3_4 _06962_ (.A(_06475_),
    .B(_06480_),
    .C(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__nand3_4 _06963_ (.A(_06475_),
    .B(_06480_),
    .C(_06483_),
    .Y(_06485_));
 sky130_fd_sc_hd__and2_2 _06964_ (.A(_05550_),
    .B(_05614_),
    .X(_06486_));
 sky130_fd_sc_hd__and3_1 _06965_ (.A(_05410_),
    .B(_05474_),
    .C(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__nand3_2 _06966_ (.A(_05410_),
    .B(_05474_),
    .C(_06486_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(_06484_),
    .B(_06487_),
    .Y(_06489_));
 sky130_fd_sc_hd__and2_1 _06968_ (.A(_05116_),
    .B(_05182_),
    .X(_06490_));
 sky130_fd_sc_hd__a31o_2 _06969_ (.A1(_06484_),
    .A2(_06487_),
    .A3(_06490_),
    .B1(net174),
    .X(_06491_));
 sky130_fd_sc_hd__xor2_4 _06970_ (.A(_05312_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__xnor2_1 _06971_ (.A(_05312_),
    .B(_06491_),
    .Y(_06493_));
 sky130_fd_sc_hd__and2_4 _06972_ (.A(net288),
    .B(net289),
    .X(_06494_));
 sky130_fd_sc_hd__nand2_4 _06973_ (.A(net288),
    .B(net289),
    .Y(_06495_));
 sky130_fd_sc_hd__a21o_1 _06974_ (.A1(_06484_),
    .A2(_06487_),
    .B1(net174),
    .X(_06496_));
 sky130_fd_sc_hd__nor2_1 _06975_ (.A(_05182_),
    .B(net174),
    .Y(_06497_));
 sky130_fd_sc_hd__a31o_2 _06976_ (.A1(_05182_),
    .A2(_06484_),
    .A3(_06487_),
    .B1(net174),
    .X(_06498_));
 sky130_fd_sc_hd__xnor2_2 _06977_ (.A(_05116_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__xor2_4 _06978_ (.A(_05116_),
    .B(_06498_),
    .X(_06500_));
 sky130_fd_sc_hd__o22a_1 _06979_ (.A1(net288),
    .A2(net67),
    .B1(net237),
    .B2(net64),
    .X(_06501_));
 sky130_fd_sc_hd__xnor2_2 _06980_ (.A(net239),
    .B(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__or4_2 _06981_ (.A(net292),
    .B(net289),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06503_));
 sky130_fd_sc_hd__nand2_1 _06982_ (.A(net263),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__o21a_1 _06983_ (.A1(reg1_val[4]),
    .A2(_06503_),
    .B1(net263),
    .X(_06505_));
 sky130_fd_sc_hd__xnor2_2 _06984_ (.A(reg1_val[5]),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__inv_4 _06985_ (.A(net194),
    .Y(_06507_));
 sky130_fd_sc_hd__o31a_1 _06986_ (.A1(net292),
    .A2(net289),
    .A3(reg1_val[2]),
    .B1(net263),
    .X(_06508_));
 sky130_fd_sc_hd__xnor2_1 _06987_ (.A(reg1_val[3]),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__xor2_2 _06988_ (.A(reg1_val[4]),
    .B(_06504_),
    .X(_06510_));
 sky130_fd_sc_hd__or2_1 _06989_ (.A(net192),
    .B(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(net192),
    .B(_06510_),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(_06511_),
    .B(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__a21o_2 _06992_ (.A1(_06484_),
    .A2(_06486_),
    .B1(net174),
    .X(_06514_));
 sky130_fd_sc_hd__xnor2_4 _06993_ (.A(_05485_),
    .B(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__xnor2_4 _06994_ (.A(_05474_),
    .B(_06514_),
    .Y(_06516_));
 sky130_fd_sc_hd__mux2_2 _06995_ (.A0(_06511_),
    .A1(_06512_),
    .S(_06507_),
    .X(_06517_));
 sky130_fd_sc_hd__nor2_1 _06996_ (.A(_05550_),
    .B(net174),
    .Y(_06518_));
 sky130_fd_sc_hd__a211o_2 _06997_ (.A1(_05550_),
    .A2(_06484_),
    .B1(net174),
    .C1(_05623_),
    .X(_06519_));
 sky130_fd_sc_hd__a211o_2 _06998_ (.A1(net175),
    .A2(_06485_),
    .B1(_06518_),
    .C1(_05614_),
    .X(_06520_));
 sky130_fd_sc_hd__and2_2 _06999_ (.A(_06519_),
    .B(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__nand2_8 _07000_ (.A(_06519_),
    .B(_06520_),
    .Y(_06522_));
 sky130_fd_sc_hd__o22a_1 _07001_ (.A1(net155),
    .A2(net62),
    .B1(net153),
    .B2(net60),
    .X(_06523_));
 sky130_fd_sc_hd__xnor2_1 _07002_ (.A(net194),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__or2_1 _07003_ (.A(_06502_),
    .B(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__o21a_1 _07004_ (.A1(net292),
    .A2(reg1_val[1]),
    .B1(net263),
    .X(_06526_));
 sky130_fd_sc_hd__xnor2_2 _07005_ (.A(reg1_val[2]),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__and2_1 _07006_ (.A(_06469_),
    .B(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _07007_ (.A(_06469_),
    .B(_06527_),
    .Y(_06529_));
 sky130_fd_sc_hd__nor2_1 _07008_ (.A(_06469_),
    .B(_06527_),
    .Y(_06530_));
 sky130_fd_sc_hd__or2_1 _07009_ (.A(_06469_),
    .B(_06527_),
    .X(_06531_));
 sky130_fd_sc_hd__nor2_2 _07010_ (.A(_06528_),
    .B(_06530_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand2_1 _07011_ (.A(_06529_),
    .B(_06531_),
    .Y(_06533_));
 sky130_fd_sc_hd__a22oi_4 _07012_ (.A1(_05182_),
    .A2(_06496_),
    .B1(_06497_),
    .B2(_06489_),
    .Y(_06534_));
 sky130_fd_sc_hd__a22o_2 _07013_ (.A1(_05182_),
    .A2(_06496_),
    .B1(_06497_),
    .B2(_06489_),
    .X(_06535_));
 sky130_fd_sc_hd__a31oi_4 _07014_ (.A1(_05474_),
    .A2(_06484_),
    .A3(_06486_),
    .B1(net174),
    .Y(_06536_));
 sky130_fd_sc_hd__xor2_4 _07015_ (.A(_05410_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__xnor2_4 _07016_ (.A(_05410_),
    .B(_06536_),
    .Y(_06538_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(_06529_),
    .A1(_06531_),
    .S(net192),
    .X(_06539_));
 sky130_fd_sc_hd__mux2_2 _07018_ (.A0(_06528_),
    .A1(_06530_),
    .S(net192),
    .X(_06540_));
 sky130_fd_sc_hd__o22a_1 _07019_ (.A1(net151),
    .A2(net58),
    .B1(net56),
    .B2(net148),
    .X(_06541_));
 sky130_fd_sc_hd__xnor2_2 _07020_ (.A(net193),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__xnor2_2 _07021_ (.A(_06502_),
    .B(_06524_),
    .Y(_06543_));
 sky130_fd_sc_hd__o21a_1 _07022_ (.A1(_06542_),
    .A2(_06543_),
    .B1(_06525_),
    .X(_06544_));
 sky130_fd_sc_hd__o22a_1 _07023_ (.A1(net64),
    .A2(net151),
    .B1(net58),
    .B2(net149),
    .X(_06545_));
 sky130_fd_sc_hd__xnor2_2 _07024_ (.A(net193),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__a41o_1 _07025_ (.A1(_05312_),
    .A2(_06484_),
    .A3(_06487_),
    .A4(_06490_),
    .B1(_05040_),
    .X(_06547_));
 sky130_fd_sc_hd__nand3_2 _07026_ (.A(_05040_),
    .B(_05312_),
    .C(_06490_),
    .Y(_06548_));
 sky130_fd_sc_hd__nor3_4 _07027_ (.A(_06485_),
    .B(_06488_),
    .C(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__or3_4 _07028_ (.A(_06485_),
    .B(_06488_),
    .C(_06548_),
    .X(_06550_));
 sky130_fd_sc_hd__nor2_1 _07029_ (.A(_05040_),
    .B(net175),
    .Y(_06551_));
 sky130_fd_sc_hd__a31oi_2 _07030_ (.A1(net175),
    .A2(_06547_),
    .A3(_06550_),
    .B1(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__a31o_4 _07031_ (.A1(net175),
    .A2(_06547_),
    .A3(_06550_),
    .B1(_06551_),
    .X(_06553_));
 sky130_fd_sc_hd__o22a_1 _07032_ (.A1(net67),
    .A2(net237),
    .B1(net55),
    .B2(net288),
    .X(_06554_));
 sky130_fd_sc_hd__xnor2_2 _07033_ (.A(net239),
    .B(_06554_),
    .Y(_06555_));
 sky130_fd_sc_hd__o22a_1 _07034_ (.A1(net62),
    .A2(net153),
    .B1(net56),
    .B2(net155),
    .X(_06556_));
 sky130_fd_sc_hd__xnor2_2 _07035_ (.A(net194),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__nor2_1 _07036_ (.A(_06555_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__xnor2_2 _07037_ (.A(_06555_),
    .B(_06557_),
    .Y(_06559_));
 sky130_fd_sc_hd__nor2_1 _07038_ (.A(_06546_),
    .B(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__xor2_2 _07039_ (.A(_06546_),
    .B(_06559_),
    .X(_00136_));
 sky130_fd_sc_hd__nand2b_1 _07040_ (.A_N(_06544_),
    .B(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__or2_1 _07041_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .X(_00138_));
 sky130_fd_sc_hd__o31a_2 _07042_ (.A1(reg1_val[6]),
    .A2(_06503_),
    .A3(_00138_),
    .B1(net263),
    .X(_00139_));
 sky130_fd_sc_hd__xnor2_4 _07043_ (.A(reg1_val[7]),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__o21a_1 _07044_ (.A1(_06503_),
    .A2(_00138_),
    .B1(net263),
    .X(_00141_));
 sky130_fd_sc_hd__xnor2_2 _07045_ (.A(reg1_val[6]),
    .B(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_2 _07046_ (.A(net194),
    .B(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__or2_1 _07047_ (.A(net194),
    .B(_00142_),
    .X(_00144_));
 sky130_fd_sc_hd__nand2_4 _07048_ (.A(_00143_),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__o21ai_4 _07049_ (.A1(_06471_),
    .A2(_06484_),
    .B1(_05550_),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_2 _07050_ (.A(_06485_),
    .B(_06518_),
    .Y(_00147_));
 sky130_fd_sc_hd__and2_4 _07051_ (.A(_00146_),
    .B(_00147_),
    .X(_00148_));
 sky130_fd_sc_hd__nand2_4 _07052_ (.A(_00146_),
    .B(_00147_),
    .Y(_00149_));
 sky130_fd_sc_hd__or3b_1 _07053_ (.A(net194),
    .B(_00142_),
    .C_N(net190),
    .X(_00150_));
 sky130_fd_sc_hd__o21a_2 _07054_ (.A1(net189),
    .A2(_00143_),
    .B1(_00150_),
    .X(_00151_));
 sky130_fd_sc_hd__a31oi_4 _07055_ (.A1(_06475_),
    .A2(_06480_),
    .A3(_06482_),
    .B1(net174),
    .Y(_00152_));
 sky130_fd_sc_hd__nor2_1 _07056_ (.A(_05757_),
    .B(net174),
    .Y(_00153_));
 sky130_fd_sc_hd__o21ai_4 _07057_ (.A1(_00152_),
    .A2(_00153_),
    .B1(_05700_),
    .Y(_00154_));
 sky130_fd_sc_hd__or3_4 _07058_ (.A(_05700_),
    .B(_00152_),
    .C(_00153_),
    .X(_00155_));
 sky130_fd_sc_hd__and2_2 _07059_ (.A(_00154_),
    .B(_00155_),
    .X(_00156_));
 sky130_fd_sc_hd__nand2_8 _07060_ (.A(_00154_),
    .B(_00155_),
    .Y(_00157_));
 sky130_fd_sc_hd__o22a_1 _07061_ (.A1(net147),
    .A2(net52),
    .B1(net145),
    .B2(net50),
    .X(_00158_));
 sky130_fd_sc_hd__xnor2_1 _07062_ (.A(net189),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__or4_2 _07063_ (.A(reg1_val[6]),
    .B(reg1_val[7]),
    .C(_06503_),
    .D(_00138_),
    .X(_00160_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(net263),
    .B(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__o21a_1 _07065_ (.A1(reg1_val[8]),
    .A2(_00160_),
    .B1(net263),
    .X(_00162_));
 sky130_fd_sc_hd__xnor2_4 _07066_ (.A(reg1_val[9]),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__xnor2_2 _07067_ (.A(_05757_),
    .B(_00152_),
    .Y(_00164_));
 sky130_fd_sc_hd__xnor2_4 _07068_ (.A(_05766_),
    .B(_00152_),
    .Y(_00165_));
 sky130_fd_sc_hd__xor2_2 _07069_ (.A(reg1_val[8]),
    .B(_00161_),
    .X(_00166_));
 sky130_fd_sc_hd__or2_1 _07070_ (.A(net190),
    .B(_00166_),
    .X(_00167_));
 sky130_fd_sc_hd__nand2_1 _07071_ (.A(net190),
    .B(_00166_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _07072_ (.A(_00167_),
    .B(_00168_),
    .Y(_00169_));
 sky130_fd_sc_hd__a21o_1 _07073_ (.A1(_06475_),
    .A2(_06480_),
    .B1(net174),
    .X(_00170_));
 sky130_fd_sc_hd__nor2_1 _07074_ (.A(_05883_),
    .B(net174),
    .Y(_00171_));
 sky130_fd_sc_hd__a31o_2 _07075_ (.A1(_05883_),
    .A2(_06475_),
    .A3(_06480_),
    .B1(net174),
    .X(_00172_));
 sky130_fd_sc_hd__xnor2_2 _07076_ (.A(_05829_),
    .B(_00172_),
    .Y(_00173_));
 sky130_fd_sc_hd__xor2_4 _07077_ (.A(_05829_),
    .B(_00172_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_2 _07078_ (.A0(_00168_),
    .A1(_00167_),
    .S(net172),
    .X(_00175_));
 sky130_fd_sc_hd__o22a_1 _07079_ (.A1(net100),
    .A2(net134),
    .B1(net98),
    .B2(net132),
    .X(_00176_));
 sky130_fd_sc_hd__xnor2_1 _07080_ (.A(net172),
    .B(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__nor2_1 _07081_ (.A(_00159_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__xnor2_1 _07082_ (.A(_06544_),
    .B(_00136_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(_00178_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_2 _07084_ (.A(_00137_),
    .B(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__or4_4 _07085_ (.A(reg1_val[8]),
    .B(reg1_val[9]),
    .C(reg1_val[10]),
    .D(_00160_),
    .X(_00182_));
 sky130_fd_sc_hd__or4_4 _07086_ (.A(reg1_val[11]),
    .B(reg1_val[12]),
    .C(reg1_val[13]),
    .D(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__or3_1 _07087_ (.A(net291),
    .B(net290),
    .C(_00183_),
    .X(_00184_));
 sky130_fd_sc_hd__or2_2 _07088_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_00185_));
 sky130_fd_sc_hd__or3_4 _07089_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_00185_),
    .X(_00186_));
 sky130_fd_sc_hd__o41a_4 _07090_ (.A1(net291),
    .A2(net290),
    .A3(_00183_),
    .A4(_00186_),
    .B1(net262),
    .X(_00187_));
 sky130_fd_sc_hd__or2_1 _07091_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .X(_00188_));
 sky130_fd_sc_hd__or2_1 _07092_ (.A(reg1_val[22]),
    .B(_00188_),
    .X(_00189_));
 sky130_fd_sc_hd__and2_1 _07093_ (.A(net263),
    .B(_00189_),
    .X(_00190_));
 sky130_fd_sc_hd__o21ai_1 _07094_ (.A1(_00187_),
    .A2(_00190_),
    .B1(reg1_val[23]),
    .Y(_00191_));
 sky130_fd_sc_hd__or3_1 _07095_ (.A(reg1_val[23]),
    .B(_00187_),
    .C(_00190_),
    .X(_00192_));
 sky130_fd_sc_hd__and2_2 _07096_ (.A(_00191_),
    .B(_00192_),
    .X(_00193_));
 sky130_fd_sc_hd__and3_1 _07097_ (.A(net294),
    .B(_05258_),
    .C(net222),
    .X(_00194_));
 sky130_fd_sc_hd__a211o_1 _07098_ (.A1(_06318_),
    .A2(_06472_),
    .B1(_06471_),
    .C1(_06310_),
    .X(_00195_));
 sky130_fd_sc_hd__a211o_1 _07099_ (.A1(net175),
    .A2(_06473_),
    .B1(_00194_),
    .C1(_06309_),
    .X(_00196_));
 sky130_fd_sc_hd__and2_1 _07100_ (.A(_00195_),
    .B(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__nand2_4 _07101_ (.A(_00195_),
    .B(_00196_),
    .Y(_00198_));
 sky130_fd_sc_hd__o311a_2 _07102_ (.A1(reg1_val[20]),
    .A2(_00184_),
    .A3(_00186_),
    .B1(reg1_val[21]),
    .C1(net262),
    .X(_00199_));
 sky130_fd_sc_hd__a211oi_4 _07103_ (.A1(reg1_val[20]),
    .A2(net262),
    .B1(_00187_),
    .C1(reg1_val[21]),
    .Y(_00200_));
 sky130_fd_sc_hd__nor2_4 _07104_ (.A(_00199_),
    .B(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _07105_ (.A(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__o311a_1 _07106_ (.A1(_00184_),
    .A2(_00186_),
    .A3(_00188_),
    .B1(net262),
    .C1(reg1_val[22]),
    .X(_00203_));
 sky130_fd_sc_hd__a211oi_2 _07107_ (.A1(net263),
    .A2(_00188_),
    .B1(_00187_),
    .C1(reg1_val[22]),
    .Y(_00204_));
 sky130_fd_sc_hd__nor2_1 _07108_ (.A(_00203_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__or4_2 _07109_ (.A(_00199_),
    .B(_00200_),
    .C(_00203_),
    .D(_00204_),
    .X(_00206_));
 sky130_fd_sc_hd__o22ai_2 _07110_ (.A1(_00199_),
    .A2(_00200_),
    .B1(_00203_),
    .B2(_00204_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_2 _07111_ (.A(_00206_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__a21o_1 _07112_ (.A1(net175),
    .A2(_06473_),
    .B1(net222),
    .X(_00209_));
 sky130_fd_sc_hd__nand2_1 _07113_ (.A(_06473_),
    .B(_00194_),
    .Y(_00210_));
 sky130_fd_sc_hd__and2_4 _07114_ (.A(_00209_),
    .B(_00210_),
    .X(_00211_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_00209_),
    .B(_00210_),
    .Y(_00212_));
 sky130_fd_sc_hd__nor2_1 _07116_ (.A(net95),
    .B(_00206_),
    .Y(_00213_));
 sky130_fd_sc_hd__mux2_1 _07117_ (.A0(_00206_),
    .A1(_00207_),
    .S(net95),
    .X(_00214_));
 sky130_fd_sc_hd__o22a_1 _07118_ (.A1(net130),
    .A2(net47),
    .B1(net127),
    .B2(net45),
    .X(_00215_));
 sky130_fd_sc_hd__xnor2_1 _07119_ (.A(net97),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__or3_4 _07120_ (.A(reg1_val[23]),
    .B(_00186_),
    .C(_00189_),
    .X(_00217_));
 sky130_fd_sc_hd__or4_4 _07121_ (.A(net291),
    .B(net290),
    .C(_00183_),
    .D(_00217_),
    .X(_00218_));
 sky130_fd_sc_hd__or2_2 _07122_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .X(_00219_));
 sky130_fd_sc_hd__or2_1 _07123_ (.A(_00217_),
    .B(_00219_),
    .X(_00220_));
 sky130_fd_sc_hd__o41a_1 _07124_ (.A1(net291),
    .A2(net290),
    .A3(_00183_),
    .A4(_00220_),
    .B1(net263),
    .X(_00221_));
 sky130_fd_sc_hd__a21oi_1 _07125_ (.A1(reg1_val[26]),
    .A2(net263),
    .B1(_00221_),
    .Y(_00222_));
 sky130_fd_sc_hd__xnor2_1 _07126_ (.A(reg1_val[27]),
    .B(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__and3_2 _07127_ (.A(net294),
    .B(_05258_),
    .C(net208),
    .X(_00224_));
 sky130_fd_sc_hd__xnor2_4 _07128_ (.A(_06336_),
    .B(_00224_),
    .Y(_00225_));
 sky130_fd_sc_hd__xnor2_1 _07129_ (.A(net213),
    .B(_00224_),
    .Y(_00226_));
 sky130_fd_sc_hd__o41a_1 _07130_ (.A1(net291),
    .A2(net290),
    .A3(_00183_),
    .A4(_00217_),
    .B1(net262),
    .X(_00227_));
 sky130_fd_sc_hd__o211ai_2 _07131_ (.A1(reg1_val[24]),
    .A2(_00218_),
    .B1(net262),
    .C1(reg1_val[25]),
    .Y(_00228_));
 sky130_fd_sc_hd__a211o_1 _07132_ (.A1(reg1_val[24]),
    .A2(net262),
    .B1(_00227_),
    .C1(reg1_val[25]),
    .X(_00229_));
 sky130_fd_sc_hd__and2_1 _07133_ (.A(_00228_),
    .B(_00229_),
    .X(_00230_));
 sky130_fd_sc_hd__xor2_2 _07134_ (.A(reg1_val[26]),
    .B(_00221_),
    .X(_00231_));
 sky130_fd_sc_hd__and3_1 _07135_ (.A(_00228_),
    .B(_00229_),
    .C(_00231_),
    .X(_00232_));
 sky130_fd_sc_hd__a21oi_1 _07136_ (.A1(_00228_),
    .A2(_00229_),
    .B1(_00231_),
    .Y(_00233_));
 sky130_fd_sc_hd__nor2_1 _07137_ (.A(_00232_),
    .B(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__and2b_1 _07138_ (.A_N(net93),
    .B(_00232_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _07139_ (.A0(_00232_),
    .A1(_00233_),
    .S(net93),
    .X(_00236_));
 sky130_fd_sc_hd__a22o_1 _07140_ (.A1(_00225_),
    .A2(net43),
    .B1(net41),
    .B2(net208),
    .X(_00237_));
 sky130_fd_sc_hd__xor2_1 _07141_ (.A(net94),
    .B(_00237_),
    .X(_00238_));
 sky130_fd_sc_hd__xor2_1 _07142_ (.A(_00216_),
    .B(_00238_),
    .X(_00239_));
 sky130_fd_sc_hd__o211a_4 _07143_ (.A1(net213),
    .A2(net208),
    .B1(net294),
    .C1(_05258_),
    .X(_00240_));
 sky130_fd_sc_hd__o311a_4 _07144_ (.A1(net216),
    .A2(net213),
    .A3(net208),
    .B1(_05258_),
    .C1(net294),
    .X(_00241_));
 sky130_fd_sc_hd__xnor2_4 _07145_ (.A(_06324_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__xnor2_4 _07146_ (.A(_06323_),
    .B(_00241_),
    .Y(_00243_));
 sky130_fd_sc_hd__xor2_2 _07147_ (.A(reg1_val[24]),
    .B(_00227_),
    .X(_00244_));
 sky130_fd_sc_hd__and3_1 _07148_ (.A(_00191_),
    .B(_00192_),
    .C(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__a21oi_1 _07149_ (.A1(_00191_),
    .A2(_00192_),
    .B1(_00244_),
    .Y(_00246_));
 sky130_fd_sc_hd__nor2_1 _07150_ (.A(_00245_),
    .B(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _07151_ (.A(net38),
    .Y(_00248_));
 sky130_fd_sc_hd__xnor2_4 _07152_ (.A(net216),
    .B(_00240_),
    .Y(_00249_));
 sky130_fd_sc_hd__xnor2_4 _07153_ (.A(_06330_),
    .B(_00240_),
    .Y(_00250_));
 sky130_fd_sc_hd__mux2_1 _07154_ (.A0(_00245_),
    .A1(_00246_),
    .S(net89),
    .X(_00251_));
 sky130_fd_sc_hd__inv_2 _07155_ (.A(net36),
    .Y(_00252_));
 sky130_fd_sc_hd__a22o_1 _07156_ (.A1(_00243_),
    .A2(net39),
    .B1(_00250_),
    .B2(net37),
    .X(_00253_));
 sky130_fd_sc_hd__xor2_1 _07157_ (.A(net91),
    .B(_00253_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_1 _07158_ (.A(_00239_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__a21bo_2 _07159_ (.A1(_00216_),
    .A2(_00238_),
    .B1_N(_00255_),
    .X(_00256_));
 sky130_fd_sc_hd__inv_2 _07160_ (.A(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__o31a_1 _07161_ (.A1(net291),
    .A2(net290),
    .A3(_00183_),
    .B1(net263),
    .X(_00258_));
 sky130_fd_sc_hd__o41a_2 _07162_ (.A1(net291),
    .A2(net290),
    .A3(reg1_val[16]),
    .A4(_00183_),
    .B1(net263),
    .X(_00259_));
 sky130_fd_sc_hd__xor2_2 _07163_ (.A(reg1_val[17]),
    .B(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__xnor2_2 _07164_ (.A(reg1_val[17]),
    .B(_00259_),
    .Y(_00261_));
 sky130_fd_sc_hd__o41a_2 _07165_ (.A1(reg1_val[11]),
    .A2(reg1_val[12]),
    .A3(reg1_val[13]),
    .A4(_00182_),
    .B1(net262),
    .X(_00262_));
 sky130_fd_sc_hd__o21a_1 _07166_ (.A1(reg1_val[14]),
    .A2(_00183_),
    .B1(net262),
    .X(_00263_));
 sky130_fd_sc_hd__xnor2_2 _07167_ (.A(net290),
    .B(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__xnor2_2 _07168_ (.A(reg1_val[16]),
    .B(_00258_),
    .Y(_00265_));
 sky130_fd_sc_hd__nor2_1 _07169_ (.A(net121),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_2 _07170_ (.A(net121),
    .B(_00265_),
    .Y(_00267_));
 sky130_fd_sc_hd__and2b_2 _07171_ (.A_N(_00266_),
    .B(_00267_),
    .X(_00268_));
 sky130_fd_sc_hd__nand2b_2 _07172_ (.A_N(_00266_),
    .B(_00267_),
    .Y(_00269_));
 sky130_fd_sc_hd__o41a_4 _07173_ (.A1(_06473_),
    .A2(_06474_),
    .A3(_06477_),
    .A4(_06478_),
    .B1(net175),
    .X(_00270_));
 sky130_fd_sc_hd__xnor2_2 _07174_ (.A(_06081_),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__xor2_4 _07175_ (.A(_06081_),
    .B(_00270_),
    .X(_00272_));
 sky130_fd_sc_hd__o31a_4 _07176_ (.A1(_06473_),
    .A2(_06474_),
    .A3(_06477_),
    .B1(net175),
    .X(_00273_));
 sky130_fd_sc_hd__o41a_4 _07177_ (.A1(_06148_),
    .A2(_06473_),
    .A3(_06474_),
    .A4(_06477_),
    .B1(net175),
    .X(_00274_));
 sky130_fd_sc_hd__xnor2_4 _07178_ (.A(_06118_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__xor2_4 _07179_ (.A(_06118_),
    .B(_00274_),
    .X(_00276_));
 sky130_fd_sc_hd__or3_4 _07180_ (.A(net125),
    .B(net121),
    .C(_00265_),
    .X(_00277_));
 sky130_fd_sc_hd__o21a_2 _07181_ (.A1(net124),
    .A2(_00267_),
    .B1(_00277_),
    .X(_00278_));
 sky130_fd_sc_hd__o21ai_4 _07182_ (.A1(net124),
    .A2(_00267_),
    .B1(_00277_),
    .Y(_00279_));
 sky130_fd_sc_hd__a22o_1 _07183_ (.A1(_00268_),
    .A2(net118),
    .B1(net115),
    .B2(_00279_),
    .X(_00280_));
 sky130_fd_sc_hd__xnor2_1 _07184_ (.A(net124),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__o41a_2 _07185_ (.A1(reg1_val[14]),
    .A2(reg1_val[15]),
    .A3(_00183_),
    .A4(_00185_),
    .B1(net263),
    .X(_00282_));
 sky130_fd_sc_hd__and3_1 _07186_ (.A(reg1_val[18]),
    .B(reg1_val[31]),
    .C(net295),
    .X(_00283_));
 sky130_fd_sc_hd__o21ai_2 _07187_ (.A1(_00282_),
    .A2(_00283_),
    .B1(reg1_val[19]),
    .Y(_00284_));
 sky130_fd_sc_hd__or3_2 _07188_ (.A(reg1_val[19]),
    .B(_00282_),
    .C(_00283_),
    .X(_00285_));
 sky130_fd_sc_hd__and2_4 _07189_ (.A(_00284_),
    .B(_00285_),
    .X(_00286_));
 sky130_fd_sc_hd__xor2_2 _07190_ (.A(reg1_val[20]),
    .B(_00187_),
    .X(_00287_));
 sky130_fd_sc_hd__a21oi_2 _07191_ (.A1(_00284_),
    .A2(_00285_),
    .B1(_00287_),
    .Y(_00288_));
 sky130_fd_sc_hd__and3_1 _07192_ (.A(_00284_),
    .B(_00285_),
    .C(_00287_),
    .X(_00289_));
 sky130_fd_sc_hd__nor2_2 _07193_ (.A(_00288_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__o21a_1 _07194_ (.A1(_06473_),
    .A2(_06474_),
    .B1(_06470_),
    .X(_00291_));
 sky130_fd_sc_hd__nand2_2 _07195_ (.A(_06241_),
    .B(_06470_),
    .Y(_00292_));
 sky130_fd_sc_hd__o22a_4 _07196_ (.A1(_06241_),
    .A2(_00291_),
    .B1(_00292_),
    .B2(_06475_),
    .X(_00293_));
 sky130_fd_sc_hd__o22ai_4 _07197_ (.A1(_06241_),
    .A2(_00291_),
    .B1(_00292_),
    .B2(_06475_),
    .Y(_00294_));
 sky130_fd_sc_hd__mux2_2 _07198_ (.A0(_00289_),
    .A1(_00288_),
    .S(_00201_),
    .X(_00295_));
 sky130_fd_sc_hd__a31o_4 _07199_ (.A1(_06309_),
    .A2(_06318_),
    .A3(_06472_),
    .B1(_06471_),
    .X(_00296_));
 sky130_fd_sc_hd__o41ai_4 _07200_ (.A1(_06302_),
    .A2(_06310_),
    .A3(net222),
    .A4(_06473_),
    .B1(net175),
    .Y(_00297_));
 sky130_fd_sc_hd__xor2_4 _07201_ (.A(_06285_),
    .B(_00297_),
    .X(_00298_));
 sky130_fd_sc_hd__xnor2_4 _07202_ (.A(_06285_),
    .B(net139),
    .Y(_00299_));
 sky130_fd_sc_hd__a22o_1 _07203_ (.A1(net30),
    .A2(_00293_),
    .B1(net28),
    .B2(net112),
    .X(_00300_));
 sky130_fd_sc_hd__xnor2_1 _07204_ (.A(net48),
    .B(_00300_),
    .Y(_00301_));
 sky130_fd_sc_hd__and2_1 _07205_ (.A(_00281_),
    .B(_00301_),
    .X(_00302_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_00281_),
    .B(_00301_),
    .Y(_00303_));
 sky130_fd_sc_hd__nor2_2 _07207_ (.A(_00302_),
    .B(_00303_),
    .Y(_00304_));
 sky130_fd_sc_hd__xnor2_2 _07208_ (.A(reg1_val[18]),
    .B(_00282_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_1 _07209_ (.A(_00261_),
    .B(_00305_),
    .Y(_00306_));
 sky130_fd_sc_hd__and2_1 _07210_ (.A(_00261_),
    .B(_00305_),
    .X(_00307_));
 sky130_fd_sc_hd__or2_2 _07211_ (.A(_00306_),
    .B(_00307_),
    .X(_00308_));
 sky130_fd_sc_hd__xor2_4 _07212_ (.A(_06148_),
    .B(_00273_),
    .X(_00309_));
 sky130_fd_sc_hd__xnor2_4 _07213_ (.A(_06148_),
    .B(_00273_),
    .Y(_00310_));
 sky130_fd_sc_hd__a211oi_2 _07214_ (.A1(_00284_),
    .A2(_00285_),
    .B1(_00305_),
    .C1(net124),
    .Y(_00311_));
 sky130_fd_sc_hd__a21oi_4 _07215_ (.A1(net88),
    .A2(_00307_),
    .B1(_00311_),
    .Y(_00312_));
 sky130_fd_sc_hd__o31a_4 _07216_ (.A1(_06241_),
    .A2(_06473_),
    .A3(_06474_),
    .B1(net175),
    .X(_00313_));
 sky130_fd_sc_hd__xnor2_4 _07217_ (.A(_06187_),
    .B(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__xnor2_4 _07218_ (.A(_06196_),
    .B(_00313_),
    .Y(_00315_));
 sky130_fd_sc_hd__o22a_2 _07219_ (.A1(net26),
    .A2(net111),
    .B1(net24),
    .B2(net108),
    .X(_00316_));
 sky130_fd_sc_hd__xnor2_4 _07220_ (.A(net87),
    .B(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__xnor2_4 _07221_ (.A(_00304_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__xor2_4 _07222_ (.A(_00256_),
    .B(_00318_),
    .X(_00319_));
 sky130_fd_sc_hd__a21o_1 _07223_ (.A1(_00137_),
    .A2(_00180_),
    .B1(_00319_),
    .X(_00320_));
 sky130_fd_sc_hd__xnor2_4 _07224_ (.A(_00181_),
    .B(_00319_),
    .Y(_00321_));
 sky130_fd_sc_hd__o31a_2 _07225_ (.A1(reg1_val[11]),
    .A2(reg1_val[12]),
    .A3(_00182_),
    .B1(net262),
    .X(_00322_));
 sky130_fd_sc_hd__xnor2_4 _07226_ (.A(reg1_val[13]),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__inv_6 _07227_ (.A(net138),
    .Y(_00324_));
 sky130_fd_sc_hd__a21oi_1 _07228_ (.A1(net262),
    .A2(_00182_),
    .B1(reg1_val[11]),
    .Y(_00325_));
 sky130_fd_sc_hd__and3_1 _07229_ (.A(reg1_val[11]),
    .B(net262),
    .C(_00182_),
    .X(_00326_));
 sky130_fd_sc_hd__or2_4 _07230_ (.A(_00325_),
    .B(_00326_),
    .X(_00327_));
 sky130_fd_sc_hd__inv_6 _07231_ (.A(net136),
    .Y(_00328_));
 sky130_fd_sc_hd__o21a_1 _07232_ (.A1(reg1_val[11]),
    .A2(_00182_),
    .B1(net262),
    .X(_00329_));
 sky130_fd_sc_hd__xnor2_2 _07233_ (.A(reg1_val[12]),
    .B(_00329_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(net135),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__or2_1 _07235_ (.A(net135),
    .B(_00330_),
    .X(_00332_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(_00331_),
    .B(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__a22oi_4 _07237_ (.A1(_05883_),
    .A2(_00170_),
    .B1(_00171_),
    .B2(_06481_),
    .Y(_00334_));
 sky130_fd_sc_hd__a22o_1 _07238_ (.A1(_05883_),
    .A2(_00170_),
    .B1(_00171_),
    .B2(_06481_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _07239_ (.A0(_00331_),
    .A1(_00332_),
    .S(net137),
    .X(_00336_));
 sky130_fd_sc_hd__o31a_2 _07240_ (.A1(_06476_),
    .A2(_06477_),
    .A3(_06479_),
    .B1(net175),
    .X(_00337_));
 sky130_fd_sc_hd__o41a_2 _07241_ (.A1(_05965_),
    .A2(_06476_),
    .A3(_06477_),
    .A4(_06479_),
    .B1(net175),
    .X(_00338_));
 sky130_fd_sc_hd__xnor2_2 _07242_ (.A(_05935_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__xor2_4 _07243_ (.A(_05935_),
    .B(_00338_),
    .X(_00340_));
 sky130_fd_sc_hd__o22a_1 _07244_ (.A1(net85),
    .A2(net83),
    .B1(net81),
    .B2(net79),
    .X(_00341_));
 sky130_fd_sc_hd__xnor2_1 _07245_ (.A(net137),
    .B(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__xnor2_4 _07246_ (.A(reg1_val[14]),
    .B(_00262_),
    .Y(_00343_));
 sky130_fd_sc_hd__or2_1 _07247_ (.A(net137),
    .B(_00343_),
    .X(_00344_));
 sky130_fd_sc_hd__nand2_1 _07248_ (.A(net137),
    .B(_00343_),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(_00344_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__xor2_4 _07250_ (.A(_05965_),
    .B(_00337_),
    .X(_00347_));
 sky130_fd_sc_hd__xnor2_2 _07251_ (.A(_05965_),
    .B(_00337_),
    .Y(_00348_));
 sky130_fd_sc_hd__mux2_1 _07252_ (.A0(_00345_),
    .A1(_00344_),
    .S(net122),
    .X(_00349_));
 sky130_fd_sc_hd__a21oi_4 _07253_ (.A1(_06081_),
    .A2(net175),
    .B1(_00270_),
    .Y(_00350_));
 sky130_fd_sc_hd__xor2_2 _07254_ (.A(_06026_),
    .B(_00350_),
    .X(_00351_));
 sky130_fd_sc_hd__xnor2_4 _07255_ (.A(_06026_),
    .B(_00350_),
    .Y(_00352_));
 sky130_fd_sc_hd__o22a_1 _07256_ (.A1(net77),
    .A2(net75),
    .B1(net73),
    .B2(net71),
    .X(_00353_));
 sky130_fd_sc_hd__xnor2_1 _07257_ (.A(net121),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__nor2_1 _07258_ (.A(_00342_),
    .B(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__and2_1 _07259_ (.A(_00342_),
    .B(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__nor2_1 _07260_ (.A(_00355_),
    .B(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__a22o_1 _07261_ (.A1(_00268_),
    .A2(net115),
    .B1(_00279_),
    .B2(_00309_),
    .X(_00358_));
 sky130_fd_sc_hd__xnor2_1 _07262_ (.A(net124),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__xnor2_4 _07263_ (.A(_06302_),
    .B(_00296_),
    .Y(_00360_));
 sky130_fd_sc_hd__xor2_4 _07264_ (.A(_06302_),
    .B(_00296_),
    .X(_00361_));
 sky130_fd_sc_hd__a22o_1 _07265_ (.A1(net30),
    .A2(net112),
    .B1(_00360_),
    .B2(net28),
    .X(_00362_));
 sky130_fd_sc_hd__xnor2_1 _07266_ (.A(net48),
    .B(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__and2_1 _07267_ (.A(_00359_),
    .B(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__xor2_1 _07268_ (.A(_00359_),
    .B(_00363_),
    .X(_00365_));
 sky130_fd_sc_hd__o22a_1 _07269_ (.A1(_00294_),
    .A2(net24),
    .B1(net109),
    .B2(net26),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_1 _07270_ (.A(net87),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__and2_1 _07271_ (.A(_00365_),
    .B(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__o21a_1 _07272_ (.A1(_00364_),
    .A2(_00368_),
    .B1(_00357_),
    .X(_00369_));
 sky130_fd_sc_hd__nor3_1 _07273_ (.A(_00357_),
    .B(_00364_),
    .C(_00368_),
    .Y(_00370_));
 sky130_fd_sc_hd__nor2_1 _07274_ (.A(_00369_),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__o31a_1 _07275_ (.A1(reg1_val[8]),
    .A2(reg1_val[9]),
    .A3(_00160_),
    .B1(net263),
    .X(_00372_));
 sky130_fd_sc_hd__xnor2_2 _07276_ (.A(reg1_val[10]),
    .B(_00372_),
    .Y(_00373_));
 sky130_fd_sc_hd__and2_1 _07277_ (.A(net173),
    .B(_00373_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _07278_ (.A(net173),
    .B(_00373_),
    .Y(_00375_));
 sky130_fd_sc_hd__nor2_1 _07279_ (.A(net173),
    .B(_00373_),
    .Y(_00376_));
 sky130_fd_sc_hd__or2_1 _07280_ (.A(net173),
    .B(_00373_),
    .X(_00377_));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(_00374_),
    .B(_00376_),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(_00375_),
    .B(_00377_),
    .Y(_00379_));
 sky130_fd_sc_hd__mux2_1 _07283_ (.A0(_00375_),
    .A1(_00377_),
    .S(net135),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _07284_ (.A0(_00374_),
    .A1(_00376_),
    .S(net135),
    .X(_00381_));
 sky130_fd_sc_hd__o22a_1 _07285_ (.A1(net98),
    .A2(net105),
    .B1(net103),
    .B2(net83),
    .X(_00382_));
 sky130_fd_sc_hd__xnor2_1 _07286_ (.A(net135),
    .B(_00382_),
    .Y(_00383_));
 sky130_fd_sc_hd__o22a_1 _07287_ (.A1(net119),
    .A2(net73),
    .B1(net71),
    .B2(net77),
    .X(_00384_));
 sky130_fd_sc_hd__xnor2_1 _07288_ (.A(net121),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__o22a_1 _07289_ (.A1(net85),
    .A2(net79),
    .B1(net75),
    .B2(net81),
    .X(_00386_));
 sky130_fd_sc_hd__xnor2_1 _07290_ (.A(net137),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__xnor2_1 _07291_ (.A(_00383_),
    .B(_00385_),
    .Y(_00388_));
 sky130_fd_sc_hd__nor2_1 _07292_ (.A(_00387_),
    .B(_00388_),
    .Y(_00389_));
 sky130_fd_sc_hd__o21bai_2 _07293_ (.A1(_00383_),
    .A2(_00385_),
    .B1_N(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__and2_1 _07294_ (.A(_00371_),
    .B(_00390_),
    .X(_00391_));
 sky130_fd_sc_hd__xnor2_1 _07295_ (.A(_00371_),
    .B(_00390_),
    .Y(_00392_));
 sky130_fd_sc_hd__o22a_1 _07296_ (.A1(net67),
    .A2(net151),
    .B1(net149),
    .B2(net64),
    .X(_00393_));
 sky130_fd_sc_hd__xnor2_2 _07297_ (.A(net193),
    .B(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__a21oi_4 _07298_ (.A1(net175),
    .A2(_06550_),
    .B1(_04899_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_4 _07299_ (.A(_04899_),
    .B(net175),
    .Y(_00396_));
 sky130_fd_sc_hd__nor2_8 _07300_ (.A(_06549_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__nor2_4 _07301_ (.A(_00395_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__or2_2 _07302_ (.A(_00395_),
    .B(_00397_),
    .X(_00399_));
 sky130_fd_sc_hd__o22a_1 _07303_ (.A1(net237),
    .A2(net55),
    .B1(net16),
    .B2(net288),
    .X(_00400_));
 sky130_fd_sc_hd__xnor2_2 _07304_ (.A(net239),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__o22a_1 _07305_ (.A1(net155),
    .A2(net58),
    .B1(net56),
    .B2(net153),
    .X(_00402_));
 sky130_fd_sc_hd__xnor2_2 _07306_ (.A(net194),
    .B(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__nor2_1 _07307_ (.A(_00401_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__xnor2_2 _07308_ (.A(_00401_),
    .B(_00403_),
    .Y(_00405_));
 sky130_fd_sc_hd__nor2_1 _07309_ (.A(_00394_),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__xnor2_2 _07310_ (.A(_00394_),
    .B(_00405_),
    .Y(_00407_));
 sky130_fd_sc_hd__o22a_1 _07311_ (.A1(net60),
    .A2(net147),
    .B1(net52),
    .B2(net145),
    .X(_00408_));
 sky130_fd_sc_hd__xnor2_1 _07312_ (.A(net189),
    .B(_00408_),
    .Y(_00409_));
 sky130_fd_sc_hd__o22a_1 _07313_ (.A1(net50),
    .A2(net134),
    .B1(net132),
    .B2(net100),
    .X(_00410_));
 sky130_fd_sc_hd__xnor2_1 _07314_ (.A(net172),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__nor2_2 _07315_ (.A(_00409_),
    .B(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__o22a_1 _07316_ (.A1(net100),
    .A2(net105),
    .B1(net103),
    .B2(net98),
    .X(_00413_));
 sky130_fd_sc_hd__xnor2_2 _07317_ (.A(net135),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__o22a_1 _07318_ (.A1(net62),
    .A2(net147),
    .B1(net145),
    .B2(net60),
    .X(_00415_));
 sky130_fd_sc_hd__xnor2_2 _07319_ (.A(net189),
    .B(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__nor2_1 _07320_ (.A(_00414_),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__xor2_2 _07321_ (.A(_00414_),
    .B(_00416_),
    .X(_00418_));
 sky130_fd_sc_hd__o22a_1 _07322_ (.A1(net52),
    .A2(net134),
    .B1(net132),
    .B2(net50),
    .X(_00419_));
 sky130_fd_sc_hd__xnor2_2 _07323_ (.A(net172),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__inv_2 _07324_ (.A(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__xnor2_2 _07325_ (.A(_00418_),
    .B(_00420_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _07326_ (.A(_00412_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__xnor2_2 _07327_ (.A(_00412_),
    .B(_00422_),
    .Y(_00424_));
 sky130_fd_sc_hd__xnor2_2 _07328_ (.A(_00407_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__a22o_1 _07329_ (.A1(_00225_),
    .A2(net41),
    .B1(_00250_),
    .B2(net43),
    .X(_00426_));
 sky130_fd_sc_hd__xor2_2 _07330_ (.A(net94),
    .B(_00426_),
    .X(_00427_));
 sky130_fd_sc_hd__o22a_1 _07331_ (.A1(net130),
    .A2(net45),
    .B1(net107),
    .B2(net47),
    .X(_00428_));
 sky130_fd_sc_hd__xnor2_1 _07332_ (.A(net97),
    .B(_00428_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(_00427_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__xor2_1 _07334_ (.A(_00427_),
    .B(_00429_),
    .X(_00431_));
 sky130_fd_sc_hd__a22o_1 _07335_ (.A1(_00211_),
    .A2(net39),
    .B1(net37),
    .B2(_00243_),
    .X(_00432_));
 sky130_fd_sc_hd__xor2_1 _07336_ (.A(net91),
    .B(_00432_),
    .X(_00433_));
 sky130_fd_sc_hd__nand2_1 _07337_ (.A(_00431_),
    .B(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__or2_1 _07338_ (.A(_00431_),
    .B(_00433_),
    .X(_00435_));
 sky130_fd_sc_hd__and2_1 _07339_ (.A(_00434_),
    .B(_00435_),
    .X(_00436_));
 sky130_fd_sc_hd__and2b_1 _07340_ (.A_N(_00425_),
    .B(_00436_),
    .X(_00437_));
 sky130_fd_sc_hd__xnor2_2 _07341_ (.A(_00425_),
    .B(_00436_),
    .Y(_00438_));
 sky130_fd_sc_hd__or3_4 _07342_ (.A(reg1_val[26]),
    .B(reg1_val[27]),
    .C(_00219_),
    .X(_00439_));
 sky130_fd_sc_hd__o21ai_2 _07343_ (.A1(_00218_),
    .A2(_00439_),
    .B1(net262),
    .Y(_00440_));
 sky130_fd_sc_hd__xnor2_4 _07344_ (.A(reg1_val[28]),
    .B(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__xor2_2 _07345_ (.A(net93),
    .B(_00441_),
    .X(_00442_));
 sky130_fd_sc_hd__xnor2_1 _07346_ (.A(net93),
    .B(_00441_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor2_1 _07347_ (.A(net210),
    .B(net23),
    .Y(_00444_));
 sky130_fd_sc_hd__or3b_2 _07348_ (.A(_06558_),
    .B(_06560_),
    .C_N(_00444_),
    .X(_00445_));
 sky130_fd_sc_hd__o21bai_1 _07349_ (.A1(_06558_),
    .A2(_06560_),
    .B1_N(_00444_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_2 _07350_ (.A(_00445_),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__xnor2_1 _07351_ (.A(_00438_),
    .B(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__nor2_1 _07352_ (.A(_00392_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _07353_ (.A(_00392_),
    .B(_00448_),
    .Y(_00450_));
 sky130_fd_sc_hd__and2b_1 _07354_ (.A_N(_00449_),
    .B(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__xor2_4 _07355_ (.A(_00321_),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__or2_1 _07356_ (.A(_00239_),
    .B(_00254_),
    .X(_00453_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_00255_),
    .B(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__nor2_1 _07358_ (.A(_00365_),
    .B(_00367_),
    .Y(_00455_));
 sky130_fd_sc_hd__or2_1 _07359_ (.A(_00368_),
    .B(_00455_),
    .X(_00456_));
 sky130_fd_sc_hd__xnor2_1 _07360_ (.A(_00178_),
    .B(_00179_),
    .Y(_00457_));
 sky130_fd_sc_hd__xnor2_1 _07361_ (.A(_00456_),
    .B(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__xnor2_1 _07362_ (.A(_00454_),
    .B(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__o22a_1 _07363_ (.A1(net83),
    .A2(net105),
    .B1(net103),
    .B2(net79),
    .X(_00460_));
 sky130_fd_sc_hd__xnor2_1 _07364_ (.A(net135),
    .B(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__o22a_1 _07365_ (.A1(net119),
    .A2(net77),
    .B1(net73),
    .B2(net117),
    .X(_00462_));
 sky130_fd_sc_hd__xnor2_1 _07366_ (.A(net121),
    .B(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__o22a_1 _07367_ (.A1(net85),
    .A2(net75),
    .B1(net71),
    .B2(net81),
    .X(_00464_));
 sky130_fd_sc_hd__xnor2_1 _07368_ (.A(net137),
    .B(_00464_),
    .Y(_00465_));
 sky130_fd_sc_hd__xnor2_1 _07369_ (.A(_00461_),
    .B(_00463_),
    .Y(_00466_));
 sky130_fd_sc_hd__nor2_1 _07370_ (.A(_00465_),
    .B(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__o21bai_2 _07371_ (.A1(_00461_),
    .A2(_00463_),
    .B1_N(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__and2_1 _07372_ (.A(_00409_),
    .B(_00411_),
    .X(_00469_));
 sky130_fd_sc_hd__nor2_1 _07373_ (.A(_00412_),
    .B(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__a22o_1 _07374_ (.A1(_00268_),
    .A2(_00309_),
    .B1(_00315_),
    .B2(_00279_),
    .X(_00471_));
 sky130_fd_sc_hd__xnor2_1 _07375_ (.A(net124),
    .B(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__a22o_1 _07376_ (.A1(_00198_),
    .A2(net28),
    .B1(_00360_),
    .B2(net30),
    .X(_00473_));
 sky130_fd_sc_hd__xnor2_1 _07377_ (.A(net48),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__and2_1 _07378_ (.A(_00472_),
    .B(_00474_),
    .X(_00475_));
 sky130_fd_sc_hd__nor2_1 _07379_ (.A(_00472_),
    .B(_00474_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_00475_),
    .B(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__o22a_1 _07381_ (.A1(_00294_),
    .A2(net26),
    .B1(net24),
    .B2(net113),
    .X(_00478_));
 sky130_fd_sc_hd__xnor2_1 _07382_ (.A(net87),
    .B(_00478_),
    .Y(_00479_));
 sky130_fd_sc_hd__and2_1 _07383_ (.A(_00477_),
    .B(_00479_),
    .X(_00480_));
 sky130_fd_sc_hd__o21a_1 _07384_ (.A1(_00475_),
    .A2(_00480_),
    .B1(_00470_),
    .X(_00481_));
 sky130_fd_sc_hd__nor3_1 _07385_ (.A(_00470_),
    .B(_00475_),
    .C(_00480_),
    .Y(_00482_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_00481_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__xnor2_1 _07387_ (.A(_00468_),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__nor2_1 _07388_ (.A(_00459_),
    .B(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__xor2_2 _07389_ (.A(_06542_),
    .B(_06543_),
    .X(_00486_));
 sky130_fd_sc_hd__and2_1 _07390_ (.A(net94),
    .B(_00486_),
    .X(_00487_));
 sky130_fd_sc_hd__o22a_1 _07391_ (.A1(net288),
    .A2(net64),
    .B1(net58),
    .B2(_06495_),
    .X(_00488_));
 sky130_fd_sc_hd__xnor2_2 _07392_ (.A(net239),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__o22a_1 _07393_ (.A1(net151),
    .A2(net56),
    .B1(net149),
    .B2(net62),
    .X(_00490_));
 sky130_fd_sc_hd__xnor2_2 _07394_ (.A(net193),
    .B(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__or2_1 _07395_ (.A(_00489_),
    .B(_00491_),
    .X(_00492_));
 sky130_fd_sc_hd__xnor2_2 _07396_ (.A(net94),
    .B(_00486_),
    .Y(_00493_));
 sky130_fd_sc_hd__nor2_1 _07397_ (.A(_00492_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__and2_1 _07398_ (.A(_00387_),
    .B(_00388_),
    .X(_00495_));
 sky130_fd_sc_hd__nor2_1 _07399_ (.A(_00389_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__o22a_1 _07400_ (.A1(net47),
    .A2(net128),
    .B1(net45),
    .B2(_00242_),
    .X(_00497_));
 sky130_fd_sc_hd__xor2_1 _07401_ (.A(net97),
    .B(_00497_),
    .X(_00498_));
 sky130_fd_sc_hd__nand2_1 _07402_ (.A(net208),
    .B(net43),
    .Y(_00499_));
 sky130_fd_sc_hd__xor2_1 _07403_ (.A(net94),
    .B(_00499_),
    .X(_00500_));
 sky130_fd_sc_hd__nor2_1 _07404_ (.A(_00498_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__and2_1 _07405_ (.A(_00498_),
    .B(_00500_),
    .X(_00502_));
 sky130_fd_sc_hd__or2_1 _07406_ (.A(_00501_),
    .B(_00502_),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _07407_ (.A1(net39),
    .A2(_00250_),
    .B1(net37),
    .B2(_00225_),
    .X(_00504_));
 sky130_fd_sc_hd__xor2_1 _07408_ (.A(net91),
    .B(_00504_),
    .X(_00505_));
 sky130_fd_sc_hd__and2b_1 _07409_ (.A_N(_00503_),
    .B(_00505_),
    .X(_00506_));
 sky130_fd_sc_hd__nor2_2 _07410_ (.A(_00501_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__xnor2_1 _07411_ (.A(_00496_),
    .B(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__o21ai_2 _07412_ (.A1(_00487_),
    .A2(_00494_),
    .B1(_00508_),
    .Y(_00509_));
 sky130_fd_sc_hd__or3_1 _07413_ (.A(_00487_),
    .B(_00494_),
    .C(_00508_),
    .X(_00510_));
 sky130_fd_sc_hd__and2_2 _07414_ (.A(_00509_),
    .B(_00510_),
    .X(_00511_));
 sky130_fd_sc_hd__nand2_1 _07415_ (.A(_00459_),
    .B(_00484_),
    .Y(_00512_));
 sky130_fd_sc_hd__and2b_1 _07416_ (.A_N(_00485_),
    .B(_00512_),
    .X(_00513_));
 sky130_fd_sc_hd__a21o_1 _07417_ (.A1(_00511_),
    .A2(_00512_),
    .B1(_00485_),
    .X(_00514_));
 sky130_fd_sc_hd__xnor2_2 _07418_ (.A(_00492_),
    .B(_00493_),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2_1 _07419_ (.A(_00477_),
    .B(_00479_),
    .Y(_00516_));
 sky130_fd_sc_hd__nor2_1 _07420_ (.A(_00480_),
    .B(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__and2b_1 _07421_ (.A_N(_00515_),
    .B(_00517_),
    .X(_00518_));
 sky130_fd_sc_hd__and2b_1 _07422_ (.A_N(_00505_),
    .B(_00503_),
    .X(_00519_));
 sky130_fd_sc_hd__or2_2 _07423_ (.A(_00506_),
    .B(_00519_),
    .X(_00520_));
 sky130_fd_sc_hd__inv_2 _07424_ (.A(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__xnor2_2 _07425_ (.A(_00515_),
    .B(_00517_),
    .Y(_00522_));
 sky130_fd_sc_hd__a21o_1 _07426_ (.A1(_00521_),
    .A2(_00522_),
    .B1(_00518_),
    .X(_00523_));
 sky130_fd_sc_hd__and2_1 _07427_ (.A(_00159_),
    .B(_00177_),
    .X(_00524_));
 sky130_fd_sc_hd__nor2_1 _07428_ (.A(_00178_),
    .B(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__o22a_1 _07429_ (.A1(net79),
    .A2(net105),
    .B1(net103),
    .B2(net75),
    .X(_00526_));
 sky130_fd_sc_hd__xnor2_1 _07430_ (.A(net135),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__o22a_1 _07431_ (.A1(net117),
    .A2(net77),
    .B1(net73),
    .B2(net111),
    .X(_00528_));
 sky130_fd_sc_hd__xnor2_1 _07432_ (.A(net121),
    .B(_00528_),
    .Y(_00529_));
 sky130_fd_sc_hd__nor2_1 _07433_ (.A(_00527_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__o22a_1 _07434_ (.A1(net119),
    .A2(net81),
    .B1(net71),
    .B2(net85),
    .X(_00531_));
 sky130_fd_sc_hd__xnor2_1 _07435_ (.A(net137),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__xnor2_1 _07436_ (.A(_00527_),
    .B(_00529_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _07437_ (.A(_00532_),
    .B(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__o21a_1 _07438_ (.A1(_00530_),
    .A2(_00534_),
    .B1(_00525_),
    .X(_00535_));
 sky130_fd_sc_hd__o22a_1 _07439_ (.A1(net134),
    .A2(net98),
    .B1(net132),
    .B2(net83),
    .X(_00536_));
 sky130_fd_sc_hd__xnor2_2 _07440_ (.A(net172),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__o22a_1 _07441_ (.A1(net155),
    .A2(net60),
    .B1(net52),
    .B2(net153),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_2 _07442_ (.A(net194),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__or2_1 _07443_ (.A(_00537_),
    .B(_00539_),
    .X(_00540_));
 sky130_fd_sc_hd__o22a_1 _07444_ (.A1(net147),
    .A2(net50),
    .B1(net100),
    .B2(net145),
    .X(_00541_));
 sky130_fd_sc_hd__xnor2_2 _07445_ (.A(net189),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__xnor2_2 _07446_ (.A(_00537_),
    .B(_00539_),
    .Y(_00543_));
 sky130_fd_sc_hd__o21ai_2 _07447_ (.A1(_00542_),
    .A2(_00543_),
    .B1(_00540_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor3_1 _07448_ (.A(_00525_),
    .B(_00530_),
    .C(_00534_),
    .Y(_00545_));
 sky130_fd_sc_hd__or2_1 _07449_ (.A(_00535_),
    .B(_00545_),
    .X(_00546_));
 sky130_fd_sc_hd__and2b_1 _07450_ (.A_N(_00546_),
    .B(_00544_),
    .X(_00547_));
 sky130_fd_sc_hd__nor2_1 _07451_ (.A(_00535_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__o21a_1 _07452_ (.A1(_00535_),
    .A2(_00547_),
    .B1(_00523_),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _07453_ (.A(_00465_),
    .B(_00466_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(_00467_),
    .B(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__a22o_1 _07455_ (.A1(_00279_),
    .A2(_00293_),
    .B1(_00315_),
    .B2(_00268_),
    .X(_00552_));
 sky130_fd_sc_hd__xnor2_1 _07456_ (.A(net124),
    .B(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__a22o_1 _07457_ (.A1(_00198_),
    .A2(net30),
    .B1(net28),
    .B2(_00211_),
    .X(_00554_));
 sky130_fd_sc_hd__xnor2_1 _07458_ (.A(net48),
    .B(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__and2_1 _07459_ (.A(_00553_),
    .B(_00555_),
    .X(_00556_));
 sky130_fd_sc_hd__xor2_1 _07460_ (.A(_00553_),
    .B(_00555_),
    .X(_00557_));
 sky130_fd_sc_hd__o22a_1 _07461_ (.A1(net113),
    .A2(net26),
    .B1(net24),
    .B2(_00361_),
    .X(_00558_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(net87),
    .B(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__and2_1 _07463_ (.A(_00557_),
    .B(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__o21a_1 _07464_ (.A1(_00556_),
    .A2(_00560_),
    .B1(_00551_),
    .X(_00561_));
 sky130_fd_sc_hd__o22a_1 _07465_ (.A1(net62),
    .A2(net151),
    .B1(net149),
    .B2(net60),
    .X(_00562_));
 sky130_fd_sc_hd__xor2_2 _07466_ (.A(net193),
    .B(_00562_),
    .X(_00563_));
 sky130_fd_sc_hd__o22a_2 _07467_ (.A1(net288),
    .A2(net58),
    .B1(net56),
    .B2(_06495_),
    .X(_00564_));
 sky130_fd_sc_hd__xnor2_4 _07468_ (.A(net240),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__o22a_1 _07469_ (.A1(net47),
    .A2(_00242_),
    .B1(_00249_),
    .B2(net45),
    .X(_00566_));
 sky130_fd_sc_hd__xnor2_1 _07470_ (.A(net97),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__and3_1 _07471_ (.A(_00563_),
    .B(_00565_),
    .C(_00567_),
    .X(_00568_));
 sky130_fd_sc_hd__a21oi_1 _07472_ (.A1(_00563_),
    .A2(_00565_),
    .B1(_00567_),
    .Y(_00569_));
 sky130_fd_sc_hd__a22o_1 _07473_ (.A1(_00225_),
    .A2(net39),
    .B1(net37),
    .B2(net208),
    .X(_00570_));
 sky130_fd_sc_hd__xor2_1 _07474_ (.A(net91),
    .B(_00570_),
    .X(_00571_));
 sky130_fd_sc_hd__or3b_1 _07475_ (.A(_00568_),
    .B(_00569_),
    .C_N(_00571_),
    .X(_00572_));
 sky130_fd_sc_hd__nand2b_1 _07476_ (.A_N(_00568_),
    .B(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__nor3_1 _07477_ (.A(_00551_),
    .B(_00556_),
    .C(_00560_),
    .Y(_00574_));
 sky130_fd_sc_hd__nor2_1 _07478_ (.A(_00561_),
    .B(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__a21o_1 _07479_ (.A1(_00573_),
    .A2(_00575_),
    .B1(_00561_),
    .X(_00576_));
 sky130_fd_sc_hd__xnor2_2 _07480_ (.A(_00523_),
    .B(_00548_),
    .Y(_00577_));
 sky130_fd_sc_hd__a21o_1 _07481_ (.A1(_00576_),
    .A2(_00577_),
    .B1(_00549_),
    .X(_00578_));
 sky130_fd_sc_hd__o31ai_4 _07482_ (.A1(_00389_),
    .A2(_00495_),
    .A3(_00507_),
    .B1(_00509_),
    .Y(_00579_));
 sky130_fd_sc_hd__o32a_2 _07483_ (.A1(_00368_),
    .A2(_00455_),
    .A3(_00457_),
    .B1(_00458_),
    .B2(_00454_),
    .X(_00580_));
 sky130_fd_sc_hd__a21oi_2 _07484_ (.A1(_00468_),
    .A2(_00483_),
    .B1(_00481_),
    .Y(_00581_));
 sky130_fd_sc_hd__nor2_1 _07485_ (.A(_00580_),
    .B(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__xor2_4 _07486_ (.A(_00580_),
    .B(_00581_),
    .X(_00583_));
 sky130_fd_sc_hd__xor2_2 _07487_ (.A(_00579_),
    .B(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__xnor2_2 _07488_ (.A(_00578_),
    .B(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2b_1 _07489_ (.A_N(_00585_),
    .B(_00514_),
    .Y(_00586_));
 sky130_fd_sc_hd__xnor2_2 _07490_ (.A(_00514_),
    .B(_00585_),
    .Y(_00587_));
 sky130_fd_sc_hd__and2_1 _07491_ (.A(_00452_),
    .B(_00587_),
    .X(_00588_));
 sky130_fd_sc_hd__xor2_2 _07492_ (.A(_00489_),
    .B(_00491_),
    .X(_00589_));
 sky130_fd_sc_hd__o22a_1 _07493_ (.A1(net75),
    .A2(net106),
    .B1(net104),
    .B2(net71),
    .X(_00590_));
 sky130_fd_sc_hd__xnor2_2 _07494_ (.A(net136),
    .B(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__o22a_1 _07495_ (.A1(net110),
    .A2(net78),
    .B1(net74),
    .B2(net109),
    .X(_00592_));
 sky130_fd_sc_hd__xnor2_2 _07496_ (.A(net121),
    .B(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__or2_1 _07497_ (.A(_00591_),
    .B(_00593_),
    .X(_00594_));
 sky130_fd_sc_hd__o22a_1 _07498_ (.A1(net119),
    .A2(net86),
    .B1(net82),
    .B2(net116),
    .X(_00595_));
 sky130_fd_sc_hd__xnor2_2 _07499_ (.A(net138),
    .B(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__xnor2_2 _07500_ (.A(_00591_),
    .B(_00593_),
    .Y(_00597_));
 sky130_fd_sc_hd__o21ai_1 _07501_ (.A1(_00596_),
    .A2(_00597_),
    .B1(_00594_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(_00589_),
    .B(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__xnor2_1 _07503_ (.A(_00589_),
    .B(_00598_),
    .Y(_00600_));
 sky130_fd_sc_hd__o22a_1 _07504_ (.A1(net155),
    .A2(net52),
    .B1(net50),
    .B2(net153),
    .X(_00601_));
 sky130_fd_sc_hd__xnor2_1 _07505_ (.A(net194),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__o22a_1 _07506_ (.A1(net133),
    .A2(net83),
    .B1(net79),
    .B2(net131),
    .X(_00603_));
 sky130_fd_sc_hd__xnor2_1 _07507_ (.A(net171),
    .B(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__or2_1 _07508_ (.A(_00602_),
    .B(_00604_),
    .X(_00605_));
 sky130_fd_sc_hd__o22a_1 _07509_ (.A1(_00145_),
    .A2(net100),
    .B1(net98),
    .B2(net145),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_1 _07510_ (.A(net189),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__xnor2_1 _07511_ (.A(_00602_),
    .B(_00604_),
    .Y(_00608_));
 sky130_fd_sc_hd__or2_1 _07512_ (.A(_00607_),
    .B(_00608_),
    .X(_00609_));
 sky130_fd_sc_hd__a21o_1 _07513_ (.A1(_00605_),
    .A2(_00609_),
    .B1(_00600_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_1 _07514_ (.A(_00599_),
    .B(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__and2_1 _07515_ (.A(_00532_),
    .B(_00533_),
    .X(_00612_));
 sky130_fd_sc_hd__nor2_1 _07516_ (.A(_00534_),
    .B(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__o21bai_1 _07517_ (.A1(_00568_),
    .A2(_00569_),
    .B1_N(_00571_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand3_1 _07518_ (.A(_00572_),
    .B(_00613_),
    .C(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__nor2_1 _07519_ (.A(_00557_),
    .B(_00559_),
    .Y(_00616_));
 sky130_fd_sc_hd__nor2_1 _07520_ (.A(_00560_),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__a21o_1 _07521_ (.A1(_00572_),
    .A2(_00614_),
    .B1(_00613_),
    .X(_00618_));
 sky130_fd_sc_hd__nand3_1 _07522_ (.A(_00615_),
    .B(_00617_),
    .C(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__a21boi_2 _07523_ (.A1(_00617_),
    .A2(_00618_),
    .B1_N(_00615_),
    .Y(_00620_));
 sky130_fd_sc_hd__a21o_1 _07524_ (.A1(_00599_),
    .A2(_00610_),
    .B1(_00620_),
    .X(_00621_));
 sky130_fd_sc_hd__xor2_1 _07525_ (.A(_00542_),
    .B(_00543_),
    .X(_00622_));
 sky130_fd_sc_hd__a22o_1 _07526_ (.A1(_00268_),
    .A2(_00293_),
    .B1(net112),
    .B2(_00279_),
    .X(_00623_));
 sky130_fd_sc_hd__xnor2_1 _07527_ (.A(net124),
    .B(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hd__a22o_1 _07528_ (.A1(_00211_),
    .A2(net30),
    .B1(net28),
    .B2(_00243_),
    .X(_00625_));
 sky130_fd_sc_hd__xnor2_1 _07529_ (.A(net48),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__and2_1 _07530_ (.A(_00624_),
    .B(_00626_),
    .X(_00627_));
 sky130_fd_sc_hd__xor2_1 _07531_ (.A(_00624_),
    .B(_00626_),
    .X(_00628_));
 sky130_fd_sc_hd__o22a_1 _07532_ (.A1(net129),
    .A2(net24),
    .B1(_00361_),
    .B2(net26),
    .X(_00629_));
 sky130_fd_sc_hd__xnor2_1 _07533_ (.A(net87),
    .B(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__and2_1 _07534_ (.A(_00628_),
    .B(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__o21a_1 _07535_ (.A1(_00627_),
    .A2(_00631_),
    .B1(_00622_),
    .X(_00632_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(net208),
    .B(net39),
    .Y(_00633_));
 sky130_fd_sc_hd__o22a_1 _07537_ (.A1(net45),
    .A2(net143),
    .B1(net140),
    .B2(net47),
    .X(_00634_));
 sky130_fd_sc_hd__xor2_1 _07538_ (.A(net97),
    .B(_00634_),
    .X(_00635_));
 sky130_fd_sc_hd__and3_1 _07539_ (.A(net208),
    .B(net39),
    .C(_00635_),
    .X(_00636_));
 sky130_fd_sc_hd__a21oi_1 _07540_ (.A1(net208),
    .A2(net39),
    .B1(net91),
    .Y(_00637_));
 sky130_fd_sc_hd__nor3_1 _07541_ (.A(_00622_),
    .B(_00627_),
    .C(_00631_),
    .Y(_00638_));
 sky130_fd_sc_hd__nor4_1 _07542_ (.A(_00632_),
    .B(_00636_),
    .C(_00637_),
    .D(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__or2_1 _07543_ (.A(_00632_),
    .B(_00639_),
    .X(_00640_));
 sky130_fd_sc_hd__xnor2_2 _07544_ (.A(_00611_),
    .B(_00620_),
    .Y(_00641_));
 sky130_fd_sc_hd__a21bo_1 _07545_ (.A1(_00640_),
    .A2(_00641_),
    .B1_N(_00621_),
    .X(_00642_));
 sky130_fd_sc_hd__xor2_2 _07546_ (.A(_00576_),
    .B(_00577_),
    .X(_00643_));
 sky130_fd_sc_hd__xnor2_2 _07547_ (.A(_00520_),
    .B(_00522_),
    .Y(_00644_));
 sky130_fd_sc_hd__xnor2_2 _07548_ (.A(_00544_),
    .B(_00546_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _07549_ (.A(_00644_),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__xnor2_2 _07550_ (.A(_00644_),
    .B(_00645_),
    .Y(_00647_));
 sky130_fd_sc_hd__xnor2_2 _07551_ (.A(_00573_),
    .B(_00575_),
    .Y(_00648_));
 sky130_fd_sc_hd__o21ai_2 _07552_ (.A1(_00647_),
    .A2(_00648_),
    .B1(_00646_),
    .Y(_00649_));
 sky130_fd_sc_hd__xnor2_2 _07553_ (.A(_00642_),
    .B(_00643_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2b_1 _07554_ (.A_N(_00650_),
    .B(_00649_),
    .Y(_00651_));
 sky130_fd_sc_hd__a21bo_2 _07555_ (.A1(_00642_),
    .A2(_00643_),
    .B1_N(_00651_),
    .X(_00652_));
 sky130_fd_sc_hd__xor2_4 _07556_ (.A(_00452_),
    .B(_00587_),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_4 _07557_ (.A1(_00652_),
    .A2(_00653_),
    .B1(_00588_),
    .Y(_00654_));
 sky130_fd_sc_hd__a21bo_2 _07558_ (.A1(_00578_),
    .A2(_00584_),
    .B1_N(_00586_),
    .X(_00655_));
 sky130_fd_sc_hd__o21a_2 _07559_ (.A1(_00407_),
    .A2(_00424_),
    .B1(_00423_),
    .X(_00656_));
 sky130_fd_sc_hd__o22a_1 _07560_ (.A1(net119),
    .A2(net32),
    .B1(net72),
    .B2(net34),
    .X(_00657_));
 sky130_fd_sc_hd__xnor2_1 _07561_ (.A(net125),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__a22o_1 _07562_ (.A1(_00293_),
    .A2(net28),
    .B1(_00315_),
    .B2(net30),
    .X(_00659_));
 sky130_fd_sc_hd__xnor2_1 _07563_ (.A(net48),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__and2_1 _07564_ (.A(_00658_),
    .B(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__nor2_1 _07565_ (.A(_00658_),
    .B(_00660_),
    .Y(_00662_));
 sky130_fd_sc_hd__nor2_1 _07566_ (.A(_00661_),
    .B(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__o22a_1 _07567_ (.A1(net117),
    .A2(net26),
    .B1(net111),
    .B2(net24),
    .X(_00664_));
 sky130_fd_sc_hd__xnor2_1 _07568_ (.A(net87),
    .B(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__xor2_1 _07569_ (.A(_00663_),
    .B(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__o31a_2 _07570_ (.A1(reg1_val[28]),
    .A2(_00218_),
    .A3(_00439_),
    .B1(net262),
    .X(_00667_));
 sky130_fd_sc_hd__xor2_4 _07571_ (.A(reg1_val[29]),
    .B(_00667_),
    .X(_00668_));
 sky130_fd_sc_hd__xnor2_1 _07572_ (.A(reg1_val[29]),
    .B(_00667_),
    .Y(_00669_));
 sky130_fd_sc_hd__or2_1 _07573_ (.A(_00444_),
    .B(_00668_),
    .X(_00670_));
 sky130_fd_sc_hd__and3_1 _07574_ (.A(_00445_),
    .B(_00666_),
    .C(_00670_),
    .X(_00671_));
 sky130_fd_sc_hd__a21oi_2 _07575_ (.A1(_00445_),
    .A2(_00670_),
    .B1(_00666_),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_2 _07576_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__xnor2_4 _07577_ (.A(_00656_),
    .B(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__a21o_1 _07578_ (.A1(_00418_),
    .A2(_00421_),
    .B1(_00417_),
    .X(_00675_));
 sky130_fd_sc_hd__a21o_1 _07579_ (.A1(net93),
    .A2(_00441_),
    .B1(_00668_),
    .X(_00676_));
 sky130_fd_sc_hd__o21ai_2 _07580_ (.A1(net93),
    .A2(_00441_),
    .B1(_00668_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(_00676_),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__o22a_1 _07582_ (.A1(net143),
    .A2(net23),
    .B1(net15),
    .B2(net210),
    .X(_00679_));
 sky130_fd_sc_hd__xnor2_1 _07583_ (.A(_00668_),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__xor2_1 _07584_ (.A(_00675_),
    .B(_00680_),
    .X(_00681_));
 sky130_fd_sc_hd__o21a_1 _07585_ (.A1(_00404_),
    .A2(_00406_),
    .B1(_00681_),
    .X(_00682_));
 sky130_fd_sc_hd__nor3_1 _07586_ (.A(_00404_),
    .B(_00406_),
    .C(_00681_),
    .Y(_00683_));
 sky130_fd_sc_hd__nor2_1 _07587_ (.A(_00682_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__o22a_1 _07588_ (.A1(net67),
    .A2(net149),
    .B1(net55),
    .B2(net151),
    .X(_00685_));
 sky130_fd_sc_hd__xnor2_2 _07589_ (.A(net192),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__a211o_4 _07590_ (.A1(_04888_),
    .A2(_06549_),
    .B1(net174),
    .C1(_04812_),
    .X(_00687_));
 sky130_fd_sc_hd__o211ai_4 _07591_ (.A1(net174),
    .A2(_06549_),
    .B1(_00396_),
    .C1(_04812_),
    .Y(_00688_));
 sky130_fd_sc_hd__and2_2 _07592_ (.A(_00687_),
    .B(_00688_),
    .X(_00689_));
 sky130_fd_sc_hd__nand2_4 _07593_ (.A(_00687_),
    .B(_00688_),
    .Y(_00690_));
 sky130_fd_sc_hd__a22o_1 _07594_ (.A1(_06494_),
    .A2(_00398_),
    .B1(_00690_),
    .B2(net292),
    .X(_00691_));
 sky130_fd_sc_hd__xnor2_2 _07595_ (.A(_06468_),
    .B(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__o22a_1 _07596_ (.A1(net64),
    .A2(net155),
    .B1(net153),
    .B2(net58),
    .X(_00693_));
 sky130_fd_sc_hd__xnor2_2 _07597_ (.A(net194),
    .B(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__or2_1 _07598_ (.A(_00692_),
    .B(_00694_),
    .X(_00695_));
 sky130_fd_sc_hd__xnor2_2 _07599_ (.A(_00692_),
    .B(_00694_),
    .Y(_00696_));
 sky130_fd_sc_hd__xnor2_2 _07600_ (.A(_00686_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__o22a_1 _07601_ (.A1(net50),
    .A2(net105),
    .B1(net103),
    .B2(net100),
    .X(_00698_));
 sky130_fd_sc_hd__xnor2_1 _07602_ (.A(net135),
    .B(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__o22a_1 _07603_ (.A1(net56),
    .A2(net147),
    .B1(net145),
    .B2(net62),
    .X(_00700_));
 sky130_fd_sc_hd__xnor2_1 _07604_ (.A(net189),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__xor2_1 _07605_ (.A(_00699_),
    .B(_00701_),
    .X(_00702_));
 sky130_fd_sc_hd__o22a_1 _07606_ (.A1(net60),
    .A2(net134),
    .B1(net132),
    .B2(net52),
    .X(_00703_));
 sky130_fd_sc_hd__xnor2_1 _07607_ (.A(net172),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__and2b_1 _07608_ (.A_N(_00704_),
    .B(_00702_),
    .X(_00705_));
 sky130_fd_sc_hd__xnor2_1 _07609_ (.A(_00702_),
    .B(_00704_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_00355_),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__xnor2_1 _07611_ (.A(_00355_),
    .B(_00706_),
    .Y(_00708_));
 sky130_fd_sc_hd__xnor2_1 _07612_ (.A(_00697_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__a22o_1 _07613_ (.A1(net43),
    .A2(_00243_),
    .B1(_00250_),
    .B2(net41),
    .X(_00710_));
 sky130_fd_sc_hd__xor2_1 _07614_ (.A(net94),
    .B(_00710_),
    .X(_00711_));
 sky130_fd_sc_hd__o22a_1 _07615_ (.A1(net47),
    .A2(_00298_),
    .B1(_00361_),
    .B2(net45),
    .X(_00712_));
 sky130_fd_sc_hd__xnor2_1 _07616_ (.A(net97),
    .B(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _07617_ (.A(_00711_),
    .B(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__or2_1 _07618_ (.A(_00711_),
    .B(_00713_),
    .X(_00715_));
 sky130_fd_sc_hd__and2_1 _07619_ (.A(_00714_),
    .B(_00715_),
    .X(_00716_));
 sky130_fd_sc_hd__a22o_1 _07620_ (.A1(_00198_),
    .A2(net39),
    .B1(net37),
    .B2(_00211_),
    .X(_00717_));
 sky130_fd_sc_hd__xor2_1 _07621_ (.A(net91),
    .B(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _07622_ (.A(_00716_),
    .B(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__or2_1 _07623_ (.A(_00716_),
    .B(_00718_),
    .X(_00720_));
 sky130_fd_sc_hd__and2_1 _07624_ (.A(_00719_),
    .B(_00720_),
    .X(_00721_));
 sky130_fd_sc_hd__and2b_1 _07625_ (.A_N(_00709_),
    .B(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__xnor2_1 _07626_ (.A(_00709_),
    .B(_00721_),
    .Y(_00723_));
 sky130_fd_sc_hd__xor2_1 _07627_ (.A(_00684_),
    .B(_00723_),
    .X(_00724_));
 sky130_fd_sc_hd__a21oi_2 _07628_ (.A1(_00304_),
    .A2(_00317_),
    .B1(_00302_),
    .Y(_00725_));
 sky130_fd_sc_hd__o22a_1 _07629_ (.A1(net98),
    .A2(net85),
    .B1(net83),
    .B2(net81),
    .X(_00726_));
 sky130_fd_sc_hd__xnor2_1 _07630_ (.A(net137),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__o22a_1 _07631_ (.A1(net79),
    .A2(net77),
    .B1(net75),
    .B2(net73),
    .X(_00728_));
 sky130_fd_sc_hd__xnor2_1 _07632_ (.A(net121),
    .B(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2_1 _07633_ (.A(_00727_),
    .B(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__and2_1 _07634_ (.A(_00727_),
    .B(_00729_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _07635_ (.A(_00730_),
    .B(_00731_),
    .X(_00732_));
 sky130_fd_sc_hd__a21oi_2 _07636_ (.A1(_00430_),
    .A2(_00434_),
    .B1(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__and3_1 _07637_ (.A(_00430_),
    .B(_00434_),
    .C(_00732_),
    .X(_00734_));
 sky130_fd_sc_hd__nor2_1 _07638_ (.A(_00733_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__and2b_1 _07639_ (.A_N(_00725_),
    .B(_00735_),
    .X(_00736_));
 sky130_fd_sc_hd__xnor2_1 _07640_ (.A(_00725_),
    .B(_00735_),
    .Y(_00737_));
 sky130_fd_sc_hd__and2_1 _07641_ (.A(_00724_),
    .B(_00737_),
    .X(_00738_));
 sky130_fd_sc_hd__nor2_1 _07642_ (.A(_00724_),
    .B(_00737_),
    .Y(_00739_));
 sky130_fd_sc_hd__nor2_2 _07643_ (.A(_00738_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__xor2_4 _07644_ (.A(_00674_),
    .B(_00740_),
    .X(_00741_));
 sky130_fd_sc_hd__a21o_1 _07645_ (.A1(_00321_),
    .A2(_00450_),
    .B1(_00449_),
    .X(_00742_));
 sky130_fd_sc_hd__o21ai_4 _07646_ (.A1(_00257_),
    .A2(_00318_),
    .B1(_00320_),
    .Y(_00743_));
 sky130_fd_sc_hd__or2_2 _07647_ (.A(_00369_),
    .B(_00391_),
    .X(_00744_));
 sky130_fd_sc_hd__a21oi_4 _07648_ (.A1(_00438_),
    .A2(_00447_),
    .B1(_00437_),
    .Y(_00745_));
 sky130_fd_sc_hd__o21ba_1 _07649_ (.A1(_00369_),
    .A2(_00391_),
    .B1_N(_00745_),
    .X(_00746_));
 sky130_fd_sc_hd__xnor2_4 _07650_ (.A(_00744_),
    .B(_00745_),
    .Y(_00747_));
 sky130_fd_sc_hd__xnor2_4 _07651_ (.A(_00743_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__a21oi_4 _07652_ (.A1(_00579_),
    .A2(_00583_),
    .B1(_00582_),
    .Y(_00749_));
 sky130_fd_sc_hd__xnor2_2 _07653_ (.A(_00748_),
    .B(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand2b_1 _07654_ (.A_N(_00750_),
    .B(_00742_),
    .Y(_00751_));
 sky130_fd_sc_hd__xnor2_2 _07655_ (.A(_00742_),
    .B(_00750_),
    .Y(_00752_));
 sky130_fd_sc_hd__and2_1 _07656_ (.A(_00741_),
    .B(_00752_),
    .X(_00753_));
 sky130_fd_sc_hd__xor2_4 _07657_ (.A(_00741_),
    .B(_00752_),
    .X(_00754_));
 sky130_fd_sc_hd__xnor2_4 _07658_ (.A(_00655_),
    .B(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__or2_1 _07659_ (.A(_00654_),
    .B(_00755_),
    .X(_00756_));
 sky130_fd_sc_hd__xnor2_2 _07660_ (.A(_00654_),
    .B(_00755_),
    .Y(_00757_));
 sky130_fd_sc_hd__xnor2_4 _07661_ (.A(_00652_),
    .B(_00653_),
    .Y(_00758_));
 sky130_fd_sc_hd__xor2_4 _07662_ (.A(_00511_),
    .B(_00513_),
    .X(_00759_));
 sky130_fd_sc_hd__xnor2_2 _07663_ (.A(_00649_),
    .B(_00650_),
    .Y(_00760_));
 sky130_fd_sc_hd__and2_1 _07664_ (.A(_00759_),
    .B(_00760_),
    .X(_00761_));
 sky130_fd_sc_hd__xnor2_2 _07665_ (.A(_00640_),
    .B(_00641_),
    .Y(_00762_));
 sky130_fd_sc_hd__xor2_2 _07666_ (.A(_00563_),
    .B(_00565_),
    .X(_00763_));
 sky130_fd_sc_hd__o22a_2 _07667_ (.A1(net71),
    .A2(net106),
    .B1(net104),
    .B2(net119),
    .X(_00764_));
 sky130_fd_sc_hd__xnor2_4 _07668_ (.A(net136),
    .B(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__o22a_2 _07669_ (.A1(net146),
    .A2(net98),
    .B1(net83),
    .B2(net144),
    .X(_00766_));
 sky130_fd_sc_hd__xnor2_4 _07670_ (.A(net188),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_1 _07671_ (.A(_00765_),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__xor2_4 _07672_ (.A(_00765_),
    .B(_00767_),
    .X(_00769_));
 sky130_fd_sc_hd__o22a_2 _07673_ (.A1(net133),
    .A2(net79),
    .B1(net75),
    .B2(net131),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_4 _07674_ (.A(net622),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_2 _07675_ (.A(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__a21oi_1 _07676_ (.A1(_00769_),
    .A2(_00772_),
    .B1(_00768_),
    .Y(_00773_));
 sky130_fd_sc_hd__and2b_1 _07677_ (.A_N(_00773_),
    .B(_00763_),
    .X(_00774_));
 sky130_fd_sc_hd__o22a_1 _07678_ (.A1(_06495_),
    .A2(net62),
    .B1(net56),
    .B2(net288),
    .X(_00775_));
 sky130_fd_sc_hd__xnor2_2 _07679_ (.A(net238),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__o22a_1 _07680_ (.A1(net155),
    .A2(net50),
    .B1(net100),
    .B2(net153),
    .X(_00777_));
 sky130_fd_sc_hd__xnor2_2 _07681_ (.A(net194),
    .B(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__or2_1 _07682_ (.A(_00776_),
    .B(_00778_),
    .X(_00779_));
 sky130_fd_sc_hd__o22a_1 _07683_ (.A1(net60),
    .A2(net150),
    .B1(net148),
    .B2(net52),
    .X(_00780_));
 sky130_fd_sc_hd__xnor2_2 _07684_ (.A(net191),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__xnor2_2 _07685_ (.A(_00776_),
    .B(_00778_),
    .Y(_00782_));
 sky130_fd_sc_hd__o21ai_1 _07686_ (.A1(_00781_),
    .A2(_00782_),
    .B1(_00779_),
    .Y(_00783_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(_00763_),
    .B(_00773_),
    .Y(_00784_));
 sky130_fd_sc_hd__a21o_1 _07688_ (.A1(_00783_),
    .A2(_00784_),
    .B1(_00774_),
    .X(_00785_));
 sky130_fd_sc_hd__xnor2_2 _07689_ (.A(_00596_),
    .B(_00597_),
    .Y(_00786_));
 sky130_fd_sc_hd__xnor2_1 _07690_ (.A(_00633_),
    .B(_00635_),
    .Y(_00787_));
 sky130_fd_sc_hd__nor2_1 _07691_ (.A(_00786_),
    .B(_00787_),
    .Y(_00788_));
 sky130_fd_sc_hd__xor2_1 _07692_ (.A(_00628_),
    .B(_00630_),
    .X(_00789_));
 sky130_fd_sc_hd__xor2_1 _07693_ (.A(_00786_),
    .B(_00787_),
    .X(_00790_));
 sky130_fd_sc_hd__a21o_1 _07694_ (.A1(_00789_),
    .A2(_00790_),
    .B1(_00788_),
    .X(_00791_));
 sky130_fd_sc_hd__nand2_1 _07695_ (.A(_00785_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__o22a_2 _07696_ (.A1(net116),
    .A2(net86),
    .B1(net82),
    .B2(net110),
    .X(_00793_));
 sky130_fd_sc_hd__xnor2_4 _07697_ (.A(net138),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__a22o_1 _07698_ (.A1(_00268_),
    .A2(net112),
    .B1(_00360_),
    .B2(_00279_),
    .X(_00795_));
 sky130_fd_sc_hd__xnor2_2 _07699_ (.A(net125),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__or2_1 _07700_ (.A(_00794_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__xnor2_4 _07701_ (.A(_00794_),
    .B(_00796_),
    .Y(_00798_));
 sky130_fd_sc_hd__o22a_2 _07702_ (.A1(net108),
    .A2(net78),
    .B1(net74),
    .B2(net114),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_4 _07703_ (.A(net123),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__o21ai_1 _07704_ (.A1(_00798_),
    .A2(_00800_),
    .B1(_00797_),
    .Y(_00801_));
 sky130_fd_sc_hd__xor2_1 _07705_ (.A(_00607_),
    .B(_00608_),
    .X(_00802_));
 sky130_fd_sc_hd__and2_1 _07706_ (.A(_00801_),
    .B(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__o22a_2 _07707_ (.A1(net130),
    .A2(net26),
    .B1(net24),
    .B2(net128),
    .X(_00804_));
 sky130_fd_sc_hd__xnor2_4 _07708_ (.A(net87),
    .B(_00804_),
    .Y(_00805_));
 sky130_fd_sc_hd__a22o_1 _07709_ (.A1(_00243_),
    .A2(net30),
    .B1(net28),
    .B2(_00250_),
    .X(_00806_));
 sky130_fd_sc_hd__xnor2_4 _07710_ (.A(net48),
    .B(_00806_),
    .Y(_00807_));
 sky130_fd_sc_hd__and2_1 _07711_ (.A(_00805_),
    .B(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__xor2_1 _07712_ (.A(_00801_),
    .B(_00802_),
    .X(_00809_));
 sky130_fd_sc_hd__a21oi_1 _07713_ (.A1(_00808_),
    .A2(_00809_),
    .B1(_00803_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor2_1 _07714_ (.A(_00785_),
    .B(_00791_),
    .Y(_00811_));
 sky130_fd_sc_hd__xor2_1 _07715_ (.A(_00785_),
    .B(_00791_),
    .X(_00812_));
 sky130_fd_sc_hd__o21a_1 _07716_ (.A1(_00810_),
    .A2(_00811_),
    .B1(_00792_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _07717_ (.A(_00762_),
    .B(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__nand3_1 _07718_ (.A(_00600_),
    .B(_00605_),
    .C(_00609_),
    .Y(_00815_));
 sky130_fd_sc_hd__and2_1 _07719_ (.A(_00610_),
    .B(_00815_),
    .X(_00816_));
 sky130_fd_sc_hd__a21o_1 _07720_ (.A1(_00615_),
    .A2(_00618_),
    .B1(_00617_),
    .X(_00817_));
 sky130_fd_sc_hd__and3_1 _07721_ (.A(_00619_),
    .B(_00816_),
    .C(_00817_),
    .X(_00818_));
 sky130_fd_sc_hd__a21oi_1 _07722_ (.A1(_00619_),
    .A2(_00817_),
    .B1(_00816_),
    .Y(_00819_));
 sky130_fd_sc_hd__nor2_1 _07723_ (.A(_00818_),
    .B(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__o22a_1 _07724_ (.A1(_00636_),
    .A2(_00637_),
    .B1(_00638_),
    .B2(_00632_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _07725_ (.A(_00639_),
    .B(_00821_),
    .X(_00822_));
 sky130_fd_sc_hd__o21ba_1 _07726_ (.A1(_00819_),
    .A2(_00822_),
    .B1_N(_00818_),
    .X(_00823_));
 sky130_fd_sc_hd__xnor2_2 _07727_ (.A(_00762_),
    .B(_00813_),
    .Y(_00824_));
 sky130_fd_sc_hd__o21ai_4 _07728_ (.A1(_00823_),
    .A2(_00824_),
    .B1(_00814_),
    .Y(_00825_));
 sky130_fd_sc_hd__xor2_4 _07729_ (.A(_00759_),
    .B(_00760_),
    .X(_00826_));
 sky130_fd_sc_hd__a21oi_4 _07730_ (.A1(_00825_),
    .A2(_00826_),
    .B1(_00761_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_00758_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__xor2_2 _07732_ (.A(_00647_),
    .B(_00648_),
    .X(_00829_));
 sky130_fd_sc_hd__xor2_1 _07733_ (.A(_00823_),
    .B(_00824_),
    .X(_00830_));
 sky130_fd_sc_hd__xnor2_1 _07734_ (.A(_00810_),
    .B(_00812_),
    .Y(_00831_));
 sky130_fd_sc_hd__xor2_4 _07735_ (.A(_00805_),
    .B(_00807_),
    .X(_00832_));
 sky130_fd_sc_hd__xnor2_4 _07736_ (.A(_00769_),
    .B(_00771_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_00832_),
    .B(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__xnor2_4 _07738_ (.A(_00832_),
    .B(_00833_),
    .Y(_00835_));
 sky130_fd_sc_hd__xnor2_4 _07739_ (.A(_00798_),
    .B(_00800_),
    .Y(_00836_));
 sky130_fd_sc_hd__or2_1 _07740_ (.A(_00835_),
    .B(_00836_),
    .X(_00837_));
 sky130_fd_sc_hd__o21ai_4 _07741_ (.A1(_00835_),
    .A2(_00836_),
    .B1(_00834_),
    .Y(_00838_));
 sky130_fd_sc_hd__o22a_2 _07742_ (.A1(net146),
    .A2(net83),
    .B1(net79),
    .B2(net144),
    .X(_00839_));
 sky130_fd_sc_hd__xnor2_4 _07743_ (.A(net188),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__o22a_2 _07744_ (.A1(net119),
    .A2(net106),
    .B1(net104),
    .B2(net116),
    .X(_00841_));
 sky130_fd_sc_hd__xnor2_4 _07745_ (.A(net136),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _07746_ (.A(_00840_),
    .B(_00842_),
    .Y(_00843_));
 sky130_fd_sc_hd__xor2_4 _07747_ (.A(_00840_),
    .B(_00842_),
    .X(_00844_));
 sky130_fd_sc_hd__o22a_1 _07748_ (.A1(net133),
    .A2(net75),
    .B1(net71),
    .B2(net131),
    .X(_00845_));
 sky130_fd_sc_hd__xnor2_2 _07749_ (.A(net622),
    .B(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _07750_ (.A(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__a21oi_4 _07751_ (.A1(_00844_),
    .A2(_00847_),
    .B1(_00843_),
    .Y(_00848_));
 sky130_fd_sc_hd__o22a_2 _07752_ (.A1(net210),
    .A2(net45),
    .B1(net143),
    .B2(net47),
    .X(_00849_));
 sky130_fd_sc_hd__xnor2_4 _07753_ (.A(net97),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__and2b_1 _07754_ (.A_N(_00848_),
    .B(_00850_),
    .X(_00851_));
 sky130_fd_sc_hd__o22a_1 _07755_ (.A1(net287),
    .A2(net62),
    .B1(net60),
    .B2(net237),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_2 _07756_ (.A(net238),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__o22a_1 _07757_ (.A1(net154),
    .A2(net100),
    .B1(net98),
    .B2(net152),
    .X(_00854_));
 sky130_fd_sc_hd__xnor2_2 _07758_ (.A(net195),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__nor2_1 _07759_ (.A(_00853_),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_00853_),
    .B(_00855_),
    .Y(_00857_));
 sky130_fd_sc_hd__xnor2_1 _07761_ (.A(_00853_),
    .B(_00855_),
    .Y(_00858_));
 sky130_fd_sc_hd__o22a_1 _07762_ (.A1(net150),
    .A2(net52),
    .B1(net50),
    .B2(net148),
    .X(_00859_));
 sky130_fd_sc_hd__xor2_1 _07763_ (.A(net191),
    .B(_00859_),
    .X(_00860_));
 sky130_fd_sc_hd__a21o_2 _07764_ (.A1(_00857_),
    .A2(_00860_),
    .B1(_00856_),
    .X(_00861_));
 sky130_fd_sc_hd__xnor2_4 _07765_ (.A(_00848_),
    .B(_00850_),
    .Y(_00862_));
 sky130_fd_sc_hd__a21oi_4 _07766_ (.A1(_00861_),
    .A2(_00862_),
    .B1(_00851_),
    .Y(_00863_));
 sky130_fd_sc_hd__a21o_1 _07767_ (.A1(_00834_),
    .A2(_00837_),
    .B1(_00863_),
    .X(_00864_));
 sky130_fd_sc_hd__xor2_2 _07768_ (.A(_00781_),
    .B(_00782_),
    .X(_00865_));
 sky130_fd_sc_hd__o22a_1 _07769_ (.A1(net110),
    .A2(net86),
    .B1(net82),
    .B2(net108),
    .X(_00866_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(net138),
    .B(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__o22a_1 _07771_ (.A1(net129),
    .A2(net32),
    .B1(net107),
    .B2(net34),
    .X(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07772_ (.A(net124),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__nor2_1 _07773_ (.A(_00867_),
    .B(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(_00867_),
    .B(_00869_),
    .Y(_00871_));
 sky130_fd_sc_hd__o22a_1 _07775_ (.A1(net114),
    .A2(net78),
    .B1(net74),
    .B2(net113),
    .X(_00872_));
 sky130_fd_sc_hd__xnor2_1 _07776_ (.A(net123),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__o21ba_1 _07777_ (.A1(_00871_),
    .A2(_00873_),
    .B1_N(_00870_),
    .X(_00874_));
 sky130_fd_sc_hd__and2b_1 _07778_ (.A_N(_00874_),
    .B(_00865_),
    .X(_00875_));
 sky130_fd_sc_hd__o22a_1 _07779_ (.A1(net127),
    .A2(net26),
    .B1(net24),
    .B2(net141),
    .X(_00876_));
 sky130_fd_sc_hd__xnor2_2 _07780_ (.A(net87),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__a22o_1 _07781_ (.A1(_00250_),
    .A2(net30),
    .B1(net28),
    .B2(_00225_),
    .X(_00878_));
 sky130_fd_sc_hd__xnor2_2 _07782_ (.A(net48),
    .B(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__and2_1 _07783_ (.A(_00877_),
    .B(_00879_),
    .X(_00880_));
 sky130_fd_sc_hd__xnor2_1 _07784_ (.A(_00865_),
    .B(_00874_),
    .Y(_00881_));
 sky130_fd_sc_hd__a21o_2 _07785_ (.A1(_00880_),
    .A2(_00881_),
    .B1(_00875_),
    .X(_00882_));
 sky130_fd_sc_hd__xnor2_4 _07786_ (.A(_00838_),
    .B(_00863_),
    .Y(_00883_));
 sky130_fd_sc_hd__a21bo_1 _07787_ (.A1(_00882_),
    .A2(_00883_),
    .B1_N(_00864_),
    .X(_00884_));
 sky130_fd_sc_hd__xnor2_1 _07788_ (.A(_00783_),
    .B(_00784_),
    .Y(_00885_));
 sky130_fd_sc_hd__xnor2_1 _07789_ (.A(_00789_),
    .B(_00790_),
    .Y(_00886_));
 sky130_fd_sc_hd__xnor2_1 _07790_ (.A(_00808_),
    .B(_00809_),
    .Y(_00887_));
 sky130_fd_sc_hd__xnor2_1 _07791_ (.A(_00885_),
    .B(_00886_),
    .Y(_00888_));
 sky130_fd_sc_hd__nor2_1 _07792_ (.A(_00887_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21ba_1 _07793_ (.A1(_00885_),
    .A2(_00886_),
    .B1_N(_00889_),
    .X(_00890_));
 sky130_fd_sc_hd__xor2_1 _07794_ (.A(_00831_),
    .B(_00884_),
    .X(_00891_));
 sky130_fd_sc_hd__nand2b_1 _07795_ (.A_N(_00890_),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__a21bo_1 _07796_ (.A1(_00831_),
    .A2(_00884_),
    .B1_N(_00892_),
    .X(_00893_));
 sky130_fd_sc_hd__xnor2_1 _07797_ (.A(_00829_),
    .B(_00830_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2b_1 _07798_ (.A_N(_00894_),
    .B(_00893_),
    .Y(_00895_));
 sky130_fd_sc_hd__a21bo_2 _07799_ (.A1(_00829_),
    .A2(_00830_),
    .B1_N(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__xor2_4 _07800_ (.A(_00825_),
    .B(_00826_),
    .X(_00897_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(_00896_),
    .B(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__a2bb2o_1 _07802_ (.A1_N(_00758_),
    .A2_N(_00827_),
    .B1(_00896_),
    .B2(_00897_),
    .X(_00899_));
 sky130_fd_sc_hd__xnor2_1 _07803_ (.A(_00820_),
    .B(_00822_),
    .Y(_00900_));
 sky130_fd_sc_hd__xnor2_1 _07804_ (.A(_00890_),
    .B(_00891_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(_00900_),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__xnor2_4 _07806_ (.A(_00882_),
    .B(_00883_),
    .Y(_00903_));
 sky130_fd_sc_hd__xor2_2 _07807_ (.A(_00877_),
    .B(_00879_),
    .X(_00904_));
 sky130_fd_sc_hd__xnor2_2 _07808_ (.A(_00844_),
    .B(_00846_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _07809_ (.A(_00904_),
    .B(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__xnor2_1 _07810_ (.A(_00871_),
    .B(_00873_),
    .Y(_00907_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(_00904_),
    .B(_00905_),
    .Y(_00908_));
 sky130_fd_sc_hd__xor2_1 _07812_ (.A(_00904_),
    .B(_00905_),
    .X(_00909_));
 sky130_fd_sc_hd__o21a_1 _07813_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00906_),
    .X(_00910_));
 sky130_fd_sc_hd__nor2_1 _07814_ (.A(net210),
    .B(net47),
    .Y(_00911_));
 sky130_fd_sc_hd__a21oi_1 _07815_ (.A1(_06519_),
    .A2(_06520_),
    .B1(net288),
    .Y(_00912_));
 sky130_fd_sc_hd__and3_1 _07816_ (.A(_06494_),
    .B(_00146_),
    .C(_00147_),
    .X(_00913_));
 sky130_fd_sc_hd__o21a_1 _07817_ (.A1(_00912_),
    .A2(_00913_),
    .B1(net240),
    .X(_00914_));
 sky130_fd_sc_hd__nor3_1 _07818_ (.A(net240),
    .B(_00912_),
    .C(_00913_),
    .Y(_00915_));
 sky130_fd_sc_hd__o22a_1 _07819_ (.A1(net155),
    .A2(net98),
    .B1(net83),
    .B2(net153),
    .X(_00916_));
 sky130_fd_sc_hd__xnor2_1 _07820_ (.A(net194),
    .B(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__or3_2 _07821_ (.A(_00914_),
    .B(_00915_),
    .C(_00917_),
    .X(_00918_));
 sky130_fd_sc_hd__o21ai_1 _07822_ (.A1(_00914_),
    .A2(_00915_),
    .B1(_00917_),
    .Y(_00919_));
 sky130_fd_sc_hd__o22a_1 _07823_ (.A1(net151),
    .A2(net50),
    .B1(net100),
    .B2(net149),
    .X(_00920_));
 sky130_fd_sc_hd__xor2_1 _07824_ (.A(net192),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_00918_),
    .B(_00919_),
    .C(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_00918_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__mux2_1 _07827_ (.A0(net97),
    .A1(_00923_),
    .S(_00911_),
    .X(_00924_));
 sky130_fd_sc_hd__nand2b_1 _07828_ (.A_N(_00910_),
    .B(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(_00858_),
    .B(_00860_),
    .Y(_00926_));
 sky130_fd_sc_hd__o22a_1 _07830_ (.A1(net116),
    .A2(net106),
    .B1(net104),
    .B2(net110),
    .X(_00927_));
 sky130_fd_sc_hd__xnor2_1 _07831_ (.A(net136),
    .B(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__o22a_1 _07832_ (.A1(net146),
    .A2(net79),
    .B1(net75),
    .B2(net144),
    .X(_00929_));
 sky130_fd_sc_hd__xnor2_1 _07833_ (.A(net188),
    .B(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__xor2_1 _07834_ (.A(_00928_),
    .B(_00930_),
    .X(_00931_));
 sky130_fd_sc_hd__o22a_1 _07835_ (.A1(net131),
    .A2(net119),
    .B1(net71),
    .B2(net133),
    .X(_00932_));
 sky130_fd_sc_hd__xnor2_1 _07836_ (.A(net171),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__and2b_1 _07837_ (.A_N(_00933_),
    .B(_00931_),
    .X(_00934_));
 sky130_fd_sc_hd__o21ba_1 _07838_ (.A1(_00928_),
    .A2(_00930_),
    .B1_N(_00934_),
    .X(_00935_));
 sky130_fd_sc_hd__and2b_1 _07839_ (.A_N(_00935_),
    .B(_00926_),
    .X(_00936_));
 sky130_fd_sc_hd__o22a_1 _07840_ (.A1(net108),
    .A2(net86),
    .B1(net82),
    .B2(net114),
    .X(_00937_));
 sky130_fd_sc_hd__xnor2_1 _07841_ (.A(net138),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__o22a_1 _07842_ (.A1(net113),
    .A2(net78),
    .B1(net74),
    .B2(net107),
    .X(_00939_));
 sky130_fd_sc_hd__xnor2_1 _07843_ (.A(net123),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nor2_1 _07844_ (.A(_00938_),
    .B(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__xnor2_1 _07845_ (.A(_00926_),
    .B(_00935_),
    .Y(_00942_));
 sky130_fd_sc_hd__a21o_1 _07846_ (.A1(_00941_),
    .A2(_00942_),
    .B1(_00936_),
    .X(_00943_));
 sky130_fd_sc_hd__xnor2_2 _07847_ (.A(_00910_),
    .B(_00924_),
    .Y(_00944_));
 sky130_fd_sc_hd__a21bo_1 _07848_ (.A1(_00943_),
    .A2(_00944_),
    .B1_N(_00925_),
    .X(_00945_));
 sky130_fd_sc_hd__and2b_1 _07849_ (.A_N(_00903_),
    .B(_00945_),
    .X(_00946_));
 sky130_fd_sc_hd__xor2_2 _07850_ (.A(_00835_),
    .B(_00836_),
    .X(_00947_));
 sky130_fd_sc_hd__xor2_2 _07851_ (.A(_00861_),
    .B(_00862_),
    .X(_00948_));
 sky130_fd_sc_hd__xnor2_1 _07852_ (.A(_00947_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__xnor2_1 _07853_ (.A(_00880_),
    .B(_00881_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_1 _07854_ (.A(_00949_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__a21oi_4 _07855_ (.A1(_00947_),
    .A2(_00948_),
    .B1(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__xnor2_4 _07856_ (.A(_00903_),
    .B(_00945_),
    .Y(_00953_));
 sky130_fd_sc_hd__and2b_1 _07857_ (.A_N(_00952_),
    .B(_00953_),
    .X(_00954_));
 sky130_fd_sc_hd__xor2_1 _07858_ (.A(_00900_),
    .B(_00901_),
    .X(_00955_));
 sky130_fd_sc_hd__o21ai_1 _07859_ (.A1(_00946_),
    .A2(_00954_),
    .B1(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__xor2_1 _07860_ (.A(_00893_),
    .B(_00894_),
    .X(_00957_));
 sky130_fd_sc_hd__and3_1 _07861_ (.A(_00902_),
    .B(_00956_),
    .C(_00957_),
    .X(_00958_));
 sky130_fd_sc_hd__and2_1 _07862_ (.A(_00887_),
    .B(_00888_),
    .X(_00959_));
 sky130_fd_sc_hd__nor2_2 _07863_ (.A(_00889_),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__xnor2_4 _07864_ (.A(_00952_),
    .B(_00953_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_1 _07865_ (.A(_00960_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__a21o_1 _07866_ (.A1(_00918_),
    .A2(_00919_),
    .B1(_00921_),
    .X(_00963_));
 sky130_fd_sc_hd__and2_1 _07867_ (.A(_00938_),
    .B(_00940_),
    .X(_00964_));
 sky130_fd_sc_hd__nor2_1 _07868_ (.A(_00941_),
    .B(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__and3_1 _07869_ (.A(_00922_),
    .B(_00963_),
    .C(_00965_),
    .X(_00966_));
 sky130_fd_sc_hd__a21oi_1 _07870_ (.A1(_00922_),
    .A2(_00963_),
    .B1(_00965_),
    .Y(_00967_));
 sky130_fd_sc_hd__and2b_1 _07871_ (.A_N(_00931_),
    .B(_00933_),
    .X(_00968_));
 sky130_fd_sc_hd__or2_1 _07872_ (.A(_00934_),
    .B(_00968_),
    .X(_00969_));
 sky130_fd_sc_hd__or3_1 _07873_ (.A(_00966_),
    .B(_00967_),
    .C(_00969_),
    .X(_00970_));
 sky130_fd_sc_hd__o21ba_1 _07874_ (.A1(_00967_),
    .A2(_00969_),
    .B1_N(_00966_),
    .X(_00971_));
 sky130_fd_sc_hd__o22a_1 _07875_ (.A1(net130),
    .A2(net34),
    .B1(net32),
    .B2(net128),
    .X(_00972_));
 sky130_fd_sc_hd__xnor2_1 _07876_ (.A(net125),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__a22o_1 _07877_ (.A1(_00225_),
    .A2(net30),
    .B1(net28),
    .B2(net208),
    .X(_00974_));
 sky130_fd_sc_hd__xnor2_1 _07878_ (.A(net48),
    .B(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__and2_1 _07879_ (.A(_00973_),
    .B(_00975_),
    .X(_00976_));
 sky130_fd_sc_hd__nor2_1 _07880_ (.A(_00973_),
    .B(_00975_),
    .Y(_00977_));
 sky130_fd_sc_hd__nor2_1 _07881_ (.A(_00976_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__o22a_1 _07882_ (.A1(_00242_),
    .A2(net26),
    .B1(net24),
    .B2(_00249_),
    .X(_00979_));
 sky130_fd_sc_hd__xnor2_1 _07883_ (.A(net87),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__a21oi_1 _07884_ (.A1(_00978_),
    .A2(_00980_),
    .B1(_00976_),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _07885_ (.A(_00971_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__o22a_1 _07886_ (.A1(net114),
    .A2(net85),
    .B1(net81),
    .B2(_00298_),
    .X(_00983_));
 sky130_fd_sc_hd__xnor2_2 _07887_ (.A(net137),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__o22a_1 _07888_ (.A1(net129),
    .A2(net73),
    .B1(net107),
    .B2(net77),
    .X(_00985_));
 sky130_fd_sc_hd__xnor2_1 _07889_ (.A(net121),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _07890_ (.A(_00984_),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__and3_1 _07891_ (.A(net292),
    .B(_00146_),
    .C(_00147_),
    .X(_00988_));
 sky130_fd_sc_hd__a21oi_1 _07892_ (.A1(_00154_),
    .A2(_00155_),
    .B1(net237),
    .Y(_00989_));
 sky130_fd_sc_hd__o21ai_1 _07893_ (.A1(_00988_),
    .A2(_00989_),
    .B1(net240),
    .Y(_00990_));
 sky130_fd_sc_hd__or3_1 _07894_ (.A(net240),
    .B(_00988_),
    .C(_00989_),
    .X(_00991_));
 sky130_fd_sc_hd__o22a_1 _07895_ (.A1(net155),
    .A2(net83),
    .B1(net79),
    .B2(net153),
    .X(_00992_));
 sky130_fd_sc_hd__xnor2_1 _07896_ (.A(_06507_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__and3_1 _07897_ (.A(_00990_),
    .B(_00991_),
    .C(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__a22o_1 _07898_ (.A1(_06532_),
    .A2(net102),
    .B1(_00174_),
    .B2(_06540_),
    .X(_00995_));
 sky130_fd_sc_hd__xnor2_1 _07899_ (.A(net192),
    .B(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__a21oi_1 _07900_ (.A1(_00990_),
    .A2(_00991_),
    .B1(_00993_),
    .Y(_00997_));
 sky130_fd_sc_hd__a21o_1 _07901_ (.A1(_00990_),
    .A2(_00991_),
    .B1(_00993_),
    .X(_00998_));
 sky130_fd_sc_hd__or3b_1 _07902_ (.A(_00994_),
    .B(_00997_),
    .C_N(_00996_),
    .X(_00999_));
 sky130_fd_sc_hd__a21oi_1 _07903_ (.A1(_00996_),
    .A2(_00998_),
    .B1(_00994_),
    .Y(_01000_));
 sky130_fd_sc_hd__o22a_1 _07904_ (.A1(net147),
    .A2(net75),
    .B1(net71),
    .B2(net145),
    .X(_01001_));
 sky130_fd_sc_hd__xnor2_1 _07905_ (.A(net190),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__o22a_1 _07906_ (.A1(net110),
    .A2(net106),
    .B1(net104),
    .B2(net109),
    .X(_01003_));
 sky130_fd_sc_hd__xnor2_1 _07907_ (.A(net136),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__xor2_1 _07908_ (.A(_01002_),
    .B(_01004_),
    .X(_01005_));
 sky130_fd_sc_hd__o22a_1 _07909_ (.A1(net134),
    .A2(net119),
    .B1(net116),
    .B2(net131),
    .X(_01006_));
 sky130_fd_sc_hd__xnor2_1 _07910_ (.A(net622),
    .B(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__and2b_1 _07911_ (.A_N(_01007_),
    .B(_01005_),
    .X(_01008_));
 sky130_fd_sc_hd__o21bai_1 _07912_ (.A1(_01002_),
    .A2(_01004_),
    .B1_N(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__xnor2_1 _07913_ (.A(_00987_),
    .B(_01000_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _07914_ (.A(_01009_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__o31ai_2 _07915_ (.A1(_00984_),
    .A2(_00986_),
    .A3(_01000_),
    .B1(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__xor2_1 _07916_ (.A(_00971_),
    .B(_00981_),
    .X(_01013_));
 sky130_fd_sc_hd__a21o_1 _07917_ (.A1(_01012_),
    .A2(_01013_),
    .B1(_00982_),
    .X(_01014_));
 sky130_fd_sc_hd__xor2_2 _07918_ (.A(_00943_),
    .B(_00944_),
    .X(_01015_));
 sky130_fd_sc_hd__xnor2_1 _07919_ (.A(_00907_),
    .B(_00909_),
    .Y(_01016_));
 sky130_fd_sc_hd__xor2_1 _07920_ (.A(_00911_),
    .B(_00923_),
    .X(_01017_));
 sky130_fd_sc_hd__xnor2_1 _07921_ (.A(_00941_),
    .B(_00942_),
    .Y(_01018_));
 sky130_fd_sc_hd__xnor2_1 _07922_ (.A(_01016_),
    .B(_01017_),
    .Y(_01019_));
 sky130_fd_sc_hd__or2_1 _07923_ (.A(_01018_),
    .B(_01019_),
    .X(_01020_));
 sky130_fd_sc_hd__a21bo_1 _07924_ (.A1(_01016_),
    .A2(_01017_),
    .B1_N(_01020_),
    .X(_01021_));
 sky130_fd_sc_hd__xnor2_2 _07925_ (.A(_01014_),
    .B(_01015_),
    .Y(_01022_));
 sky130_fd_sc_hd__and2b_1 _07926_ (.A_N(_01022_),
    .B(_01021_),
    .X(_01023_));
 sky130_fd_sc_hd__a21o_2 _07927_ (.A1(_01014_),
    .A2(_01015_),
    .B1(_01023_),
    .X(_01024_));
 sky130_fd_sc_hd__xnor2_4 _07928_ (.A(_00960_),
    .B(_00961_),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2b_1 _07929_ (.A_N(_01025_),
    .B(_01024_),
    .Y(_01026_));
 sky130_fd_sc_hd__or3_1 _07930_ (.A(_00946_),
    .B(_00954_),
    .C(_00955_),
    .X(_01027_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_00956_),
    .B(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__and3_1 _07932_ (.A(_00962_),
    .B(_01026_),
    .C(_01028_),
    .X(_01029_));
 sky130_fd_sc_hd__a21o_1 _07933_ (.A1(_00962_),
    .A2(_01026_),
    .B1(_01028_),
    .X(_01030_));
 sky130_fd_sc_hd__nand2b_4 _07934_ (.A_N(_01029_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__and2_1 _07935_ (.A(_00949_),
    .B(_00950_),
    .X(_01032_));
 sky130_fd_sc_hd__nor2_1 _07936_ (.A(_00951_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__xnor2_2 _07937_ (.A(_01021_),
    .B(_01022_),
    .Y(_01034_));
 sky130_fd_sc_hd__and2_1 _07938_ (.A(_01033_),
    .B(_01034_),
    .X(_01035_));
 sky130_fd_sc_hd__or2_1 _07939_ (.A(_01033_),
    .B(_01034_),
    .X(_01036_));
 sky130_fd_sc_hd__xnor2_2 _07940_ (.A(_01033_),
    .B(_01034_),
    .Y(_01037_));
 sky130_fd_sc_hd__xnor2_1 _07941_ (.A(_01012_),
    .B(_01013_),
    .Y(_01038_));
 sky130_fd_sc_hd__o22a_1 _07942_ (.A1(net127),
    .A2(net34),
    .B1(net32),
    .B2(net141),
    .X(_01039_));
 sky130_fd_sc_hd__xnor2_1 _07943_ (.A(net125),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand2_1 _07944_ (.A(net208),
    .B(net30),
    .Y(_01041_));
 sky130_fd_sc_hd__xnor2_1 _07945_ (.A(net48),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__and2b_1 _07946_ (.A_N(_01042_),
    .B(_01040_),
    .X(_01043_));
 sky130_fd_sc_hd__xor2_1 _07947_ (.A(_01040_),
    .B(_01042_),
    .X(_01044_));
 sky130_fd_sc_hd__o22a_1 _07948_ (.A1(net140),
    .A2(net26),
    .B1(net24),
    .B2(net142),
    .X(_01045_));
 sky130_fd_sc_hd__xnor2_1 _07949_ (.A(net87),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__and2b_1 _07950_ (.A_N(_01044_),
    .B(_01046_),
    .X(_01047_));
 sky130_fd_sc_hd__or2_1 _07951_ (.A(_01043_),
    .B(_01047_),
    .X(_01048_));
 sky130_fd_sc_hd__o21bai_1 _07952_ (.A1(_00994_),
    .A2(_00997_),
    .B1_N(_00996_),
    .Y(_01049_));
 sky130_fd_sc_hd__and2_1 _07953_ (.A(_00984_),
    .B(_00986_),
    .X(_01050_));
 sky130_fd_sc_hd__nor2_1 _07954_ (.A(_00987_),
    .B(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__and3_1 _07955_ (.A(_00999_),
    .B(_01049_),
    .C(_01051_),
    .X(_01052_));
 sky130_fd_sc_hd__and2b_1 _07956_ (.A_N(_01005_),
    .B(_01007_),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _07957_ (.A(_01008_),
    .B(_01053_),
    .X(_01054_));
 sky130_fd_sc_hd__a21oi_1 _07958_ (.A1(_00999_),
    .A2(_01049_),
    .B1(_01051_),
    .Y(_01055_));
 sky130_fd_sc_hd__or3_1 _07959_ (.A(_01052_),
    .B(_01054_),
    .C(_01055_),
    .X(_01056_));
 sky130_fd_sc_hd__o21ba_1 _07960_ (.A1(_01054_),
    .A2(_01055_),
    .B1_N(_01052_),
    .X(_01057_));
 sky130_fd_sc_hd__o21ba_1 _07961_ (.A1(_01043_),
    .A2(_01047_),
    .B1_N(_01057_),
    .X(_01058_));
 sky130_fd_sc_hd__o22a_1 _07962_ (.A1(net144),
    .A2(net119),
    .B1(net71),
    .B2(net146),
    .X(_01059_));
 sky130_fd_sc_hd__xnor2_1 _07963_ (.A(net188),
    .B(_01059_),
    .Y(_01060_));
 sky130_fd_sc_hd__o22a_1 _07964_ (.A1(net133),
    .A2(net116),
    .B1(net110),
    .B2(net131),
    .X(_01061_));
 sky130_fd_sc_hd__xnor2_1 _07965_ (.A(net171),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__or2_1 _07966_ (.A(_01060_),
    .B(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__a21o_1 _07967_ (.A1(_00154_),
    .A2(_00155_),
    .B1(net287),
    .X(_01064_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(_06494_),
    .B(net102),
    .Y(_01065_));
 sky130_fd_sc_hd__a21oi_1 _07969_ (.A1(_01064_),
    .A2(_01065_),
    .B1(net238),
    .Y(_01066_));
 sky130_fd_sc_hd__and3_1 _07970_ (.A(net238),
    .B(_01064_),
    .C(_01065_),
    .X(_01067_));
 sky130_fd_sc_hd__o22a_1 _07971_ (.A1(net154),
    .A2(net79),
    .B1(net75),
    .B2(net152),
    .X(_01068_));
 sky130_fd_sc_hd__xnor2_1 _07972_ (.A(net195),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__or3_2 _07973_ (.A(_01066_),
    .B(_01067_),
    .C(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__o22a_1 _07974_ (.A1(net150),
    .A2(net98),
    .B1(net83),
    .B2(net148),
    .X(_01071_));
 sky130_fd_sc_hd__xnor2_1 _07975_ (.A(net193),
    .B(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__o21ai_1 _07976_ (.A1(_01066_),
    .A2(_01067_),
    .B1(_01069_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand3b_2 _07977_ (.A_N(_01072_),
    .B(_01073_),
    .C(_01070_),
    .Y(_01074_));
 sky130_fd_sc_hd__xnor2_1 _07978_ (.A(net48),
    .B(_01063_),
    .Y(_01075_));
 sky130_fd_sc_hd__a21o_1 _07979_ (.A1(_01070_),
    .A2(_01074_),
    .B1(_01075_),
    .X(_01076_));
 sky130_fd_sc_hd__o21ai_1 _07980_ (.A1(net48),
    .A2(_01063_),
    .B1(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__xnor2_1 _07981_ (.A(_01048_),
    .B(_01057_),
    .Y(_01078_));
 sky130_fd_sc_hd__a21o_1 _07982_ (.A1(_01077_),
    .A2(_01078_),
    .B1(_01058_),
    .X(_01079_));
 sky130_fd_sc_hd__nand2b_1 _07983_ (.A_N(_01038_),
    .B(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__o21ai_1 _07984_ (.A1(_00966_),
    .A2(_00967_),
    .B1(_00969_),
    .Y(_01081_));
 sky130_fd_sc_hd__xor2_1 _07985_ (.A(_00978_),
    .B(_00980_),
    .X(_01082_));
 sky130_fd_sc_hd__and3_1 _07986_ (.A(_00970_),
    .B(_01081_),
    .C(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__a21oi_1 _07987_ (.A1(_00970_),
    .A2(_01081_),
    .B1(_01082_),
    .Y(_01084_));
 sky130_fd_sc_hd__xnor2_1 _07988_ (.A(_01009_),
    .B(_01010_),
    .Y(_01085_));
 sky130_fd_sc_hd__nor3_1 _07989_ (.A(_01083_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nor2_1 _07990_ (.A(_01083_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__xnor2_1 _07991_ (.A(_01038_),
    .B(_01079_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2b_1 _07992_ (.A_N(_01087_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_2 _07993_ (.A(_01080_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__a21o_2 _07994_ (.A1(_01036_),
    .A2(_01090_),
    .B1(_01035_),
    .X(_01091_));
 sky130_fd_sc_hd__xnor2_4 _07995_ (.A(_01024_),
    .B(_01025_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _07996_ (.A(_01091_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__xnor2_4 _07997_ (.A(_01091_),
    .B(_01092_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(_01018_),
    .B(_01019_),
    .Y(_01095_));
 sky130_fd_sc_hd__and2_1 _07999_ (.A(_01020_),
    .B(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__xnor2_1 _08000_ (.A(_01087_),
    .B(_01088_),
    .Y(_01097_));
 sky130_fd_sc_hd__and2_1 _08001_ (.A(_01096_),
    .B(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__o22a_1 _08002_ (.A1(net146),
    .A2(net119),
    .B1(net116),
    .B2(net144),
    .X(_01099_));
 sky130_fd_sc_hd__xnor2_1 _08003_ (.A(net188),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__o22a_1 _08004_ (.A1(net133),
    .A2(net110),
    .B1(net108),
    .B2(net131),
    .X(_01101_));
 sky130_fd_sc_hd__xnor2_1 _08005_ (.A(net171),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__or2_1 _08006_ (.A(_01100_),
    .B(_01102_),
    .X(_01103_));
 sky130_fd_sc_hd__xnor2_1 _08007_ (.A(_01060_),
    .B(_01062_),
    .Y(_01104_));
 sky130_fd_sc_hd__nor2_1 _08008_ (.A(_01103_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__xor2_1 _08009_ (.A(_01103_),
    .B(_01104_),
    .X(_01106_));
 sky130_fd_sc_hd__a21bo_1 _08010_ (.A1(_01070_),
    .A2(_01073_),
    .B1_N(_01072_),
    .X(_01107_));
 sky130_fd_sc_hd__nand3_1 _08011_ (.A(_01074_),
    .B(_01106_),
    .C(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__and2b_1 _08012_ (.A_N(_01105_),
    .B(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__a31o_1 _08013_ (.A1(_01074_),
    .A2(_01106_),
    .A3(_01107_),
    .B1(_01105_),
    .X(_01110_));
 sky130_fd_sc_hd__o22a_1 _08014_ (.A1(net108),
    .A2(net106),
    .B1(net104),
    .B2(net114),
    .X(_01111_));
 sky130_fd_sc_hd__xnor2_1 _08015_ (.A(net136),
    .B(_01111_),
    .Y(_01112_));
 sky130_fd_sc_hd__o22a_1 _08016_ (.A1(net129),
    .A2(net78),
    .B1(net74),
    .B2(net127),
    .X(_01113_));
 sky130_fd_sc_hd__xnor2_1 _08017_ (.A(net123),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__o22a_1 _08018_ (.A1(net113),
    .A2(net86),
    .B1(net82),
    .B2(net107),
    .X(_01115_));
 sky130_fd_sc_hd__xnor2_1 _08019_ (.A(net138),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__xnor2_1 _08020_ (.A(_01112_),
    .B(_01114_),
    .Y(_01117_));
 sky130_fd_sc_hd__or2_1 _08021_ (.A(_01116_),
    .B(_01117_),
    .X(_01118_));
 sky130_fd_sc_hd__o21a_1 _08022_ (.A1(_01112_),
    .A2(_01114_),
    .B1(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__o22a_1 _08023_ (.A1(net287),
    .A2(net100),
    .B1(net98),
    .B2(net237),
    .X(_01120_));
 sky130_fd_sc_hd__xnor2_2 _08024_ (.A(net238),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__o22a_1 _08025_ (.A1(net154),
    .A2(net75),
    .B1(net71),
    .B2(net152),
    .X(_01122_));
 sky130_fd_sc_hd__xnor2_2 _08026_ (.A(net195),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__or2_1 _08027_ (.A(_01121_),
    .B(_01123_),
    .X(_01124_));
 sky130_fd_sc_hd__o22a_1 _08028_ (.A1(net150),
    .A2(net83),
    .B1(net79),
    .B2(net148),
    .X(_01125_));
 sky130_fd_sc_hd__xnor2_2 _08029_ (.A(net191),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__xnor2_2 _08030_ (.A(_01121_),
    .B(_01123_),
    .Y(_01127_));
 sky130_fd_sc_hd__o21ai_2 _08031_ (.A1(_01126_),
    .A2(_01127_),
    .B1(_01124_),
    .Y(_01128_));
 sky130_fd_sc_hd__o22a_1 _08032_ (.A1(net141),
    .A2(net34),
    .B1(net32),
    .B2(net140),
    .X(_01129_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(net125),
    .B(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(_01128_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__xnor2_1 _08035_ (.A(_01128_),
    .B(_01130_),
    .Y(_01132_));
 sky130_fd_sc_hd__o22a_1 _08036_ (.A1(net142),
    .A2(net26),
    .B1(net24),
    .B2(net209),
    .X(_01133_));
 sky130_fd_sc_hd__xnor2_1 _08037_ (.A(net87),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__inv_2 _08038_ (.A(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__o21a_1 _08039_ (.A1(_01132_),
    .A2(_01135_),
    .B1(_01131_),
    .X(_01136_));
 sky130_fd_sc_hd__xnor2_2 _08040_ (.A(_01110_),
    .B(_01119_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2b_1 _08041_ (.A_N(_01136_),
    .B(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__o21ai_1 _08042_ (.A1(_01109_),
    .A2(_01119_),
    .B1(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__xnor2_1 _08043_ (.A(_01077_),
    .B(_01078_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2b_1 _08044_ (.A_N(_01140_),
    .B(_01139_),
    .Y(_01141_));
 sky130_fd_sc_hd__and2b_1 _08045_ (.A_N(_01046_),
    .B(_01044_),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_1 _08046_ (.A(_01047_),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__o21ai_1 _08047_ (.A1(_01052_),
    .A2(_01055_),
    .B1(_01054_),
    .Y(_01144_));
 sky130_fd_sc_hd__and3_1 _08048_ (.A(_01056_),
    .B(_01143_),
    .C(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__nand3_1 _08049_ (.A(_01070_),
    .B(_01074_),
    .C(_01075_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_01076_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__a21oi_1 _08051_ (.A1(_01056_),
    .A2(_01144_),
    .B1(_01143_),
    .Y(_01148_));
 sky130_fd_sc_hd__or3_1 _08052_ (.A(_01145_),
    .B(_01147_),
    .C(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__and2b_1 _08053_ (.A_N(_01145_),
    .B(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__xnor2_1 _08054_ (.A(_01139_),
    .B(_01140_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2b_1 _08055_ (.A_N(_01150_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _08056_ (.A(_01141_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__xor2_1 _08057_ (.A(_01096_),
    .B(_01097_),
    .X(_01154_));
 sky130_fd_sc_hd__a21o_1 _08058_ (.A1(_01153_),
    .A2(_01154_),
    .B1(_01098_),
    .X(_01155_));
 sky130_fd_sc_hd__xnor2_4 _08059_ (.A(_01037_),
    .B(_01090_),
    .Y(_01156_));
 sky130_fd_sc_hd__xnor2_2 _08060_ (.A(_01155_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__or2_1 _08061_ (.A(_01094_),
    .B(_01157_),
    .X(_01158_));
 sky130_fd_sc_hd__o21ai_1 _08062_ (.A1(_01145_),
    .A2(_01148_),
    .B1(_01147_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_2 _08063_ (.A(_01149_),
    .B(_01159_),
    .Y(_01160_));
 sky130_fd_sc_hd__a21o_1 _08064_ (.A1(_01074_),
    .A2(_01107_),
    .B1(_01106_),
    .X(_01161_));
 sky130_fd_sc_hd__nand2_1 _08065_ (.A(_01116_),
    .B(_01117_),
    .Y(_01162_));
 sky130_fd_sc_hd__and2_1 _08066_ (.A(_01118_),
    .B(_01162_),
    .X(_01163_));
 sky130_fd_sc_hd__and3_1 _08067_ (.A(_01108_),
    .B(_01161_),
    .C(_01163_),
    .X(_01164_));
 sky130_fd_sc_hd__a21oi_1 _08068_ (.A1(_01108_),
    .A2(_01161_),
    .B1(_01163_),
    .Y(_01165_));
 sky130_fd_sc_hd__xnor2_1 _08069_ (.A(_01132_),
    .B(_01135_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor3_1 _08070_ (.A(_01164_),
    .B(_01165_),
    .C(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__or2_1 _08071_ (.A(_01164_),
    .B(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__xnor2_2 _08072_ (.A(_01136_),
    .B(_01137_),
    .Y(_01169_));
 sky130_fd_sc_hd__o22a_1 _08073_ (.A1(net287),
    .A2(net98),
    .B1(net83),
    .B2(net237),
    .X(_01170_));
 sky130_fd_sc_hd__xnor2_1 _08074_ (.A(net238),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__o22a_1 _08075_ (.A1(net150),
    .A2(net79),
    .B1(net75),
    .B2(net148),
    .X(_01172_));
 sky130_fd_sc_hd__xnor2_1 _08076_ (.A(net191),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__or2_1 _08077_ (.A(_01171_),
    .B(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_01100_),
    .B(_01102_),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _08079_ (.A(_01103_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _08080_ (.A(_01174_),
    .B(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_01174_),
    .B(_01176_),
    .Y(_01178_));
 sky130_fd_sc_hd__xnor2_1 _08082_ (.A(_01174_),
    .B(_01176_),
    .Y(_01179_));
 sky130_fd_sc_hd__xor2_2 _08083_ (.A(_01126_),
    .B(_01127_),
    .X(_01180_));
 sky130_fd_sc_hd__a21o_1 _08084_ (.A1(_01178_),
    .A2(_01180_),
    .B1(_01177_),
    .X(_01181_));
 sky130_fd_sc_hd__o22a_1 _08085_ (.A1(net114),
    .A2(net106),
    .B1(net104),
    .B2(net113),
    .X(_01182_));
 sky130_fd_sc_hd__xnor2_1 _08086_ (.A(net136),
    .B(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__o22a_1 _08087_ (.A1(net127),
    .A2(net78),
    .B1(net74),
    .B2(net141),
    .X(_01184_));
 sky130_fd_sc_hd__xnor2_1 _08088_ (.A(net123),
    .B(_01184_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _08089_ (.A(_01183_),
    .B(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__o22a_1 _08090_ (.A1(net129),
    .A2(net82),
    .B1(net107),
    .B2(net86),
    .X(_01187_));
 sky130_fd_sc_hd__xnor2_1 _08091_ (.A(net138),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__xnor2_1 _08092_ (.A(_01183_),
    .B(_01185_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_1 _08093_ (.A(_01188_),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _08094_ (.A(_01186_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__o21a_1 _08095_ (.A1(_01186_),
    .A2(_01190_),
    .B1(_01181_),
    .X(_01192_));
 sky130_fd_sc_hd__nor2_1 _08096_ (.A(net209),
    .B(net26),
    .Y(_01193_));
 sky130_fd_sc_hd__o22a_1 _08097_ (.A1(net140),
    .A2(net34),
    .B1(net32),
    .B2(net142),
    .X(_01194_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(net125),
    .B(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__mux2_2 _08099_ (.A0(net87),
    .A1(_01195_),
    .S(_01193_),
    .X(_01196_));
 sky130_fd_sc_hd__xnor2_2 _08100_ (.A(_01181_),
    .B(_01191_),
    .Y(_01197_));
 sky130_fd_sc_hd__a21oi_2 _08101_ (.A1(_01196_),
    .A2(_01197_),
    .B1(_01192_),
    .Y(_01198_));
 sky130_fd_sc_hd__and2b_1 _08102_ (.A_N(_01198_),
    .B(_01169_),
    .X(_01199_));
 sky130_fd_sc_hd__xnor2_2 _08103_ (.A(_01169_),
    .B(_01198_),
    .Y(_01200_));
 sky130_fd_sc_hd__xnor2_2 _08104_ (.A(_01168_),
    .B(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__xor2_2 _08105_ (.A(_01196_),
    .B(_01197_),
    .X(_01202_));
 sky130_fd_sc_hd__xor2_1 _08106_ (.A(_01171_),
    .B(_01173_),
    .X(_01203_));
 sky130_fd_sc_hd__o22a_1 _08107_ (.A1(net142),
    .A2(net34),
    .B1(net32),
    .B2(net209),
    .X(_01204_));
 sky130_fd_sc_hd__xnor2_1 _08108_ (.A(net125),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__and2_1 _08109_ (.A(_01203_),
    .B(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__o22a_1 _08110_ (.A1(net287),
    .A2(net83),
    .B1(net79),
    .B2(net237),
    .X(_01207_));
 sky130_fd_sc_hd__xnor2_2 _08111_ (.A(net238),
    .B(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__o22a_1 _08112_ (.A1(net150),
    .A2(net75),
    .B1(net71),
    .B2(net148),
    .X(_01209_));
 sky130_fd_sc_hd__xnor2_2 _08113_ (.A(net191),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _08114_ (.A(_01208_),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__xor2_1 _08115_ (.A(_01203_),
    .B(_01205_),
    .X(_01212_));
 sky130_fd_sc_hd__and2_1 _08116_ (.A(_01211_),
    .B(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__a21o_1 _08117_ (.A1(_01211_),
    .A2(_01212_),
    .B1(_01206_),
    .X(_01214_));
 sky130_fd_sc_hd__o22a_1 _08118_ (.A1(net131),
    .A2(net114),
    .B1(net108),
    .B2(net133),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_1 _08119_ (.A(net171),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__o22a_1 _08120_ (.A1(net152),
    .A2(net119),
    .B1(net71),
    .B2(net154),
    .X(_01217_));
 sky130_fd_sc_hd__xnor2_1 _08121_ (.A(net195),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__o22a_1 _08122_ (.A1(net146),
    .A2(net116),
    .B1(net110),
    .B2(net144),
    .X(_01219_));
 sky130_fd_sc_hd__xnor2_1 _08123_ (.A(net188),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__xnor2_1 _08124_ (.A(_01216_),
    .B(_01218_),
    .Y(_01221_));
 sky130_fd_sc_hd__or2_1 _08125_ (.A(_01220_),
    .B(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__o21a_1 _08126_ (.A1(_01216_),
    .A2(_01218_),
    .B1(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__o21ba_1 _08127_ (.A1(_01206_),
    .A2(_01213_),
    .B1_N(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__o22a_1 _08128_ (.A1(net113),
    .A2(net106),
    .B1(net104),
    .B2(net107),
    .X(_01225_));
 sky130_fd_sc_hd__xnor2_2 _08129_ (.A(net136),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__o22a_1 _08130_ (.A1(net141),
    .A2(net78),
    .B1(net74),
    .B2(net140),
    .X(_01227_));
 sky130_fd_sc_hd__xnor2_1 _08131_ (.A(net123),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__o22a_1 _08132_ (.A1(net129),
    .A2(net86),
    .B1(net82),
    .B2(net127),
    .X(_01229_));
 sky130_fd_sc_hd__xnor2_1 _08133_ (.A(net138),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__xnor2_1 _08134_ (.A(_01226_),
    .B(_01228_),
    .Y(_01231_));
 sky130_fd_sc_hd__or2_1 _08135_ (.A(_01230_),
    .B(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__o21ai_2 _08136_ (.A1(_01226_),
    .A2(_01228_),
    .B1(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2b_1 _08137_ (.A_N(_01214_),
    .B(_01223_),
    .Y(_01234_));
 sky130_fd_sc_hd__xor2_1 _08138_ (.A(_01214_),
    .B(_01223_),
    .X(_01235_));
 sky130_fd_sc_hd__a21o_1 _08139_ (.A1(_01233_),
    .A2(_01234_),
    .B1(_01224_),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_2 _08140_ (.A(_01179_),
    .B(_01180_),
    .Y(_01237_));
 sky130_fd_sc_hd__and2_1 _08141_ (.A(_01188_),
    .B(_01189_),
    .X(_01238_));
 sky130_fd_sc_hd__nor2_1 _08142_ (.A(_01190_),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__xnor2_1 _08143_ (.A(_01237_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__xnor2_1 _08144_ (.A(_01193_),
    .B(_01195_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_1 _08145_ (.A(_01240_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__a21oi_2 _08146_ (.A1(_01237_),
    .A2(_01239_),
    .B1(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__xor2_2 _08147_ (.A(_01202_),
    .B(_01236_),
    .X(_01244_));
 sky130_fd_sc_hd__nand2b_1 _08148_ (.A_N(_01243_),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__a21bo_1 _08149_ (.A1(_01202_),
    .A2(_01236_),
    .B1_N(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_2 _08150_ (.A(_01160_),
    .B(_01201_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2b_1 _08151_ (.A_N(_01247_),
    .B(_01246_),
    .Y(_01248_));
 sky130_fd_sc_hd__o21ai_2 _08152_ (.A1(_01160_),
    .A2(_01201_),
    .B1(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__o21a_1 _08153_ (.A1(_01083_),
    .A2(_01084_),
    .B1(_01085_),
    .X(_01250_));
 sky130_fd_sc_hd__nor2_2 _08154_ (.A(_01086_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__xnor2_1 _08155_ (.A(_01150_),
    .B(_01151_),
    .Y(_01252_));
 sky130_fd_sc_hd__and2_1 _08156_ (.A(_01251_),
    .B(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__xor2_2 _08157_ (.A(_01251_),
    .B(_01252_),
    .X(_01254_));
 sky130_fd_sc_hd__a21o_1 _08158_ (.A1(_01168_),
    .A2(_01200_),
    .B1(_01199_),
    .X(_01255_));
 sky130_fd_sc_hd__xor2_2 _08159_ (.A(_01254_),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__nor2_1 _08160_ (.A(_01249_),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_01249_),
    .B(_01256_),
    .Y(_01258_));
 sky130_fd_sc_hd__xnor2_1 _08162_ (.A(_01249_),
    .B(_01256_),
    .Y(_01259_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_01254_),
    .A2(_01255_),
    .B1(_01253_),
    .X(_01260_));
 sky130_fd_sc_hd__xnor2_1 _08164_ (.A(_01153_),
    .B(_01154_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2b_1 _08165_ (.A_N(_01261_),
    .B(_01260_),
    .Y(_01262_));
 sky130_fd_sc_hd__and2b_1 _08166_ (.A_N(_01260_),
    .B(_01261_),
    .X(_01263_));
 sky130_fd_sc_hd__xor2_1 _08167_ (.A(_01260_),
    .B(_01261_),
    .X(_01264_));
 sky130_fd_sc_hd__or2_1 _08168_ (.A(_01259_),
    .B(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__o21a_1 _08169_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_01166_),
    .X(_01266_));
 sky130_fd_sc_hd__nor2_1 _08170_ (.A(_01167_),
    .B(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__xnor2_2 _08171_ (.A(_01243_),
    .B(_01244_),
    .Y(_01268_));
 sky130_fd_sc_hd__and2_1 _08172_ (.A(_01267_),
    .B(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__xor2_2 _08173_ (.A(_01267_),
    .B(_01268_),
    .X(_01270_));
 sky130_fd_sc_hd__o22a_1 _08174_ (.A1(net133),
    .A2(net114),
    .B1(net113),
    .B2(net131),
    .X(_01271_));
 sky130_fd_sc_hd__xnor2_1 _08175_ (.A(net171),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__o22a_1 _08176_ (.A1(net154),
    .A2(net119),
    .B1(net116),
    .B2(net152),
    .X(_01273_));
 sky130_fd_sc_hd__xnor2_1 _08177_ (.A(net195),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__xnor2_1 _08178_ (.A(_01272_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__o22a_1 _08179_ (.A1(net146),
    .A2(net110),
    .B1(net108),
    .B2(net144),
    .X(_01276_));
 sky130_fd_sc_hd__xnor2_1 _08180_ (.A(net188),
    .B(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_1 _08181_ (.A(_01275_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__o21ba_1 _08182_ (.A1(_01272_),
    .A2(_01274_),
    .B1_N(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__xor2_2 _08183_ (.A(_01208_),
    .B(_01210_),
    .X(_01280_));
 sky130_fd_sc_hd__nor2_1 _08184_ (.A(net209),
    .B(net34),
    .Y(_01281_));
 sky130_fd_sc_hd__mux2_1 _08185_ (.A0(net125),
    .A1(_01280_),
    .S(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__and2b_1 _08186_ (.A_N(_01279_),
    .B(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__o22a_1 _08187_ (.A1(net107),
    .A2(net106),
    .B1(net104),
    .B2(net129),
    .X(_01284_));
 sky130_fd_sc_hd__xnor2_2 _08188_ (.A(net136),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__o22a_1 _08189_ (.A1(net140),
    .A2(net78),
    .B1(net74),
    .B2(net142),
    .X(_01286_));
 sky130_fd_sc_hd__xnor2_2 _08190_ (.A(net123),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__o22a_1 _08191_ (.A1(net127),
    .A2(net86),
    .B1(net82),
    .B2(net141),
    .X(_01288_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(net138),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__xnor2_1 _08193_ (.A(_01285_),
    .B(_01287_),
    .Y(_01290_));
 sky130_fd_sc_hd__or2_1 _08194_ (.A(_01289_),
    .B(_01290_),
    .X(_01291_));
 sky130_fd_sc_hd__o21ai_2 _08195_ (.A1(_01285_),
    .A2(_01287_),
    .B1(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__xnor2_2 _08196_ (.A(_01279_),
    .B(_01282_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21oi_2 _08197_ (.A1(_01292_),
    .A2(_01293_),
    .B1(_01283_),
    .Y(_01294_));
 sky130_fd_sc_hd__xnor2_2 _08198_ (.A(_01233_),
    .B(_01235_),
    .Y(_01295_));
 sky130_fd_sc_hd__and2b_1 _08199_ (.A_N(_01294_),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__nor2_1 _08200_ (.A(_01211_),
    .B(_01212_),
    .Y(_01297_));
 sky130_fd_sc_hd__or2_1 _08201_ (.A(_01213_),
    .B(_01297_),
    .X(_01298_));
 sky130_fd_sc_hd__nand2_1 _08202_ (.A(_01220_),
    .B(_01221_),
    .Y(_01299_));
 sky130_fd_sc_hd__and2_1 _08203_ (.A(_01222_),
    .B(_01299_),
    .X(_01300_));
 sky130_fd_sc_hd__or3b_1 _08204_ (.A(_01213_),
    .B(_01297_),
    .C_N(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(_01230_),
    .B(_01231_),
    .Y(_01302_));
 sky130_fd_sc_hd__and2_1 _08206_ (.A(_01232_),
    .B(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__xnor2_1 _08207_ (.A(_01298_),
    .B(_01300_),
    .Y(_01304_));
 sky130_fd_sc_hd__a21bo_1 _08208_ (.A1(_01303_),
    .A2(_01304_),
    .B1_N(_01301_),
    .X(_01305_));
 sky130_fd_sc_hd__xnor2_2 _08209_ (.A(_01294_),
    .B(_01295_),
    .Y(_01306_));
 sky130_fd_sc_hd__a21o_1 _08210_ (.A1(_01305_),
    .A2(_01306_),
    .B1(_01296_),
    .X(_01307_));
 sky130_fd_sc_hd__a21oi_2 _08211_ (.A1(_01270_),
    .A2(_01307_),
    .B1(_01269_),
    .Y(_01308_));
 sky130_fd_sc_hd__xor2_2 _08212_ (.A(_01246_),
    .B(_01247_),
    .X(_01309_));
 sky130_fd_sc_hd__and2_1 _08213_ (.A(_01308_),
    .B(_01309_),
    .X(_01310_));
 sky130_fd_sc_hd__or2_1 _08214_ (.A(_01308_),
    .B(_01309_),
    .X(_01311_));
 sky130_fd_sc_hd__and2_1 _08215_ (.A(_01240_),
    .B(_01241_),
    .X(_01312_));
 sky130_fd_sc_hd__or2_1 _08216_ (.A(_01242_),
    .B(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__xnor2_2 _08217_ (.A(_01305_),
    .B(_01306_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _08218_ (.A(_01313_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__xor2_2 _08219_ (.A(_01313_),
    .B(_01314_),
    .X(_01316_));
 sky130_fd_sc_hd__xnor2_1 _08220_ (.A(_01292_),
    .B(_01293_),
    .Y(_01317_));
 sky130_fd_sc_hd__o22a_1 _08221_ (.A1(net141),
    .A2(net86),
    .B1(net82),
    .B2(net140),
    .X(_01318_));
 sky130_fd_sc_hd__xnor2_1 _08222_ (.A(net138),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__o22a_1 _08223_ (.A1(net142),
    .A2(net78),
    .B1(net74),
    .B2(net209),
    .X(_01320_));
 sky130_fd_sc_hd__xnor2_1 _08224_ (.A(net123),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_1 _08225_ (.A(_01319_),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__o22a_1 _08226_ (.A1(net287),
    .A2(net79),
    .B1(net75),
    .B2(net237),
    .X(_01323_));
 sky130_fd_sc_hd__xnor2_2 _08227_ (.A(net238),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__o22a_1 _08228_ (.A1(net154),
    .A2(net116),
    .B1(net110),
    .B2(net152),
    .X(_01325_));
 sky130_fd_sc_hd__xnor2_2 _08229_ (.A(net195),
    .B(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(_01324_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__xnor2_2 _08231_ (.A(_01324_),
    .B(_01326_),
    .Y(_01328_));
 sky130_fd_sc_hd__o22a_1 _08232_ (.A1(net148),
    .A2(net119),
    .B1(net71),
    .B2(net150),
    .X(_01329_));
 sky130_fd_sc_hd__xnor2_2 _08233_ (.A(net191),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__o21bai_2 _08234_ (.A1(_01328_),
    .A2(_01330_),
    .B1_N(_01327_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_01322_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__o22a_1 _08236_ (.A1(net129),
    .A2(net106),
    .B1(net104),
    .B2(net127),
    .X(_01333_));
 sky130_fd_sc_hd__xnor2_2 _08237_ (.A(net136),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__o22a_1 _08238_ (.A1(net144),
    .A2(net114),
    .B1(net108),
    .B2(net146),
    .X(_01335_));
 sky130_fd_sc_hd__xnor2_2 _08239_ (.A(net188),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__xor2_2 _08240_ (.A(_01334_),
    .B(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__o22a_1 _08241_ (.A1(net133),
    .A2(net113),
    .B1(net107),
    .B2(net131),
    .X(_01338_));
 sky130_fd_sc_hd__xnor2_2 _08242_ (.A(net171),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2b_1 _08243_ (.A_N(_01339_),
    .B(_01337_),
    .Y(_01340_));
 sky130_fd_sc_hd__o21ai_2 _08244_ (.A1(_01334_),
    .A2(_01336_),
    .B1(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__xor2_2 _08245_ (.A(_01322_),
    .B(_01331_),
    .X(_01342_));
 sky130_fd_sc_hd__a21boi_1 _08246_ (.A1(_01341_),
    .A2(_01342_),
    .B1_N(_01332_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _08247_ (.A(_01317_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__and2_1 _08248_ (.A(_01275_),
    .B(_01277_),
    .X(_01345_));
 sky130_fd_sc_hd__nor2_1 _08249_ (.A(_01278_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__xnor2_2 _08250_ (.A(_01280_),
    .B(_01281_),
    .Y(_01347_));
 sky130_fd_sc_hd__xnor2_1 _08251_ (.A(_01346_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_01289_),
    .B(_01290_),
    .Y(_01349_));
 sky130_fd_sc_hd__and2_1 _08253_ (.A(_01291_),
    .B(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_01348_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__o31ai_2 _08255_ (.A1(_01278_),
    .A2(_01345_),
    .A3(_01347_),
    .B1(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__xor2_1 _08256_ (.A(_01317_),
    .B(_01343_),
    .X(_01353_));
 sky130_fd_sc_hd__a21o_1 _08257_ (.A1(_01352_),
    .A2(_01353_),
    .B1(_01344_),
    .X(_01354_));
 sky130_fd_sc_hd__a21o_1 _08258_ (.A1(_01316_),
    .A2(_01354_),
    .B1(_01315_),
    .X(_01355_));
 sky130_fd_sc_hd__xor2_2 _08259_ (.A(_01270_),
    .B(_01307_),
    .X(_01356_));
 sky130_fd_sc_hd__nand2_1 _08260_ (.A(_01355_),
    .B(_01356_),
    .Y(_01357_));
 sky130_fd_sc_hd__a21o_1 _08261_ (.A1(_01311_),
    .A2(_01357_),
    .B1(_01310_),
    .X(_01358_));
 sky130_fd_sc_hd__xnor2_2 _08262_ (.A(_01308_),
    .B(_01309_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _08263_ (.A(_01355_),
    .B(_01356_),
    .Y(_01360_));
 sky130_fd_sc_hd__xor2_1 _08264_ (.A(_01355_),
    .B(_01356_),
    .X(_01361_));
 sky130_fd_sc_hd__xnor2_1 _08265_ (.A(_01355_),
    .B(_01356_),
    .Y(_01362_));
 sky130_fd_sc_hd__or2_1 _08266_ (.A(_01359_),
    .B(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__xor2_2 _08267_ (.A(_01316_),
    .B(_01354_),
    .X(_01364_));
 sky130_fd_sc_hd__xnor2_1 _08268_ (.A(_01303_),
    .B(_01304_),
    .Y(_01365_));
 sky130_fd_sc_hd__xnor2_1 _08269_ (.A(_01352_),
    .B(_01353_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _08270_ (.A(_01365_),
    .B(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__xnor2_2 _08271_ (.A(_01341_),
    .B(_01342_),
    .Y(_01368_));
 sky130_fd_sc_hd__o22a_1 _08272_ (.A1(net140),
    .A2(net86),
    .B1(net82),
    .B2(net142),
    .X(_01369_));
 sky130_fd_sc_hd__xnor2_1 _08273_ (.A(net138),
    .B(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _08274_ (.A(net209),
    .B(net78),
    .Y(_01371_));
 sky130_fd_sc_hd__xnor2_1 _08275_ (.A(net123),
    .B(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2b_1 _08276_ (.A_N(_01370_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__o22a_1 _08277_ (.A1(net287),
    .A2(net75),
    .B1(net71),
    .B2(net237),
    .X(_01374_));
 sky130_fd_sc_hd__xnor2_2 _08278_ (.A(net238),
    .B(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__o22a_1 _08279_ (.A1(net154),
    .A2(net110),
    .B1(net108),
    .B2(net152),
    .X(_01376_));
 sky130_fd_sc_hd__xnor2_2 _08280_ (.A(net195),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__or2_1 _08281_ (.A(_01375_),
    .B(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__xnor2_2 _08282_ (.A(_01375_),
    .B(_01377_),
    .Y(_01379_));
 sky130_fd_sc_hd__o22a_1 _08283_ (.A1(net150),
    .A2(net119),
    .B1(net116),
    .B2(net148),
    .X(_01380_));
 sky130_fd_sc_hd__xnor2_2 _08284_ (.A(net191),
    .B(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__o21a_1 _08285_ (.A1(_01379_),
    .A2(_01381_),
    .B1(_01378_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_1 _08286_ (.A(_01373_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__o22a_1 _08287_ (.A1(net127),
    .A2(net106),
    .B1(net104),
    .B2(net141),
    .X(_01384_));
 sky130_fd_sc_hd__xnor2_2 _08288_ (.A(net136),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__o22a_1 _08289_ (.A1(net146),
    .A2(net114),
    .B1(net113),
    .B2(net144),
    .X(_01386_));
 sky130_fd_sc_hd__xnor2_2 _08290_ (.A(net188),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_1 _08291_ (.A(_01385_),
    .B(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__o22a_1 _08292_ (.A1(net131),
    .A2(net129),
    .B1(net107),
    .B2(net133),
    .X(_01389_));
 sky130_fd_sc_hd__xnor2_1 _08293_ (.A(net171),
    .B(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__nand2b_1 _08294_ (.A_N(_01390_),
    .B(_01388_),
    .Y(_01391_));
 sky130_fd_sc_hd__o21ai_2 _08295_ (.A1(_01385_),
    .A2(_01387_),
    .B1(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__xor2_2 _08296_ (.A(_01373_),
    .B(_01382_),
    .X(_01393_));
 sky130_fd_sc_hd__a21oi_2 _08297_ (.A1(_01392_),
    .A2(_01393_),
    .B1(_01383_),
    .Y(_01394_));
 sky130_fd_sc_hd__xnor2_2 _08298_ (.A(_01328_),
    .B(_01330_),
    .Y(_01395_));
 sky130_fd_sc_hd__and2_1 _08299_ (.A(_01319_),
    .B(_01321_),
    .X(_01396_));
 sky130_fd_sc_hd__or2_2 _08300_ (.A(_01322_),
    .B(_01396_),
    .X(_01397_));
 sky130_fd_sc_hd__xnor2_2 _08301_ (.A(_01395_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__xnor2_2 _08302_ (.A(_01337_),
    .B(_01339_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2b_1 _08303_ (.A_N(_01398_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__o21ai_2 _08304_ (.A1(_01395_),
    .A2(_01397_),
    .B1(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__xnor2_2 _08305_ (.A(_01368_),
    .B(_01394_),
    .Y(_01402_));
 sky130_fd_sc_hd__and2b_1 _08306_ (.A_N(_01402_),
    .B(_01401_),
    .X(_01403_));
 sky130_fd_sc_hd__o21bai_2 _08307_ (.A1(_01368_),
    .A2(_01394_),
    .B1_N(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__xor2_1 _08308_ (.A(_01365_),
    .B(_01366_),
    .X(_01405_));
 sky130_fd_sc_hd__a21o_1 _08309_ (.A1(_01404_),
    .A2(_01405_),
    .B1(_01367_),
    .X(_01406_));
 sky130_fd_sc_hd__nor2_1 _08310_ (.A(_01364_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__nand2_1 _08311_ (.A(_01364_),
    .B(_01406_),
    .Y(_01408_));
 sky130_fd_sc_hd__or2_1 _08312_ (.A(_01348_),
    .B(_01350_),
    .X(_01409_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(_01351_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__xor2_2 _08314_ (.A(_01401_),
    .B(_01402_),
    .X(_01411_));
 sky130_fd_sc_hd__or2_1 _08315_ (.A(_01410_),
    .B(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__o22a_1 _08316_ (.A1(net146),
    .A2(net113),
    .B1(net107),
    .B2(net144),
    .X(_01413_));
 sky130_fd_sc_hd__xnor2_1 _08317_ (.A(net188),
    .B(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__o22a_1 _08318_ (.A1(net133),
    .A2(net129),
    .B1(net127),
    .B2(net131),
    .X(_01415_));
 sky130_fd_sc_hd__xnor2_1 _08319_ (.A(net171),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__or3_1 _08320_ (.A(net123),
    .B(_01414_),
    .C(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__a22o_1 _08321_ (.A1(_06494_),
    .A2(net118),
    .B1(_00352_),
    .B2(net292),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_4 _08322_ (.A(net240),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__o22a_1 _08323_ (.A1(net152),
    .A2(net114),
    .B1(net108),
    .B2(net154),
    .X(_01420_));
 sky130_fd_sc_hd__xnor2_1 _08324_ (.A(net195),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__or2_1 _08325_ (.A(_01419_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__o22a_1 _08326_ (.A1(net150),
    .A2(net116),
    .B1(net110),
    .B2(net148),
    .X(_01423_));
 sky130_fd_sc_hd__xnor2_1 _08327_ (.A(net191),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__xnor2_1 _08328_ (.A(_01419_),
    .B(_01421_),
    .Y(_01425_));
 sky130_fd_sc_hd__o21a_2 _08329_ (.A1(_01424_),
    .A2(_01425_),
    .B1(_01422_),
    .X(_01426_));
 sky130_fd_sc_hd__o21ai_1 _08330_ (.A1(_01414_),
    .A2(_01416_),
    .B1(net123),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _08331_ (.A(_01417_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__o21ai_2 _08332_ (.A1(_01426_),
    .A2(_01428_),
    .B1(_01417_),
    .Y(_01429_));
 sky130_fd_sc_hd__xnor2_2 _08333_ (.A(_01392_),
    .B(_01393_),
    .Y(_01430_));
 sky130_fd_sc_hd__and2b_1 _08334_ (.A_N(_01430_),
    .B(_01429_),
    .X(_01431_));
 sky130_fd_sc_hd__xor2_2 _08335_ (.A(_01379_),
    .B(_01381_),
    .X(_01432_));
 sky130_fd_sc_hd__xnor2_1 _08336_ (.A(_01370_),
    .B(_01372_),
    .Y(_01433_));
 sky130_fd_sc_hd__xnor2_1 _08337_ (.A(_01432_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__xnor2_1 _08338_ (.A(_01388_),
    .B(_01390_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2b_1 _08339_ (.A_N(_01434_),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__a21bo_1 _08340_ (.A1(_01432_),
    .A2(_01433_),
    .B1_N(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__xor2_2 _08341_ (.A(_01429_),
    .B(_01430_),
    .X(_01438_));
 sky130_fd_sc_hd__and2b_1 _08342_ (.A_N(_01438_),
    .B(_01437_),
    .X(_01439_));
 sky130_fd_sc_hd__or2_1 _08343_ (.A(_01431_),
    .B(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__xor2_2 _08344_ (.A(_01410_),
    .B(_01411_),
    .X(_01441_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(_01440_),
    .B(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__xnor2_1 _08346_ (.A(_01404_),
    .B(_01405_),
    .Y(_01443_));
 sky130_fd_sc_hd__a21oi_2 _08347_ (.A1(_01412_),
    .A2(_01442_),
    .B1(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__inv_2 _08348_ (.A(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__a21o_1 _08349_ (.A1(_01408_),
    .A2(_01445_),
    .B1(_01407_),
    .X(_01446_));
 sky130_fd_sc_hd__xnor2_2 _08350_ (.A(_01398_),
    .B(_01399_),
    .Y(_01447_));
 sky130_fd_sc_hd__xnor2_2 _08351_ (.A(_01437_),
    .B(_01438_),
    .Y(_01448_));
 sky130_fd_sc_hd__and2_1 _08352_ (.A(_01447_),
    .B(_01448_),
    .X(_01449_));
 sky130_fd_sc_hd__xor2_2 _08353_ (.A(_01426_),
    .B(_01428_),
    .X(_01450_));
 sky130_fd_sc_hd__o22a_1 _08354_ (.A1(net287),
    .A2(net119),
    .B1(net116),
    .B2(net237),
    .X(_01451_));
 sky130_fd_sc_hd__xnor2_1 _08355_ (.A(net238),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__o22a_1 _08356_ (.A1(net154),
    .A2(net114),
    .B1(net113),
    .B2(net152),
    .X(_01453_));
 sky130_fd_sc_hd__xnor2_1 _08357_ (.A(net195),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__or2_1 _08358_ (.A(_01452_),
    .B(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__o22a_1 _08359_ (.A1(net150),
    .A2(net110),
    .B1(net108),
    .B2(net148),
    .X(_01456_));
 sky130_fd_sc_hd__xnor2_2 _08360_ (.A(net191),
    .B(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__xnor2_1 _08361_ (.A(_01452_),
    .B(_01454_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _08362_ (.A(_01457_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__o21ai_2 _08363_ (.A1(_01457_),
    .A2(_01458_),
    .B1(_01455_),
    .Y(_01460_));
 sky130_fd_sc_hd__o22a_1 _08364_ (.A1(net141),
    .A2(net106),
    .B1(net104),
    .B2(net140),
    .X(_01461_));
 sky130_fd_sc_hd__xnor2_2 _08365_ (.A(_00328_),
    .B(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _08366_ (.A(_01460_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__o22a_1 _08367_ (.A1(net142),
    .A2(net86),
    .B1(net82),
    .B2(net209),
    .X(_01464_));
 sky130_fd_sc_hd__xnor2_2 _08368_ (.A(net138),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _08369_ (.A(_01460_),
    .B(_01462_),
    .Y(_01466_));
 sky130_fd_sc_hd__xor2_1 _08370_ (.A(_01460_),
    .B(_01462_),
    .X(_01467_));
 sky130_fd_sc_hd__o21a_1 _08371_ (.A1(_01465_),
    .A2(_01466_),
    .B1(_01463_),
    .X(_01468_));
 sky130_fd_sc_hd__and2b_1 _08372_ (.A_N(_01468_),
    .B(_01450_),
    .X(_01469_));
 sky130_fd_sc_hd__o22a_1 _08373_ (.A1(net144),
    .A2(net129),
    .B1(net107),
    .B2(net146),
    .X(_01470_));
 sky130_fd_sc_hd__xnor2_1 _08374_ (.A(net188),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__o22a_1 _08375_ (.A1(net133),
    .A2(net127),
    .B1(net141),
    .B2(net131),
    .X(_01472_));
 sky130_fd_sc_hd__xnor2_1 _08376_ (.A(net171),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__or2_1 _08377_ (.A(_01471_),
    .B(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__xnor2_1 _08378_ (.A(_01414_),
    .B(_01416_),
    .Y(_01475_));
 sky130_fd_sc_hd__or2_1 _08379_ (.A(_01474_),
    .B(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__xnor2_1 _08380_ (.A(_01424_),
    .B(_01425_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(_01474_),
    .B(_01475_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _08382_ (.A(_01476_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__or2_1 _08383_ (.A(_01477_),
    .B(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(_01476_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__xnor2_2 _08385_ (.A(_01450_),
    .B(_01468_),
    .Y(_01482_));
 sky130_fd_sc_hd__a21o_1 _08386_ (.A1(_01481_),
    .A2(_01482_),
    .B1(_01469_),
    .X(_01483_));
 sky130_fd_sc_hd__xor2_2 _08387_ (.A(_01447_),
    .B(_01448_),
    .X(_01484_));
 sky130_fd_sc_hd__a21oi_2 _08388_ (.A1(_01483_),
    .A2(_01484_),
    .B1(_01449_),
    .Y(_01485_));
 sky130_fd_sc_hd__xnor2_2 _08389_ (.A(_01440_),
    .B(_01441_),
    .Y(_01486_));
 sky130_fd_sc_hd__and2_1 _08390_ (.A(_01485_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__or2_1 _08391_ (.A(_01485_),
    .B(_01486_),
    .X(_01488_));
 sky130_fd_sc_hd__xnor2_1 _08392_ (.A(_01434_),
    .B(_01435_),
    .Y(_01489_));
 sky130_fd_sc_hd__inv_2 _08393_ (.A(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__xnor2_2 _08394_ (.A(_01481_),
    .B(_01482_),
    .Y(_01491_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(_01490_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__xnor2_2 _08396_ (.A(_01490_),
    .B(_01491_),
    .Y(_01493_));
 sky130_fd_sc_hd__xnor2_2 _08397_ (.A(_01465_),
    .B(_01467_),
    .Y(_01494_));
 sky130_fd_sc_hd__o22a_1 _08398_ (.A1(net140),
    .A2(net106),
    .B1(net104),
    .B2(net142),
    .X(_01495_));
 sky130_fd_sc_hd__xnor2_1 _08399_ (.A(net136),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__nor2_1 _08400_ (.A(net209),
    .B(net86),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_1 _08401_ (.A(_01496_),
    .B(_01497_),
    .Y(_01498_));
 sky130_fd_sc_hd__o21a_1 _08402_ (.A1(_00324_),
    .A2(_01497_),
    .B1(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__nand2_1 _08403_ (.A(_01494_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__o22a_1 _08404_ (.A1(net287),
    .A2(net116),
    .B1(net110),
    .B2(net237),
    .X(_01501_));
 sky130_fd_sc_hd__xnor2_1 _08405_ (.A(net238),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__o22a_1 _08406_ (.A1(net148),
    .A2(net114),
    .B1(net108),
    .B2(net150),
    .X(_01503_));
 sky130_fd_sc_hd__xnor2_1 _08407_ (.A(net191),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__or2_1 _08408_ (.A(_01502_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__nand2_1 _08409_ (.A(_01471_),
    .B(_01473_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(_01474_),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__or2_1 _08411_ (.A(_01505_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__xnor2_1 _08412_ (.A(_01505_),
    .B(_01507_),
    .Y(_01509_));
 sky130_fd_sc_hd__and2_1 _08413_ (.A(_01457_),
    .B(_01458_),
    .X(_01510_));
 sky130_fd_sc_hd__nor2_1 _08414_ (.A(_01459_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__o31a_1 _08415_ (.A1(_01459_),
    .A2(_01509_),
    .A3(_01510_),
    .B1(_01508_),
    .X(_01512_));
 sky130_fd_sc_hd__xnor2_2 _08416_ (.A(_01494_),
    .B(_01499_),
    .Y(_01513_));
 sky130_fd_sc_hd__o21a_1 _08417_ (.A1(_01512_),
    .A2(_01513_),
    .B1(_01500_),
    .X(_01514_));
 sky130_fd_sc_hd__nor2_1 _08418_ (.A(_01493_),
    .B(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _08419_ (.A(_01492_),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__xor2_2 _08420_ (.A(_01483_),
    .B(_01484_),
    .X(_01517_));
 sky130_fd_sc_hd__nand2b_1 _08421_ (.A_N(_01516_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21o_1 _08422_ (.A1(_01488_),
    .A2(_01518_),
    .B1(_01487_),
    .X(_01519_));
 sky130_fd_sc_hd__xnor2_2 _08423_ (.A(_01485_),
    .B(_01486_),
    .Y(_01520_));
 sky130_fd_sc_hd__or3_1 _08424_ (.A(_01492_),
    .B(_01515_),
    .C(_01517_),
    .X(_01521_));
 sky130_fd_sc_hd__xnor2_2 _08425_ (.A(_01516_),
    .B(_01517_),
    .Y(_01522_));
 sky130_fd_sc_hd__xnor2_2 _08426_ (.A(_01493_),
    .B(_01514_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _08427_ (.A(_01477_),
    .B(_01479_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(_01480_),
    .B(_01524_),
    .Y(_01525_));
 sky130_fd_sc_hd__xnor2_2 _08429_ (.A(_01512_),
    .B(_01513_),
    .Y(_01526_));
 sky130_fd_sc_hd__or2_1 _08430_ (.A(_01525_),
    .B(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__o22a_1 _08431_ (.A1(net133),
    .A2(net141),
    .B1(net140),
    .B2(net131),
    .X(_01528_));
 sky130_fd_sc_hd__xnor2_1 _08432_ (.A(net171),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__o22a_1 _08433_ (.A1(net154),
    .A2(net113),
    .B1(net107),
    .B2(net152),
    .X(_01530_));
 sky130_fd_sc_hd__xnor2_1 _08434_ (.A(net195),
    .B(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__or2_1 _08435_ (.A(_01529_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__o22a_1 _08436_ (.A1(net146),
    .A2(net129),
    .B1(net127),
    .B2(net144),
    .X(_01533_));
 sky130_fd_sc_hd__xnor2_1 _08437_ (.A(net188),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__xnor2_1 _08438_ (.A(_01529_),
    .B(_01531_),
    .Y(_01535_));
 sky130_fd_sc_hd__o21a_1 _08439_ (.A1(_01534_),
    .A2(_01535_),
    .B1(_01532_),
    .X(_01536_));
 sky130_fd_sc_hd__or2_1 _08440_ (.A(_01496_),
    .B(_01497_),
    .X(_01537_));
 sky130_fd_sc_hd__nand2_1 _08441_ (.A(_01498_),
    .B(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand2b_1 _08442_ (.A_N(_01536_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__xnor2_1 _08443_ (.A(_01502_),
    .B(_01504_),
    .Y(_01540_));
 sky130_fd_sc_hd__o22a_1 _08444_ (.A1(net142),
    .A2(net106),
    .B1(net104),
    .B2(net209),
    .X(_01541_));
 sky130_fd_sc_hd__xnor2_1 _08445_ (.A(net136),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__o22a_1 _08446_ (.A1(net150),
    .A2(net114),
    .B1(net113),
    .B2(net148),
    .X(_01543_));
 sky130_fd_sc_hd__xnor2_1 _08447_ (.A(net191),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__o22a_1 _08448_ (.A1(net287),
    .A2(net110),
    .B1(net108),
    .B2(net237),
    .X(_01545_));
 sky130_fd_sc_hd__xnor2_2 _08449_ (.A(net238),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__or2_1 _08450_ (.A(_01544_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__xnor2_1 _08451_ (.A(_01540_),
    .B(_01542_),
    .Y(_01548_));
 sky130_fd_sc_hd__o32a_1 _08452_ (.A1(_01544_),
    .A2(_01546_),
    .A3(_01548_),
    .B1(_01542_),
    .B2(_01540_),
    .X(_01549_));
 sky130_fd_sc_hd__xnor2_1 _08453_ (.A(_01536_),
    .B(_01538_),
    .Y(_01550_));
 sky130_fd_sc_hd__nand2b_1 _08454_ (.A_N(_01549_),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _08455_ (.A(_01539_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__xor2_2 _08456_ (.A(_01525_),
    .B(_01526_),
    .X(_01553_));
 sky130_fd_sc_hd__nand2_1 _08457_ (.A(_01552_),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__and3_1 _08458_ (.A(_01523_),
    .B(_01527_),
    .C(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__nand3_2 _08459_ (.A(_01523_),
    .B(_01527_),
    .C(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__xnor2_1 _08460_ (.A(_01509_),
    .B(_01511_),
    .Y(_01557_));
 sky130_fd_sc_hd__xnor2_1 _08461_ (.A(_01549_),
    .B(_01550_),
    .Y(_01558_));
 sky130_fd_sc_hd__xnor2_1 _08462_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__xor2_1 _08463_ (.A(_01534_),
    .B(_01535_),
    .X(_01560_));
 sky130_fd_sc_hd__o22a_1 _08464_ (.A1(net131),
    .A2(net142),
    .B1(net140),
    .B2(net133),
    .X(_01561_));
 sky130_fd_sc_hd__xnor2_1 _08465_ (.A(net171),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__o22a_1 _08466_ (.A1(net152),
    .A2(net129),
    .B1(net107),
    .B2(net154),
    .X(_01563_));
 sky130_fd_sc_hd__xnor2_1 _08467_ (.A(net195),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__or2_1 _08468_ (.A(_01562_),
    .B(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__o22a_1 _08469_ (.A1(net146),
    .A2(net127),
    .B1(net141),
    .B2(net144),
    .X(_01566_));
 sky130_fd_sc_hd__xor2_1 _08470_ (.A(net188),
    .B(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__inv_2 _08471_ (.A(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__xnor2_1 _08472_ (.A(_01562_),
    .B(_01564_),
    .Y(_01569_));
 sky130_fd_sc_hd__o21a_1 _08473_ (.A1(_01568_),
    .A2(_01569_),
    .B1(_01565_),
    .X(_01570_));
 sky130_fd_sc_hd__nand2b_1 _08474_ (.A_N(_01570_),
    .B(_01560_),
    .Y(_01571_));
 sky130_fd_sc_hd__xnor2_1 _08475_ (.A(_01560_),
    .B(_01570_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_2 _08476_ (.A(net208),
    .B(_00378_),
    .Y(_01573_));
 sky130_fd_sc_hd__xor2_1 _08477_ (.A(_01544_),
    .B(_01546_),
    .X(_01574_));
 sky130_fd_sc_hd__nor2_1 _08478_ (.A(_01573_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__a21oi_1 _08479_ (.A1(net136),
    .A2(_01573_),
    .B1(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__a21bo_1 _08480_ (.A1(_01572_),
    .A2(_01576_),
    .B1_N(_01571_),
    .X(_01577_));
 sky130_fd_sc_hd__nand2b_1 _08481_ (.A_N(_01559_),
    .B(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hd__a21bo_1 _08482_ (.A1(_01557_),
    .A2(_01558_),
    .B1_N(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__xor2_2 _08483_ (.A(_01552_),
    .B(_01553_),
    .X(_01580_));
 sky130_fd_sc_hd__and2_1 _08484_ (.A(_01579_),
    .B(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__a21oi_2 _08485_ (.A1(_01527_),
    .A2(_01554_),
    .B1(_01523_),
    .Y(_01582_));
 sky130_fd_sc_hd__inv_2 _08486_ (.A(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__or2_1 _08487_ (.A(_01579_),
    .B(_01580_),
    .X(_01584_));
 sky130_fd_sc_hd__xor2_2 _08488_ (.A(_01579_),
    .B(_01580_),
    .X(_01585_));
 sky130_fd_sc_hd__xor2_1 _08489_ (.A(_01559_),
    .B(_01577_),
    .X(_01586_));
 sky130_fd_sc_hd__xnor2_1 _08490_ (.A(_01547_),
    .B(_01548_),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_1 _08491_ (.A(_01572_),
    .B(_01576_),
    .Y(_01588_));
 sky130_fd_sc_hd__or2_1 _08492_ (.A(_01587_),
    .B(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__xnor2_1 _08493_ (.A(_01587_),
    .B(_01588_),
    .Y(_01590_));
 sky130_fd_sc_hd__o22a_1 _08494_ (.A1(net237),
    .A2(net114),
    .B1(net108),
    .B2(net287),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08495_ (.A(net238),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__o22a_1 _08496_ (.A1(net154),
    .A2(net129),
    .B1(net127),
    .B2(net152),
    .X(_01593_));
 sky130_fd_sc_hd__xnor2_1 _08497_ (.A(net195),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__or2_1 _08498_ (.A(_01592_),
    .B(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_1 _08499_ (.A(_01592_),
    .B(_01594_),
    .Y(_01596_));
 sky130_fd_sc_hd__a22o_1 _08500_ (.A1(_06532_),
    .A2(net112),
    .B1(_00360_),
    .B2(_06540_),
    .X(_01597_));
 sky130_fd_sc_hd__xnor2_2 _08501_ (.A(net191),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__inv_2 _08502_ (.A(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__o21a_1 _08503_ (.A1(_01596_),
    .A2(_01599_),
    .B1(_01595_),
    .X(_01600_));
 sky130_fd_sc_hd__xnor2_1 _08504_ (.A(_01568_),
    .B(_01569_),
    .Y(_01601_));
 sky130_fd_sc_hd__o22a_1 _08505_ (.A1(net146),
    .A2(net141),
    .B1(net140),
    .B2(net144),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_1 _08506_ (.A(net188),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__o22a_1 _08507_ (.A1(net209),
    .A2(net131),
    .B1(net142),
    .B2(net133),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _08508_ (.A(net171),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _08509_ (.A(_01603_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__xor2_1 _08510_ (.A(_01600_),
    .B(_01601_),
    .X(_01607_));
 sky130_fd_sc_hd__nand2_1 _08511_ (.A(_01606_),
    .B(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__o21ai_1 _08512_ (.A1(_01600_),
    .A2(_01601_),
    .B1(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2b_1 _08513_ (.A_N(_01590_),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__and3_1 _08514_ (.A(_01586_),
    .B(_01589_),
    .C(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__xnor2_1 _08515_ (.A(_01590_),
    .B(_01609_),
    .Y(_01612_));
 sky130_fd_sc_hd__xnor2_1 _08516_ (.A(_01606_),
    .B(_01607_),
    .Y(_01613_));
 sky130_fd_sc_hd__and2_1 _08517_ (.A(_01573_),
    .B(_01574_),
    .X(_01614_));
 sky130_fd_sc_hd__nor2_1 _08518_ (.A(_01575_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _08519_ (.A(_01613_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__xnor2_1 _08520_ (.A(_01596_),
    .B(_01598_),
    .Y(_01617_));
 sky130_fd_sc_hd__o22a_1 _08521_ (.A1(net287),
    .A2(net114),
    .B1(net113),
    .B2(net237),
    .X(_01618_));
 sky130_fd_sc_hd__xnor2_2 _08522_ (.A(net238),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__o22a_1 _08523_ (.A1(net154),
    .A2(net127),
    .B1(net141),
    .B2(net152),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_2 _08524_ (.A(net195),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__or2_1 _08525_ (.A(_01619_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__o22a_1 _08526_ (.A1(net148),
    .A2(net129),
    .B1(net107),
    .B2(net150),
    .X(_01623_));
 sky130_fd_sc_hd__xnor2_2 _08527_ (.A(net191),
    .B(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__xnor2_2 _08528_ (.A(_01619_),
    .B(_01621_),
    .Y(_01625_));
 sky130_fd_sc_hd__o21a_1 _08529_ (.A1(_01624_),
    .A2(_01625_),
    .B1(_01622_),
    .X(_01626_));
 sky130_fd_sc_hd__nand2b_1 _08530_ (.A_N(_01626_),
    .B(_01617_),
    .Y(_01627_));
 sky130_fd_sc_hd__o22a_1 _08531_ (.A1(net144),
    .A2(net142),
    .B1(net140),
    .B2(net146),
    .X(_01628_));
 sky130_fd_sc_hd__xnor2_2 _08532_ (.A(net188),
    .B(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__nor2_1 _08533_ (.A(net209),
    .B(net133),
    .Y(_01630_));
 sky130_fd_sc_hd__xnor2_2 _08534_ (.A(net171),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__and2b_1 _08535_ (.A_N(_01629_),
    .B(_01631_),
    .X(_01632_));
 sky130_fd_sc_hd__xnor2_1 _08536_ (.A(_01617_),
    .B(_01626_),
    .Y(_01633_));
 sky130_fd_sc_hd__a21bo_1 _08537_ (.A1(_01632_),
    .A2(_01633_),
    .B1_N(_01627_),
    .X(_01634_));
 sky130_fd_sc_hd__xnor2_1 _08538_ (.A(_01613_),
    .B(_01615_),
    .Y(_01635_));
 sky130_fd_sc_hd__and2b_1 _08539_ (.A_N(_01635_),
    .B(_01634_),
    .X(_01636_));
 sky130_fd_sc_hd__o21a_1 _08540_ (.A1(_01616_),
    .A2(_01636_),
    .B1(_01612_),
    .X(_01637_));
 sky130_fd_sc_hd__a21oi_2 _08541_ (.A1(_01589_),
    .A2(_01610_),
    .B1(_01586_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor3_1 _08542_ (.A(_01612_),
    .B(_01616_),
    .C(_01636_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_01637_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__and2_1 _08544_ (.A(_01603_),
    .B(_01605_),
    .X(_01641_));
 sky130_fd_sc_hd__or2_1 _08545_ (.A(_01606_),
    .B(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__xnor2_1 _08546_ (.A(_01632_),
    .B(_01633_),
    .Y(_01643_));
 sky130_fd_sc_hd__or2_1 _08547_ (.A(_01642_),
    .B(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__xor2_1 _08548_ (.A(_01642_),
    .B(_01643_),
    .X(_01645_));
 sky130_fd_sc_hd__xor2_2 _08549_ (.A(_01624_),
    .B(_01625_),
    .X(_01646_));
 sky130_fd_sc_hd__and2b_1 _08550_ (.A_N(net171),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__o22a_1 _08551_ (.A1(net287),
    .A2(net113),
    .B1(net107),
    .B2(net237),
    .X(_01648_));
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(net238),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__o22a_1 _08553_ (.A1(net150),
    .A2(net129),
    .B1(net127),
    .B2(net148),
    .X(_01650_));
 sky130_fd_sc_hd__xnor2_1 _08554_ (.A(net191),
    .B(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__nor2_2 _08555_ (.A(_01649_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__xnor2_2 _08556_ (.A(net171),
    .B(_01646_),
    .Y(_01653_));
 sky130_fd_sc_hd__a21o_1 _08557_ (.A1(_01652_),
    .A2(_01653_),
    .B1(_01647_),
    .X(_01654_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_01645_),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__xor2_1 _08559_ (.A(_01634_),
    .B(_01635_),
    .X(_01656_));
 sky130_fd_sc_hd__and3_1 _08560_ (.A(_01644_),
    .B(_01655_),
    .C(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__nand3_1 _08561_ (.A(_01644_),
    .B(_01655_),
    .C(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__xnor2_2 _08562_ (.A(_01629_),
    .B(_01631_),
    .Y(_01659_));
 sky130_fd_sc_hd__xor2_2 _08563_ (.A(_01652_),
    .B(_01653_),
    .X(_01660_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(_01659_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__a22o_1 _08565_ (.A1(_06494_),
    .A2(_00198_),
    .B1(_00360_),
    .B2(net292),
    .X(_01662_));
 sky130_fd_sc_hd__xnor2_2 _08566_ (.A(net238),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a22o_1 _08567_ (.A1(_06532_),
    .A2(_00211_),
    .B1(_00243_),
    .B2(_06540_),
    .X(_01664_));
 sky130_fd_sc_hd__xnor2_2 _08568_ (.A(net193),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__o22a_1 _08569_ (.A1(net154),
    .A2(net141),
    .B1(net140),
    .B2(net152),
    .X(_01666_));
 sky130_fd_sc_hd__xnor2_1 _08570_ (.A(_06507_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand3_2 _08571_ (.A(_01663_),
    .B(_01665_),
    .C(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__o22a_1 _08572_ (.A1(net209),
    .A2(net144),
    .B1(net142),
    .B2(net147),
    .X(_01669_));
 sky130_fd_sc_hd__xor2_1 _08573_ (.A(net188),
    .B(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__a21o_1 _08574_ (.A1(_01663_),
    .A2(_01665_),
    .B1(_01667_),
    .X(_01671_));
 sky130_fd_sc_hd__nand3_2 _08575_ (.A(_01668_),
    .B(_01670_),
    .C(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_2 _08576_ (.A(_01668_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__inv_2 _08577_ (.A(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__xnor2_2 _08578_ (.A(_01659_),
    .B(_01660_),
    .Y(_01675_));
 sky130_fd_sc_hd__o21ai_2 _08579_ (.A1(_01674_),
    .A2(_01675_),
    .B1(_01661_),
    .Y(_01676_));
 sky130_fd_sc_hd__xor2_1 _08580_ (.A(_01645_),
    .B(_01654_),
    .X(_01677_));
 sky130_fd_sc_hd__and2_1 _08581_ (.A(_01676_),
    .B(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__a21oi_1 _08582_ (.A1(_01644_),
    .A2(_01655_),
    .B1(_01656_),
    .Y(_01679_));
 sky130_fd_sc_hd__or2_1 _08583_ (.A(_01676_),
    .B(_01677_),
    .X(_01680_));
 sky130_fd_sc_hd__xor2_1 _08584_ (.A(_01676_),
    .B(_01677_),
    .X(_01681_));
 sky130_fd_sc_hd__and2_1 _08585_ (.A(_01649_),
    .B(_01651_),
    .X(_01682_));
 sky130_fd_sc_hd__nor2_1 _08586_ (.A(_01652_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__a21o_1 _08587_ (.A1(_01668_),
    .A2(_01671_),
    .B1(_01670_),
    .X(_01684_));
 sky130_fd_sc_hd__nand3_1 _08588_ (.A(_01672_),
    .B(_01683_),
    .C(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21o_1 _08589_ (.A1(_01672_),
    .A2(_01684_),
    .B1(_01683_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_1 _08590_ (.A(net210),
    .B(net147),
    .Y(_01687_));
 sky130_fd_sc_hd__o22a_1 _08591_ (.A1(net152),
    .A2(net142),
    .B1(net140),
    .B2(net154),
    .X(_01688_));
 sky130_fd_sc_hd__xnor2_1 _08592_ (.A(net195),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _08593_ (.A(_01687_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__o21ai_1 _08594_ (.A1(net210),
    .A2(net146),
    .B1(_00140_),
    .Y(_01691_));
 sky130_fd_sc_hd__and4_1 _08595_ (.A(_01685_),
    .B(_01686_),
    .C(_01690_),
    .D(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__a31o_2 _08596_ (.A1(_01672_),
    .A2(_01683_),
    .A3(_01684_),
    .B1(_01692_),
    .X(_01693_));
 sky130_fd_sc_hd__xnor2_2 _08597_ (.A(_01673_),
    .B(_01675_),
    .Y(_01694_));
 sky130_fd_sc_hd__or2_1 _08598_ (.A(_01693_),
    .B(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__and2_1 _08599_ (.A(_01693_),
    .B(_01694_),
    .X(_01696_));
 sky130_fd_sc_hd__xor2_1 _08600_ (.A(_01663_),
    .B(_01665_),
    .X(_01697_));
 sky130_fd_sc_hd__or2_1 _08601_ (.A(_01687_),
    .B(_01689_),
    .X(_01698_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_01690_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _08603_ (.A(_01697_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__a21oi_1 _08604_ (.A1(_00195_),
    .A2(_00196_),
    .B1(net288),
    .Y(_01701_));
 sky130_fd_sc_hd__and3_1 _08605_ (.A(_06494_),
    .B(_00209_),
    .C(_00210_),
    .X(_01702_));
 sky130_fd_sc_hd__o21ai_1 _08606_ (.A1(_01701_),
    .A2(_01702_),
    .B1(net240),
    .Y(_01703_));
 sky130_fd_sc_hd__or3_1 _08607_ (.A(net240),
    .B(_01701_),
    .C(_01702_),
    .X(_01704_));
 sky130_fd_sc_hd__a22o_1 _08608_ (.A1(_06532_),
    .A2(_00243_),
    .B1(_00250_),
    .B2(_06540_),
    .X(_01705_));
 sky130_fd_sc_hd__xnor2_1 _08609_ (.A(net192),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__and3_2 _08610_ (.A(_01703_),
    .B(_01704_),
    .C(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__xor2_1 _08611_ (.A(_01697_),
    .B(_01699_),
    .X(_01708_));
 sky130_fd_sc_hd__nand2_1 _08612_ (.A(_01707_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__a22oi_2 _08613_ (.A1(_01685_),
    .A2(_01686_),
    .B1(_01690_),
    .B2(_01691_),
    .Y(_01710_));
 sky130_fd_sc_hd__a211oi_1 _08614_ (.A1(_01700_),
    .A2(_01709_),
    .B1(_01710_),
    .C1(_01692_),
    .Y(_01711_));
 sky130_fd_sc_hd__o211a_1 _08615_ (.A1(_01692_),
    .A2(_01710_),
    .B1(_01709_),
    .C1(_01700_),
    .X(_01712_));
 sky130_fd_sc_hd__nor2_1 _08616_ (.A(_01711_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__xnor2_1 _08617_ (.A(_01707_),
    .B(_01708_),
    .Y(_01714_));
 sky130_fd_sc_hd__a21oi_1 _08618_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_01706_),
    .Y(_01715_));
 sky130_fd_sc_hd__o22a_1 _08619_ (.A1(net210),
    .A2(net152),
    .B1(net142),
    .B2(net154),
    .X(_01716_));
 sky130_fd_sc_hd__xnor2_1 _08620_ (.A(_06507_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__nor3b_1 _08621_ (.A(_01707_),
    .B(_01715_),
    .C_N(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__or3b_1 _08622_ (.A(_01707_),
    .B(_01715_),
    .C_N(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__a22o_1 _08623_ (.A1(_06540_),
    .A2(_00225_),
    .B1(_00250_),
    .B2(_06532_),
    .X(_01720_));
 sky130_fd_sc_hd__xor2_1 _08624_ (.A(net191),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__a32o_1 _08625_ (.A1(net292),
    .A2(_00209_),
    .A3(_00210_),
    .B1(_00243_),
    .B2(_06494_),
    .X(_01722_));
 sky130_fd_sc_hd__xnor2_1 _08626_ (.A(net240),
    .B(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__or2_1 _08627_ (.A(_01721_),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__o21ba_1 _08628_ (.A1(_01707_),
    .A2(_01715_),
    .B1_N(_01717_),
    .X(_01725_));
 sky130_fd_sc_hd__or3_2 _08629_ (.A(_01718_),
    .B(_01724_),
    .C(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__and3_1 _08630_ (.A(_01714_),
    .B(_01719_),
    .C(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__a21oi_1 _08631_ (.A1(_01719_),
    .A2(_01726_),
    .B1(_01714_),
    .Y(_01728_));
 sky130_fd_sc_hd__xor2_1 _08632_ (.A(_01721_),
    .B(_01723_),
    .X(_01729_));
 sky130_fd_sc_hd__nor2_1 _08633_ (.A(net210),
    .B(net155),
    .Y(_01730_));
 sky130_fd_sc_hd__mux2_1 _08634_ (.A0(_06507_),
    .A1(_01729_),
    .S(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__o21ai_1 _08635_ (.A1(_01718_),
    .A2(_01725_),
    .B1(_01724_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21oi_1 _08636_ (.A1(_01726_),
    .A2(_01732_),
    .B1(_01731_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21o_1 _08637_ (.A1(_01726_),
    .A2(_01732_),
    .B1(_01731_),
    .X(_01734_));
 sky130_fd_sc_hd__and3_1 _08638_ (.A(_01726_),
    .B(_01731_),
    .C(_01732_),
    .X(_01735_));
 sky130_fd_sc_hd__a22o_1 _08639_ (.A1(net292),
    .A2(_00243_),
    .B1(_00250_),
    .B2(_06494_),
    .X(_01736_));
 sky130_fd_sc_hd__xnor2_1 _08640_ (.A(net240),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__o22a_1 _08641_ (.A1(net209),
    .A2(net148),
    .B1(net143),
    .B2(net150),
    .X(_01738_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(net193),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _08643_ (.A(_01737_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__xnor2_1 _08644_ (.A(_01729_),
    .B(_01730_),
    .Y(_01741_));
 sky130_fd_sc_hd__and2b_1 _08645_ (.A_N(_01741_),
    .B(_01740_),
    .X(_01742_));
 sky130_fd_sc_hd__xnor2_1 _08646_ (.A(_01740_),
    .B(_01741_),
    .Y(_01743_));
 sky130_fd_sc_hd__a22o_1 _08647_ (.A1(_06494_),
    .A2(_00225_),
    .B1(_00250_),
    .B2(net292),
    .X(_01744_));
 sky130_fd_sc_hd__xnor2_2 _08648_ (.A(net240),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _08649_ (.A(net209),
    .B(net150),
    .Y(_01746_));
 sky130_fd_sc_hd__xnor2_1 _08650_ (.A(net193),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__and2b_1 _08651_ (.A_N(_01745_),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__and2b_1 _08652_ (.A_N(_01747_),
    .B(_01745_),
    .X(_01749_));
 sky130_fd_sc_hd__xor2_1 _08653_ (.A(_01745_),
    .B(_01746_),
    .X(_01750_));
 sky130_fd_sc_hd__a22o_1 _08654_ (.A1(net208),
    .A2(_06494_),
    .B1(_00225_),
    .B2(net292),
    .X(_01751_));
 sky130_fd_sc_hd__or2_1 _08655_ (.A(_06416_),
    .B(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__or3_1 _08656_ (.A(net239),
    .B(_01750_),
    .C(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__xor2_1 _08657_ (.A(_01737_),
    .B(_01739_),
    .X(_01754_));
 sky130_fd_sc_hd__xnor2_1 _08658_ (.A(_01748_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__mux2_1 _08659_ (.A0(net193),
    .A1(_01745_),
    .S(_01746_),
    .X(_01756_));
 sky130_fd_sc_hd__inv_2 _08660_ (.A(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__a2bb2o_1 _08661_ (.A1_N(_01753_),
    .A2_N(_01755_),
    .B1(_01757_),
    .B2(_01754_),
    .X(_01758_));
 sky130_fd_sc_hd__a21o_1 _08662_ (.A1(_01743_),
    .A2(_01758_),
    .B1(_01742_),
    .X(_01759_));
 sky130_fd_sc_hd__nor2_1 _08663_ (.A(_01733_),
    .B(_01735_),
    .Y(_01760_));
 sky130_fd_sc_hd__a21o_1 _08664_ (.A1(_01734_),
    .A2(_01759_),
    .B1(_01735_),
    .X(_01761_));
 sky130_fd_sc_hd__o21ba_1 _08665_ (.A1(_01728_),
    .A2(_01761_),
    .B1_N(_01727_),
    .X(_01762_));
 sky130_fd_sc_hd__or2_1 _08666_ (.A(_01727_),
    .B(_01728_),
    .X(_01763_));
 sky130_fd_sc_hd__o21ba_2 _08667_ (.A1(_01711_),
    .A2(_01762_),
    .B1_N(_01712_),
    .X(_01764_));
 sky130_fd_sc_hd__a21o_1 _08668_ (.A1(_01693_),
    .A2(_01694_),
    .B1(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__xor2_2 _08669_ (.A(_01693_),
    .B(_01694_),
    .X(_01766_));
 sky130_fd_sc_hd__and3_1 _08670_ (.A(_01681_),
    .B(_01695_),
    .C(_01765_),
    .X(_01767_));
 sky130_fd_sc_hd__a311o_1 _08671_ (.A1(_01681_),
    .A2(_01695_),
    .A3(_01765_),
    .B1(_01679_),
    .C1(_01678_),
    .X(_01768_));
 sky130_fd_sc_hd__nor2_1 _08672_ (.A(_01657_),
    .B(_01679_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand3_1 _08673_ (.A(_01640_),
    .B(_01658_),
    .C(_01768_),
    .Y(_01770_));
 sky130_fd_sc_hd__o21ba_1 _08674_ (.A1(_01637_),
    .A2(_01638_),
    .B1_N(_01611_),
    .X(_01771_));
 sky130_fd_sc_hd__nor2_2 _08675_ (.A(_01611_),
    .B(_01638_),
    .Y(_01772_));
 sky130_fd_sc_hd__a41o_1 _08676_ (.A1(_01640_),
    .A2(_01658_),
    .A3(_01768_),
    .A4(_01772_),
    .B1(_01771_),
    .X(_01773_));
 sky130_fd_sc_hd__a211o_1 _08677_ (.A1(_01585_),
    .A2(_01773_),
    .B1(_01581_),
    .C1(_01582_),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _08678_ (.A(_01555_),
    .B(_01582_),
    .Y(_01775_));
 sky130_fd_sc_hd__nand3_1 _08679_ (.A(_01522_),
    .B(_01556_),
    .C(_01774_),
    .Y(_01776_));
 sky130_fd_sc_hd__nand4b_2 _08680_ (.A_N(_01520_),
    .B(_01522_),
    .C(_01556_),
    .D(_01774_),
    .Y(_01777_));
 sky130_fd_sc_hd__and2_1 _08681_ (.A(_01519_),
    .B(_01777_),
    .X(_01778_));
 sky130_fd_sc_hd__xnor2_2 _08682_ (.A(_01364_),
    .B(_01406_),
    .Y(_01779_));
 sky130_fd_sc_hd__and3_1 _08683_ (.A(_01412_),
    .B(_01442_),
    .C(_01443_),
    .X(_01780_));
 sky130_fd_sc_hd__nor2_1 _08684_ (.A(_01444_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2_1 _08685_ (.A(_01444_),
    .B(_01780_),
    .X(_01782_));
 sky130_fd_sc_hd__a211o_1 _08686_ (.A1(_01519_),
    .A2(_01777_),
    .B1(_01779_),
    .C1(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__or4_1 _08687_ (.A(_01359_),
    .B(_01362_),
    .C(_01779_),
    .D(_01782_),
    .X(_01784_));
 sky130_fd_sc_hd__o221a_1 _08688_ (.A1(_01363_),
    .A2(_01446_),
    .B1(_01778_),
    .B2(_01784_),
    .C1(_01358_),
    .X(_01785_));
 sky130_fd_sc_hd__a22o_1 _08689_ (.A1(_01091_),
    .A2(_01092_),
    .B1(_01155_),
    .B2(_01156_),
    .X(_01786_));
 sky130_fd_sc_hd__o21ai_1 _08690_ (.A1(_01091_),
    .A2(_01092_),
    .B1(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__a21o_1 _08691_ (.A1(_01258_),
    .A2(_01262_),
    .B1(_01263_),
    .X(_01788_));
 sky130_fd_sc_hd__a2111o_1 _08692_ (.A1(_01258_),
    .A2(_01262_),
    .B1(_01263_),
    .C1(_01157_),
    .D1(_01094_),
    .X(_01789_));
 sky130_fd_sc_hd__o311a_2 _08693_ (.A1(_01158_),
    .A2(_01265_),
    .A3(_01785_),
    .B1(_01787_),
    .C1(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__a21o_1 _08694_ (.A1(_00902_),
    .A2(_00956_),
    .B1(_00957_),
    .X(_01791_));
 sky130_fd_sc_hd__a21o_1 _08695_ (.A1(_01030_),
    .A2(_01791_),
    .B1(_00958_),
    .X(_01792_));
 sky130_fd_sc_hd__nand2b_4 _08696_ (.A_N(_00958_),
    .B(_01791_),
    .Y(_01793_));
 sky130_fd_sc_hd__o31ai_4 _08697_ (.A1(_01031_),
    .A2(_01790_),
    .A3(_01793_),
    .B1(_01792_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _08698_ (.A(_00896_),
    .B(_00897_),
    .Y(_01795_));
 sky130_fd_sc_hd__xor2_2 _08699_ (.A(_00896_),
    .B(_00897_),
    .X(_01796_));
 sky130_fd_sc_hd__xnor2_1 _08700_ (.A(_00896_),
    .B(_00897_),
    .Y(_01797_));
 sky130_fd_sc_hd__xor2_1 _08701_ (.A(_00758_),
    .B(_00827_),
    .X(_01798_));
 sky130_fd_sc_hd__xnor2_1 _08702_ (.A(_00758_),
    .B(_00827_),
    .Y(_01799_));
 sky130_fd_sc_hd__a32o_2 _08703_ (.A1(_01794_),
    .A2(_01796_),
    .A3(_01798_),
    .B1(_00899_),
    .B2(_00828_),
    .X(_01800_));
 sky130_fd_sc_hd__xnor2_2 _08704_ (.A(_00757_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__xor2_2 _08705_ (.A(_01031_),
    .B(_01790_),
    .X(_01802_));
 sky130_fd_sc_hd__o21ai_1 _08706_ (.A1(net239),
    .A2(_01752_),
    .B1(_01750_),
    .Y(_01803_));
 sky130_fd_sc_hd__and2_1 _08707_ (.A(_01753_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_1 _08708_ (.A(_01752_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__o31ai_1 _08709_ (.A1(net191),
    .A2(_01748_),
    .A3(_01749_),
    .B1(_01753_),
    .Y(_01806_));
 sky130_fd_sc_hd__xor2_1 _08710_ (.A(_01755_),
    .B(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_01805_),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__xor2_1 _08712_ (.A(_01743_),
    .B(_01758_),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_1 _08713_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(_01759_),
    .B(_01760_),
    .Y(_01811_));
 sky130_fd_sc_hd__and2_1 _08715_ (.A(_01810_),
    .B(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__xor2_1 _08716_ (.A(_01761_),
    .B(_01763_),
    .X(_01813_));
 sky130_fd_sc_hd__and2_1 _08717_ (.A(_01812_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__xnor2_1 _08718_ (.A(_01713_),
    .B(_01762_),
    .Y(_01815_));
 sky130_fd_sc_hd__and2_1 _08719_ (.A(_01814_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_2 _08720_ (.A(_01764_),
    .B(_01766_),
    .Y(_01817_));
 sky130_fd_sc_hd__and2_1 _08721_ (.A(_01816_),
    .B(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__a21oi_1 _08722_ (.A1(_01695_),
    .A2(_01765_),
    .B1(_01681_),
    .Y(_01819_));
 sky130_fd_sc_hd__or2_1 _08723_ (.A(_01767_),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__o211ai_2 _08724_ (.A1(_01767_),
    .A2(_01819_),
    .B1(_01817_),
    .C1(_01816_),
    .Y(_01821_));
 sky130_fd_sc_hd__a211o_1 _08725_ (.A1(_01764_),
    .A2(_01766_),
    .B1(_01678_),
    .C1(_01696_),
    .X(_01822_));
 sky130_fd_sc_hd__nand3_1 _08726_ (.A(_01680_),
    .B(_01769_),
    .C(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__a21o_1 _08727_ (.A1(_01680_),
    .A2(_01822_),
    .B1(_01769_),
    .X(_01824_));
 sky130_fd_sc_hd__nand2_1 _08728_ (.A(_01823_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _08729_ (.A1(_01658_),
    .A2(_01768_),
    .B1(_01640_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _08730_ (.A(_01770_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a221o_1 _08731_ (.A1(_01823_),
    .A2(_01824_),
    .B1(_01826_),
    .B2(_01770_),
    .C1(_01821_),
    .X(_01828_));
 sky130_fd_sc_hd__o21ba_1 _08732_ (.A1(_01637_),
    .A2(_01679_),
    .B1_N(_01639_),
    .X(_01829_));
 sky130_fd_sc_hd__a41o_1 _08733_ (.A1(_01640_),
    .A2(_01680_),
    .A3(_01769_),
    .A4(_01822_),
    .B1(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_2 _08734_ (.A(_01772_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__and2b_1 _08735_ (.A_N(_01828_),
    .B(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_2 _08736_ (.A(_01585_),
    .B(_01773_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand3b_2 _08737_ (.A_N(_01828_),
    .B(_01831_),
    .C(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__a211o_1 _08738_ (.A1(_01772_),
    .A2(_01830_),
    .B1(_01581_),
    .C1(_01638_),
    .X(_01835_));
 sky130_fd_sc_hd__a21o_1 _08739_ (.A1(_01584_),
    .A2(_01835_),
    .B1(_01775_),
    .X(_01836_));
 sky130_fd_sc_hd__nand3_2 _08740_ (.A(_01584_),
    .B(_01775_),
    .C(_01835_),
    .Y(_01837_));
 sky130_fd_sc_hd__a21o_1 _08741_ (.A1(_01836_),
    .A2(_01837_),
    .B1(_01834_),
    .X(_01838_));
 sky130_fd_sc_hd__a21o_1 _08742_ (.A1(_01556_),
    .A2(_01774_),
    .B1(_01522_),
    .X(_01839_));
 sky130_fd_sc_hd__and2_1 _08743_ (.A(_01776_),
    .B(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__a221o_2 _08744_ (.A1(_01836_),
    .A2(_01837_),
    .B1(_01839_),
    .B2(_01776_),
    .C1(_01834_),
    .X(_01841_));
 sky130_fd_sc_hd__a21bo_1 _08745_ (.A1(_01518_),
    .A2(_01583_),
    .B1_N(_01521_),
    .X(_01842_));
 sky130_fd_sc_hd__nand4_2 _08746_ (.A(_01522_),
    .B(_01584_),
    .C(_01775_),
    .D(_01835_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21o_1 _08747_ (.A1(_01842_),
    .A2(_01843_),
    .B1(_01520_),
    .X(_01844_));
 sky130_fd_sc_hd__nand3_1 _08748_ (.A(_01520_),
    .B(_01842_),
    .C(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__and2_1 _08749_ (.A(_01844_),
    .B(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__nor2_1 _08750_ (.A(_01841_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__and3_1 _08751_ (.A(_01519_),
    .B(_01777_),
    .C(_01781_),
    .X(_01848_));
 sky130_fd_sc_hd__a21oi_1 _08752_ (.A1(_01519_),
    .A2(_01777_),
    .B1(_01781_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _08753_ (.A(_01848_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__a2111o_1 _08754_ (.A1(_01844_),
    .A2(_01845_),
    .B1(_01848_),
    .C1(_01849_),
    .D1(_01841_),
    .X(_01851_));
 sky130_fd_sc_hd__a21o_1 _08755_ (.A1(_01445_),
    .A2(_01488_),
    .B1(_01780_),
    .X(_01852_));
 sky130_fd_sc_hd__a211o_1 _08756_ (.A1(_01842_),
    .A2(_01843_),
    .B1(_01520_),
    .C1(_01782_),
    .X(_01853_));
 sky130_fd_sc_hd__a21o_1 _08757_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01779_),
    .X(_01854_));
 sky130_fd_sc_hd__nand3_1 _08758_ (.A(_01779_),
    .B(_01852_),
    .C(_01853_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(_01854_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__and3_1 _08760_ (.A(_01847_),
    .B(_01850_),
    .C(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__and3_1 _08761_ (.A(_01361_),
    .B(_01446_),
    .C(_01783_),
    .X(_01858_));
 sky130_fd_sc_hd__a21oi_1 _08762_ (.A1(_01446_),
    .A2(_01783_),
    .B1(_01361_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _08763_ (.A(_01858_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__a2111o_1 _08764_ (.A1(_01854_),
    .A2(_01855_),
    .B1(_01858_),
    .C1(_01859_),
    .D1(_01851_),
    .X(_01861_));
 sky130_fd_sc_hd__a21o_1 _08765_ (.A1(_01357_),
    .A2(_01408_),
    .B1(_01360_),
    .X(_01862_));
 sky130_fd_sc_hd__a211o_1 _08766_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01362_),
    .C1(_01779_),
    .X(_01863_));
 sky130_fd_sc_hd__nand3_1 _08767_ (.A(_01359_),
    .B(_01862_),
    .C(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21o_1 _08768_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01359_),
    .X(_01865_));
 sky130_fd_sc_hd__nand2_2 _08769_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__and3_1 _08770_ (.A(_01857_),
    .B(_01860_),
    .C(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__or2_1 _08771_ (.A(_01259_),
    .B(_01785_),
    .X(_01868_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(_01259_),
    .B(_01785_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__a221o_1 _08774_ (.A1(_01864_),
    .A2(_01865_),
    .B1(_01868_),
    .B2(_01869_),
    .C1(_01861_),
    .X(_01871_));
 sky130_fd_sc_hd__a21o_1 _08775_ (.A1(_01258_),
    .A2(_01311_),
    .B1(_01257_),
    .X(_01872_));
 sky130_fd_sc_hd__or2_1 _08776_ (.A(_01259_),
    .B(_01359_),
    .X(_01873_));
 sky130_fd_sc_hd__a21o_1 _08777_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__nand3_1 _08778_ (.A(_01264_),
    .B(_01872_),
    .C(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21o_1 _08779_ (.A1(_01872_),
    .A2(_01874_),
    .B1(_01264_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2_1 _08780_ (.A(_01875_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__o21a_1 _08781_ (.A1(_01265_),
    .A2(_01785_),
    .B1(_01788_),
    .X(_01878_));
 sky130_fd_sc_hd__xor2_1 _08782_ (.A(_01157_),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__a211o_2 _08783_ (.A1(_01875_),
    .A2(_01876_),
    .B1(_01879_),
    .C1(_01871_),
    .X(_01880_));
 sky130_fd_sc_hd__a21bo_1 _08784_ (.A1(_01155_),
    .A2(_01156_),
    .B1_N(_01262_),
    .X(_01881_));
 sky130_fd_sc_hd__o21ai_1 _08785_ (.A1(_01155_),
    .A2(_01156_),
    .B1(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__or2_1 _08786_ (.A(_01157_),
    .B(_01264_),
    .X(_01883_));
 sky130_fd_sc_hd__or2_1 _08787_ (.A(_01872_),
    .B(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__a211o_1 _08788_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01873_),
    .C1(_01883_),
    .X(_01885_));
 sky130_fd_sc_hd__and3_1 _08789_ (.A(_01882_),
    .B(_01884_),
    .C(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__xor2_4 _08790_ (.A(_01094_),
    .B(_01886_),
    .X(_01887_));
 sky130_fd_sc_hd__or2_1 _08791_ (.A(_01880_),
    .B(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__nor2_1 _08792_ (.A(_01802_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__a21o_1 _08793_ (.A1(_01030_),
    .A2(_01093_),
    .B1(_01029_),
    .X(_01890_));
 sky130_fd_sc_hd__a311o_2 _08794_ (.A1(_01882_),
    .A2(_01884_),
    .A3(_01885_),
    .B1(_01094_),
    .C1(_01031_),
    .X(_01891_));
 sky130_fd_sc_hd__a21o_1 _08795_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01793_),
    .X(_01892_));
 sky130_fd_sc_hd__nand3_1 _08796_ (.A(_01793_),
    .B(_01890_),
    .C(_01891_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a2111o_1 _08798_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_01802_),
    .C1(_01880_),
    .D1(_01887_),
    .X(_01895_));
 sky130_fd_sc_hd__xnor2_2 _08799_ (.A(_01794_),
    .B(_01796_),
    .Y(_01896_));
 sky130_fd_sc_hd__and3_1 _08800_ (.A(_01889_),
    .B(_01894_),
    .C(_01896_),
    .X(_01897_));
 sky130_fd_sc_hd__nand2b_1 _08801_ (.A_N(_01895_),
    .B(_01896_),
    .Y(_01898_));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(_00898_),
    .A2(_01791_),
    .B1(_01795_),
    .X(_01899_));
 sky130_fd_sc_hd__or2_1 _08803_ (.A(_01793_),
    .B(_01797_),
    .X(_01900_));
 sky130_fd_sc_hd__a211o_1 _08804_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01793_),
    .C1(_01797_),
    .X(_01901_));
 sky130_fd_sc_hd__and3_1 _08805_ (.A(_01798_),
    .B(_01899_),
    .C(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__a21oi_1 _08806_ (.A1(_01899_),
    .A2(_01901_),
    .B1(_01798_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _08807_ (.A(_01902_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_01897_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__or3_1 _08809_ (.A(_01801_),
    .B(_01902_),
    .C(_01903_),
    .X(_01906_));
 sky130_fd_sc_hd__a21oi_4 _08810_ (.A1(_00655_),
    .A2(_00754_),
    .B1(_00753_),
    .Y(_01907_));
 sky130_fd_sc_hd__o21ai_4 _08811_ (.A1(_00748_),
    .A2(_00749_),
    .B1(_00751_),
    .Y(_01908_));
 sky130_fd_sc_hd__o21ai_1 _08812_ (.A1(_00697_),
    .A2(_00708_),
    .B1(_00707_),
    .Y(_01909_));
 sky130_fd_sc_hd__a21o_1 _08813_ (.A1(_00675_),
    .A2(_00680_),
    .B1(_00682_),
    .X(_01910_));
 sky130_fd_sc_hd__o22a_1 _08814_ (.A1(net47),
    .A2(_00294_),
    .B1(_00298_),
    .B2(net45),
    .X(_01911_));
 sky130_fd_sc_hd__xnor2_1 _08815_ (.A(net97),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__a22o_1 _08816_ (.A1(_00211_),
    .A2(net43),
    .B1(net41),
    .B2(_00243_),
    .X(_01913_));
 sky130_fd_sc_hd__xor2_1 _08817_ (.A(net94),
    .B(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__and2_1 _08818_ (.A(_01912_),
    .B(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__nor2_1 _08819_ (.A(_01912_),
    .B(_01914_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _08820_ (.A(_01915_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a22o_1 _08821_ (.A1(_00198_),
    .A2(net37),
    .B1(_00360_),
    .B2(net39),
    .X(_01918_));
 sky130_fd_sc_hd__xor2_1 _08822_ (.A(net91),
    .B(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__xor2_1 _08823_ (.A(_01917_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__xnor2_1 _08824_ (.A(_01910_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__and2b_1 _08825_ (.A_N(_01921_),
    .B(_01909_),
    .X(_01922_));
 sky130_fd_sc_hd__and2b_1 _08826_ (.A_N(_01909_),
    .B(_01921_),
    .X(_01923_));
 sky130_fd_sc_hd__nor2_1 _08827_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__o21bai_1 _08828_ (.A1(_00699_),
    .A2(_00701_),
    .B1_N(_00705_),
    .Y(_01925_));
 sky130_fd_sc_hd__o21ai_2 _08829_ (.A1(_00686_),
    .A2(_00696_),
    .B1(_00695_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _08830_ (.A(_00730_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__xor2_1 _08831_ (.A(_00730_),
    .B(_01926_),
    .X(_01928_));
 sky130_fd_sc_hd__xnor2_1 _08832_ (.A(_01925_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__o22a_1 _08833_ (.A1(net52),
    .A2(net105),
    .B1(net103),
    .B2(net50),
    .X(_01930_));
 sky130_fd_sc_hd__xnor2_2 _08834_ (.A(net135),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__o22a_1 _08835_ (.A1(net58),
    .A2(_00145_),
    .B1(net145),
    .B2(net56),
    .X(_01932_));
 sky130_fd_sc_hd__xnor2_2 _08836_ (.A(net189),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_01931_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xor2_2 _08838_ (.A(_01931_),
    .B(_01933_),
    .X(_01935_));
 sky130_fd_sc_hd__o22a_1 _08839_ (.A1(net62),
    .A2(net134),
    .B1(net132),
    .B2(net60),
    .X(_01936_));
 sky130_fd_sc_hd__xnor2_2 _08840_ (.A(net172),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__inv_2 _08841_ (.A(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__xnor2_1 _08842_ (.A(_01935_),
    .B(_01937_),
    .Y(_01939_));
 sky130_fd_sc_hd__o22a_1 _08843_ (.A1(net100),
    .A2(net85),
    .B1(net81),
    .B2(net98),
    .X(_01940_));
 sky130_fd_sc_hd__xnor2_1 _08844_ (.A(net137),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__o22a_1 _08845_ (.A1(net34),
    .A2(net76),
    .B1(net72),
    .B2(net32),
    .X(_01942_));
 sky130_fd_sc_hd__xnor2_1 _08846_ (.A(net125),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__and2b_1 _08847_ (.A_N(_01941_),
    .B(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__xor2_1 _08848_ (.A(_01941_),
    .B(_01943_),
    .X(_01945_));
 sky130_fd_sc_hd__o22a_1 _08849_ (.A1(net83),
    .A2(net77),
    .B1(net73),
    .B2(net79),
    .X(_01946_));
 sky130_fd_sc_hd__xnor2_1 _08850_ (.A(net121),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__or2_1 _08851_ (.A(_01945_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_01945_),
    .B(_01947_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _08853_ (.A(_01948_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__o22a_1 _08854_ (.A1(net149),
    .A2(net55),
    .B1(net16),
    .B2(net151),
    .X(_01951_));
 sky130_fd_sc_hd__xnor2_2 _08855_ (.A(net192),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__a31o_2 _08856_ (.A1(_04801_),
    .A2(_04888_),
    .A3(_06549_),
    .B1(net174),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_4 _08857_ (.A(_04975_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__xnor2_2 _08858_ (.A(_04964_),
    .B(_01953_),
    .Y(_01955_));
 sky130_fd_sc_hd__a22o_1 _08859_ (.A1(_06494_),
    .A2(_00690_),
    .B1(_01954_),
    .B2(net292),
    .X(_01956_));
 sky130_fd_sc_hd__xnor2_2 _08860_ (.A(_06468_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__o22a_1 _08861_ (.A1(net67),
    .A2(net155),
    .B1(net153),
    .B2(net64),
    .X(_01958_));
 sky130_fd_sc_hd__xnor2_2 _08862_ (.A(net194),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__or2_1 _08863_ (.A(_01957_),
    .B(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__xnor2_2 _08864_ (.A(_01957_),
    .B(_01959_),
    .Y(_01961_));
 sky130_fd_sc_hd__xor2_2 _08865_ (.A(_01952_),
    .B(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__xnor2_1 _08866_ (.A(_01950_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_1 _08867_ (.A(_01939_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__or4_2 _08868_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_00218_),
    .D(_00439_),
    .X(_01965_));
 sky130_fd_sc_hd__o41a_1 _08869_ (.A1(reg1_val[28]),
    .A2(reg1_val[29]),
    .A3(_00218_),
    .A4(_00439_),
    .B1(net262),
    .X(_01966_));
 sky130_fd_sc_hd__xnor2_2 _08870_ (.A(reg1_val[30]),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__or2_2 _08871_ (.A(net68),
    .B(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_1 _08872_ (.A(net68),
    .B(_01967_),
    .Y(_01969_));
 sky130_fd_sc_hd__and2_1 _08873_ (.A(_01968_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_01968_),
    .B(_01969_),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_2 _08875_ (.A(net210),
    .B(net10),
    .Y(_01972_));
 sky130_fd_sc_hd__o22a_1 _08876_ (.A1(_00249_),
    .A2(net23),
    .B1(net15),
    .B2(net143),
    .X(_01973_));
 sky130_fd_sc_hd__xnor2_2 _08877_ (.A(net70),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__xor2_2 _08878_ (.A(_01972_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__or2_1 _08879_ (.A(_01964_),
    .B(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__xnor2_1 _08880_ (.A(_01964_),
    .B(_01975_),
    .Y(_01977_));
 sky130_fd_sc_hd__xor2_1 _08881_ (.A(_01929_),
    .B(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__a21oi_1 _08882_ (.A1(_00663_),
    .A2(_00665_),
    .B1(_00661_),
    .Y(_01979_));
 sky130_fd_sc_hd__o22a_1 _08883_ (.A1(net120),
    .A2(net26),
    .B1(net24),
    .B2(net117),
    .X(_01980_));
 sky130_fd_sc_hd__xnor2_1 _08884_ (.A(net87),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a22o_1 _08885_ (.A1(net30),
    .A2(_00309_),
    .B1(_00315_),
    .B2(net28),
    .X(_01982_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(net48),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__and2_1 _08887_ (.A(_01981_),
    .B(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__nor2_1 _08888_ (.A(_01981_),
    .B(_01983_),
    .Y(_01985_));
 sky130_fd_sc_hd__or2_1 _08889_ (.A(_01984_),
    .B(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__a21oi_1 _08890_ (.A1(_00714_),
    .A2(_00719_),
    .B1(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__and3_1 _08891_ (.A(_00714_),
    .B(_00719_),
    .C(_01986_),
    .X(_01988_));
 sky130_fd_sc_hd__nor2_1 _08892_ (.A(_01987_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__and2b_1 _08893_ (.A_N(_01979_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__xnor2_1 _08894_ (.A(_01979_),
    .B(_01989_),
    .Y(_01991_));
 sky130_fd_sc_hd__and2_1 _08895_ (.A(_01978_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__nor2_1 _08896_ (.A(_01978_),
    .B(_01991_),
    .Y(_01993_));
 sky130_fd_sc_hd__nor2_1 _08897_ (.A(_01992_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__xor2_2 _08898_ (.A(_01924_),
    .B(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__a21o_1 _08899_ (.A1(_00674_),
    .A2(_00740_),
    .B1(_00738_),
    .X(_01996_));
 sky130_fd_sc_hd__o21bai_4 _08900_ (.A1(_00656_),
    .A2(_00672_),
    .B1_N(_00671_),
    .Y(_01997_));
 sky130_fd_sc_hd__a21o_2 _08901_ (.A1(_00684_),
    .A2(_00723_),
    .B1(_00722_),
    .X(_01998_));
 sky130_fd_sc_hd__nor2_2 _08902_ (.A(_00733_),
    .B(_00736_),
    .Y(_01999_));
 sky130_fd_sc_hd__o21ai_1 _08903_ (.A1(_00733_),
    .A2(_00736_),
    .B1(_01998_),
    .Y(_02000_));
 sky130_fd_sc_hd__xnor2_4 _08904_ (.A(_01998_),
    .B(_01999_),
    .Y(_02001_));
 sky130_fd_sc_hd__xnor2_2 _08905_ (.A(_01997_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__a21oi_2 _08906_ (.A1(_00743_),
    .A2(_00747_),
    .B1(_00746_),
    .Y(_02003_));
 sky130_fd_sc_hd__xnor2_1 _08907_ (.A(_02002_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2b_1 _08908_ (.A_N(_02004_),
    .B(_01996_),
    .Y(_02005_));
 sky130_fd_sc_hd__xnor2_2 _08909_ (.A(_01996_),
    .B(_02004_),
    .Y(_02006_));
 sky130_fd_sc_hd__xnor2_2 _08910_ (.A(_01995_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2b_1 _08911_ (.A_N(_02007_),
    .B(_01908_),
    .Y(_02008_));
 sky130_fd_sc_hd__xor2_4 _08912_ (.A(_01908_),
    .B(_02007_),
    .X(_02009_));
 sky130_fd_sc_hd__or2_1 _08913_ (.A(_01907_),
    .B(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__and2_1 _08914_ (.A(_01907_),
    .B(_02009_),
    .X(_02011_));
 sky130_fd_sc_hd__xnor2_4 _08915_ (.A(_01907_),
    .B(_02009_),
    .Y(_02012_));
 sky130_fd_sc_hd__o22a_1 _08916_ (.A1(_00654_),
    .A2(_00755_),
    .B1(_00758_),
    .B2(_00827_),
    .X(_02013_));
 sky130_fd_sc_hd__a21o_1 _08917_ (.A1(_00654_),
    .A2(_00755_),
    .B1(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__or2_1 _08918_ (.A(_00757_),
    .B(_01799_),
    .X(_02015_));
 sky130_fd_sc_hd__a211o_1 _08919_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_00757_),
    .C1(_01799_),
    .X(_02016_));
 sky130_fd_sc_hd__o221a_2 _08920_ (.A1(_01899_),
    .A2(_02015_),
    .B1(_02016_),
    .B2(_01900_),
    .C1(_02014_),
    .X(_02017_));
 sky130_fd_sc_hd__xor2_2 _08921_ (.A(_02012_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__or3_1 _08922_ (.A(_01898_),
    .B(_01906_),
    .C(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__a21bo_2 _08923_ (.A1(_01995_),
    .A2(_02006_),
    .B1_N(_02008_),
    .X(_02020_));
 sky130_fd_sc_hd__o21ai_4 _08924_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_02005_),
    .Y(_02021_));
 sky130_fd_sc_hd__a32o_1 _08925_ (.A1(_01948_),
    .A2(_01949_),
    .A3(_01962_),
    .B1(_01963_),
    .B2(_01939_),
    .X(_02022_));
 sky130_fd_sc_hd__o22a_1 _08926_ (.A1(net45),
    .A2(_00294_),
    .B1(net108),
    .B2(net47),
    .X(_02023_));
 sky130_fd_sc_hd__xnor2_1 _08927_ (.A(net97),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__a22o_1 _08928_ (.A1(_00198_),
    .A2(net43),
    .B1(net41),
    .B2(_00211_),
    .X(_02025_));
 sky130_fd_sc_hd__xor2_1 _08929_ (.A(net94),
    .B(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__and2_1 _08930_ (.A(_02024_),
    .B(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__nor2_1 _08931_ (.A(_02024_),
    .B(_02026_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _08932_ (.A(_02027_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__a22o_1 _08933_ (.A1(net39),
    .A2(net112),
    .B1(_00360_),
    .B2(net37),
    .X(_02030_));
 sky130_fd_sc_hd__xor2_2 _08934_ (.A(net91),
    .B(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__xor2_2 _08935_ (.A(_02029_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__a21bo_1 _08936_ (.A1(_01925_),
    .A2(_01928_),
    .B1_N(_01927_),
    .X(_02033_));
 sky130_fd_sc_hd__xnor2_1 _08937_ (.A(_02032_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__and2b_1 _08938_ (.A_N(_02034_),
    .B(_02022_),
    .X(_02035_));
 sky130_fd_sc_hd__and2b_1 _08939_ (.A_N(_02022_),
    .B(_02034_),
    .X(_02036_));
 sky130_fd_sc_hd__nor2_2 _08940_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__and2b_1 _08941_ (.A_N(_01944_),
    .B(_01948_),
    .X(_02038_));
 sky130_fd_sc_hd__a21oi_2 _08942_ (.A1(_01935_),
    .A2(_01938_),
    .B1(_01934_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2b_1 _08943_ (.A_N(_02039_),
    .B(_01984_),
    .Y(_02040_));
 sky130_fd_sc_hd__xnor2_2 _08944_ (.A(_01984_),
    .B(_02039_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2b_1 _08945_ (.A_N(_02038_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__xnor2_2 _08946_ (.A(_02038_),
    .B(_02041_),
    .Y(_02043_));
 sky130_fd_sc_hd__o22a_1 _08947_ (.A1(net60),
    .A2(net105),
    .B1(net103),
    .B2(net52),
    .X(_02044_));
 sky130_fd_sc_hd__xnor2_1 _08948_ (.A(net135),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__o22a_1 _08949_ (.A1(net64),
    .A2(net147),
    .B1(net145),
    .B2(net58),
    .X(_02046_));
 sky130_fd_sc_hd__xnor2_1 _08950_ (.A(net189),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _08951_ (.A(_02045_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__xor2_1 _08952_ (.A(_02045_),
    .B(_02047_),
    .X(_02049_));
 sky130_fd_sc_hd__o22a_1 _08953_ (.A1(net56),
    .A2(net134),
    .B1(net132),
    .B2(net62),
    .X(_02050_));
 sky130_fd_sc_hd__xnor2_1 _08954_ (.A(net172),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__and2b_1 _08955_ (.A_N(_02051_),
    .B(_02049_),
    .X(_02052_));
 sky130_fd_sc_hd__and2b_1 _08956_ (.A_N(_02049_),
    .B(_02051_),
    .X(_02053_));
 sky130_fd_sc_hd__nor2_1 _08957_ (.A(_02052_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__o22a_1 _08958_ (.A1(net50),
    .A2(net85),
    .B1(net81),
    .B2(net100),
    .X(_02055_));
 sky130_fd_sc_hd__xnor2_1 _08959_ (.A(net137),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__o22a_1 _08960_ (.A1(net34),
    .A2(net80),
    .B1(net76),
    .B2(net32),
    .X(_02057_));
 sky130_fd_sc_hd__xnor2_1 _08961_ (.A(net125),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__and2b_1 _08962_ (.A_N(_02056_),
    .B(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__xor2_1 _08963_ (.A(_02056_),
    .B(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__o22a_1 _08964_ (.A1(net98),
    .A2(net77),
    .B1(net73),
    .B2(net84),
    .X(_02061_));
 sky130_fd_sc_hd__xnor2_1 _08965_ (.A(net121),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__or2_1 _08966_ (.A(_02060_),
    .B(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(_02060_),
    .B(_02062_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(_02063_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__o22a_2 _08969_ (.A1(net149),
    .A2(net16),
    .B1(net13),
    .B2(net151),
    .X(_02066_));
 sky130_fd_sc_hd__xnor2_4 _08970_ (.A(net192),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__or4_1 _08971_ (.A(_04812_),
    .B(_04899_),
    .C(_04975_),
    .D(_06550_),
    .X(_02068_));
 sky130_fd_sc_hd__a21oi_2 _08972_ (.A1(net295),
    .A2(_02068_),
    .B1(_05247_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21o_1 _08973_ (.A1(net295),
    .A2(_02068_),
    .B1(_05247_),
    .X(_02070_));
 sky130_fd_sc_hd__o22a_2 _08974_ (.A1(_06495_),
    .A2(net11),
    .B1(net7),
    .B2(net288),
    .X(_02071_));
 sky130_fd_sc_hd__xnor2_4 _08975_ (.A(net239),
    .B(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__o22a_2 _08976_ (.A1(net67),
    .A2(net153),
    .B1(net55),
    .B2(net155),
    .X(_02073_));
 sky130_fd_sc_hd__xnor2_4 _08977_ (.A(net194),
    .B(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__or2_1 _08978_ (.A(_02072_),
    .B(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__xnor2_4 _08979_ (.A(_02072_),
    .B(_02074_),
    .Y(_02076_));
 sky130_fd_sc_hd__xor2_4 _08980_ (.A(_02067_),
    .B(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__xnor2_2 _08981_ (.A(_02065_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__xnor2_2 _08982_ (.A(_02054_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(reg1_val[30]),
    .B(_01965_),
    .Y(_02080_));
 sky130_fd_sc_hd__o21a_4 _08984_ (.A1(net286),
    .A2(_02080_),
    .B1(reg1_val[31]),
    .X(_02081_));
 sky130_fd_sc_hd__o21ai_4 _08985_ (.A1(net286),
    .A2(_02080_),
    .B1(reg1_val[31]),
    .Y(_02082_));
 sky130_fd_sc_hd__a2111o_1 _08986_ (.A1(net295),
    .A2(_01965_),
    .B1(_00668_),
    .C1(reg1_val[30]),
    .D1(_04427_),
    .X(_02083_));
 sky130_fd_sc_hd__o21a_1 _08987_ (.A1(_01968_),
    .A2(net21),
    .B1(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__o21ai_2 _08988_ (.A1(_01968_),
    .A2(net21),
    .B1(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__o22a_1 _08989_ (.A1(net143),
    .A2(net10),
    .B1(net5),
    .B2(net210),
    .X(_02086_));
 sky130_fd_sc_hd__xnor2_2 _08990_ (.A(net20),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__o21a_1 _08991_ (.A1(_01952_),
    .A2(_01961_),
    .B1(_01960_),
    .X(_02088_));
 sky130_fd_sc_hd__o22a_1 _08992_ (.A1(_00242_),
    .A2(net23),
    .B1(net15),
    .B2(_00249_),
    .X(_02089_));
 sky130_fd_sc_hd__xnor2_2 _08993_ (.A(_00668_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__and2b_1 _08994_ (.A_N(_02088_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__xor2_2 _08995_ (.A(_02088_),
    .B(_02090_),
    .X(_02092_));
 sky130_fd_sc_hd__xnor2_2 _08996_ (.A(_02087_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_1 _08997_ (.A(_02079_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__xor2_2 _08998_ (.A(_02079_),
    .B(_02093_),
    .X(_02095_));
 sky130_fd_sc_hd__xor2_1 _08999_ (.A(_02043_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__a21o_1 _09000_ (.A1(_01917_),
    .A2(_01919_),
    .B1(_01915_),
    .X(_02097_));
 sky130_fd_sc_hd__o22a_1 _09001_ (.A1(net120),
    .A2(net24),
    .B1(net72),
    .B2(net26),
    .X(_02098_));
 sky130_fd_sc_hd__xnor2_1 _09002_ (.A(net87),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__a22o_1 _09003_ (.A1(net115),
    .A2(net30),
    .B1(net28),
    .B2(_00309_),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_1 _09004_ (.A(net48),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__and2_1 _09005_ (.A(_02099_),
    .B(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_1 _09006_ (.A(_02099_),
    .B(_02101_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _09007_ (.A(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _09008_ (.A(_01972_),
    .B(net21),
    .Y(_02105_));
 sky130_fd_sc_hd__a21oi_2 _09009_ (.A1(_01972_),
    .A2(_01974_),
    .B1(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__xnor2_1 _09010_ (.A(_02104_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__and2b_1 _09011_ (.A_N(_02107_),
    .B(_02097_),
    .X(_02108_));
 sky130_fd_sc_hd__xnor2_1 _09012_ (.A(_02097_),
    .B(_02107_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(_02096_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__or2_1 _09014_ (.A(_02096_),
    .B(_02109_),
    .X(_02111_));
 sky130_fd_sc_hd__and2_2 _09015_ (.A(_02110_),
    .B(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__xor2_4 _09016_ (.A(_02037_),
    .B(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__a21o_1 _09017_ (.A1(_01924_),
    .A2(_01994_),
    .B1(_01992_),
    .X(_02114_));
 sky130_fd_sc_hd__a21o_2 _09018_ (.A1(_01910_),
    .A2(_01920_),
    .B1(_01922_),
    .X(_02115_));
 sky130_fd_sc_hd__o21a_2 _09019_ (.A1(_01929_),
    .A2(_01977_),
    .B1(_01976_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_2 _09020_ (.A(_01987_),
    .B(_01990_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _09021_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__xor2_4 _09022_ (.A(_02116_),
    .B(_02117_),
    .X(_02119_));
 sky130_fd_sc_hd__xnor2_4 _09023_ (.A(_02115_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21boi_4 _09024_ (.A1(_01997_),
    .A2(_02001_),
    .B1_N(_02000_),
    .Y(_02121_));
 sky130_fd_sc_hd__xnor2_2 _09025_ (.A(_02120_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2b_1 _09026_ (.A_N(_02122_),
    .B(_02114_),
    .Y(_02123_));
 sky130_fd_sc_hd__xnor2_2 _09027_ (.A(_02114_),
    .B(_02122_),
    .Y(_02124_));
 sky130_fd_sc_hd__and2_1 _09028_ (.A(_02113_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__xor2_4 _09029_ (.A(_02113_),
    .B(_02124_),
    .X(_02126_));
 sky130_fd_sc_hd__xor2_4 _09030_ (.A(_02021_),
    .B(_02126_),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _09031_ (.A(_02020_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__xor2_2 _09032_ (.A(_02020_),
    .B(_02127_),
    .X(_02129_));
 sky130_fd_sc_hd__xnor2_2 _09033_ (.A(_02020_),
    .B(_02127_),
    .Y(_02130_));
 sky130_fd_sc_hd__a21oi_1 _09034_ (.A1(_00756_),
    .A2(_02010_),
    .B1(_02011_),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2_1 _09035_ (.A(_00757_),
    .B(_02012_),
    .Y(_02132_));
 sky130_fd_sc_hd__a21oi_2 _09036_ (.A1(_01800_),
    .A2(_02132_),
    .B1(_02131_),
    .Y(_02133_));
 sky130_fd_sc_hd__xnor2_2 _09037_ (.A(_02129_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__or4_2 _09038_ (.A(_01898_),
    .B(_01906_),
    .C(_02018_),
    .D(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__a2111o_1 _09039_ (.A1(_01899_),
    .A2(_01901_),
    .B1(_02012_),
    .C1(_02015_),
    .D1(_02130_),
    .X(_02136_));
 sky130_fd_sc_hd__a21boi_1 _09040_ (.A1(_02020_),
    .A2(_02127_),
    .B1_N(_02010_),
    .Y(_02137_));
 sky130_fd_sc_hd__o32a_1 _09041_ (.A1(_02012_),
    .A2(_02014_),
    .A3(_02130_),
    .B1(_02137_),
    .B2(_02128_),
    .X(_02138_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_02136_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__a21oi_4 _09043_ (.A1(_02021_),
    .A2(_02126_),
    .B1(_02125_),
    .Y(_02140_));
 sky130_fd_sc_hd__o21ai_4 _09044_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_02123_),
    .Y(_02141_));
 sky130_fd_sc_hd__a32o_2 _09045_ (.A1(_02063_),
    .A2(_02064_),
    .A3(_02077_),
    .B1(_02078_),
    .B2(_02054_),
    .X(_02142_));
 sky130_fd_sc_hd__o22a_1 _09046_ (.A1(net128),
    .A2(net23),
    .B1(net15),
    .B2(_00242_),
    .X(_02143_));
 sky130_fd_sc_hd__xnor2_1 _09047_ (.A(net70),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__inv_2 _09048_ (.A(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__a22o_1 _09049_ (.A1(net39),
    .A2(_00293_),
    .B1(net112),
    .B2(net37),
    .X(_02146_));
 sky130_fd_sc_hd__xor2_1 _09050_ (.A(net91),
    .B(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__xor2_1 _09051_ (.A(_02144_),
    .B(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_1 _09052_ (.A1(_00198_),
    .A2(net41),
    .B1(_00360_),
    .B2(net43),
    .X(_02149_));
 sky130_fd_sc_hd__xor2_1 _09053_ (.A(net94),
    .B(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__and2b_1 _09054_ (.A_N(_02148_),
    .B(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__and2b_1 _09055_ (.A_N(_02150_),
    .B(_02148_),
    .X(_02152_));
 sky130_fd_sc_hd__or2_1 _09056_ (.A(_02151_),
    .B(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__a21o_1 _09057_ (.A1(_02040_),
    .A2(_02042_),
    .B1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__nand3_1 _09058_ (.A(_02040_),
    .B(_02042_),
    .C(_02153_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_2 _09059_ (.A(_02154_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2b_1 _09060_ (.A_N(_02156_),
    .B(_02142_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_4 _09061_ (.A(_02142_),
    .B(_02156_),
    .Y(_02158_));
 sky130_fd_sc_hd__and2b_1 _09062_ (.A_N(_02059_),
    .B(_02063_),
    .X(_02159_));
 sky130_fd_sc_hd__o21ai_1 _09063_ (.A1(_02048_),
    .A2(_02052_),
    .B1(_02102_),
    .Y(_02160_));
 sky130_fd_sc_hd__or3_1 _09064_ (.A(_02048_),
    .B(_02052_),
    .C(_02102_),
    .X(_02161_));
 sky130_fd_sc_hd__and2_1 _09065_ (.A(_02160_),
    .B(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__nand2b_1 _09066_ (.A_N(_02159_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__xnor2_2 _09067_ (.A(_02159_),
    .B(_02162_),
    .Y(_02164_));
 sky130_fd_sc_hd__o22a_1 _09068_ (.A1(net67),
    .A2(net147),
    .B1(net145),
    .B2(net64),
    .X(_02165_));
 sky130_fd_sc_hd__xnor2_2 _09069_ (.A(net189),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__o22a_1 _09070_ (.A1(net62),
    .A2(net105),
    .B1(net103),
    .B2(net60),
    .X(_02167_));
 sky130_fd_sc_hd__xnor2_2 _09071_ (.A(net135),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _09072_ (.A(_02166_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__xor2_2 _09073_ (.A(_02166_),
    .B(_02168_),
    .X(_02170_));
 sky130_fd_sc_hd__o22a_1 _09074_ (.A1(net58),
    .A2(net134),
    .B1(net132),
    .B2(net56),
    .X(_02171_));
 sky130_fd_sc_hd__xnor2_2 _09075_ (.A(net172),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__inv_2 _09076_ (.A(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__xnor2_2 _09077_ (.A(_02170_),
    .B(_02172_),
    .Y(_02174_));
 sky130_fd_sc_hd__o22a_1 _09078_ (.A1(net52),
    .A2(net85),
    .B1(net81),
    .B2(net50),
    .X(_02175_));
 sky130_fd_sc_hd__xnor2_1 _09079_ (.A(net137),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__o22a_1 _09080_ (.A1(net34),
    .A2(net84),
    .B1(net80),
    .B2(net32),
    .X(_02177_));
 sky130_fd_sc_hd__xnor2_1 _09081_ (.A(net125),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__and2b_1 _09082_ (.A_N(_02176_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__xor2_1 _09083_ (.A(_02176_),
    .B(_02178_),
    .X(_02180_));
 sky130_fd_sc_hd__o22a_1 _09084_ (.A1(net100),
    .A2(net77),
    .B1(net73),
    .B2(net99),
    .X(_02181_));
 sky130_fd_sc_hd__xnor2_1 _09085_ (.A(net121),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _09086_ (.A(_02180_),
    .B(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(_02180_),
    .B(_02182_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(_02183_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__o22a_1 _09089_ (.A1(net149),
    .A2(net13),
    .B1(net11),
    .B2(net151),
    .X(_02186_));
 sky130_fd_sc_hd__xor2_1 _09090_ (.A(net192),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__o32a_1 _09091_ (.A1(net155),
    .A2(_00395_),
    .A3(_00397_),
    .B1(net153),
    .B2(net55),
    .X(_02188_));
 sky130_fd_sc_hd__xnor2_1 _09092_ (.A(_06507_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_1 _09093_ (.A1(net287),
    .A2(net8),
    .B1(net239),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_02189_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__xor2_1 _09095_ (.A(_02189_),
    .B(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_02187_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__or2_1 _09097_ (.A(_02187_),
    .B(_02192_),
    .X(_02194_));
 sky130_fd_sc_hd__and2_2 _09098_ (.A(_02193_),
    .B(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__xnor2_2 _09099_ (.A(_02185_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__xnor2_2 _09100_ (.A(_02174_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _09101_ (.A(_06341_),
    .B(net20),
    .Y(_02198_));
 sky130_fd_sc_hd__o21ai_2 _09102_ (.A1(_02067_),
    .A2(_02076_),
    .B1(_02075_),
    .Y(_02199_));
 sky130_fd_sc_hd__o22a_1 _09103_ (.A1(_00249_),
    .A2(net10),
    .B1(net5),
    .B2(net143),
    .X(_02200_));
 sky130_fd_sc_hd__xnor2_2 _09104_ (.A(net21),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(_02199_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__xor2_2 _09106_ (.A(_02199_),
    .B(_02201_),
    .X(_02203_));
 sky130_fd_sc_hd__xnor2_2 _09107_ (.A(_02198_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _09108_ (.A(_02197_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__xor2_2 _09109_ (.A(_02197_),
    .B(_02204_),
    .X(_02206_));
 sky130_fd_sc_hd__xnor2_1 _09110_ (.A(_02164_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a21o_1 _09111_ (.A1(_02029_),
    .A2(_02031_),
    .B1(_02027_),
    .X(_02208_));
 sky130_fd_sc_hd__o22a_1 _09112_ (.A1(net26),
    .A2(net76),
    .B1(net72),
    .B2(net24),
    .X(_02209_));
 sky130_fd_sc_hd__xnor2_1 _09113_ (.A(_00286_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__o22a_1 _09114_ (.A1(net47),
    .A2(net111),
    .B1(net109),
    .B2(net45),
    .X(_02211_));
 sky130_fd_sc_hd__xnor2_1 _09115_ (.A(net97),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__and2_1 _09116_ (.A(_02210_),
    .B(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__xor2_1 _09117_ (.A(_02210_),
    .B(_02212_),
    .X(_02214_));
 sky130_fd_sc_hd__a22o_1 _09118_ (.A1(net118),
    .A2(net30),
    .B1(net28),
    .B2(net115),
    .X(_02215_));
 sky130_fd_sc_hd__xnor2_1 _09119_ (.A(net49),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__xor2_1 _09120_ (.A(_02214_),
    .B(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__o21ba_1 _09121_ (.A1(_02087_),
    .A2(_02092_),
    .B1_N(_02091_),
    .X(_02218_));
 sky130_fd_sc_hd__and2b_1 _09122_ (.A_N(_02218_),
    .B(_02217_),
    .X(_02219_));
 sky130_fd_sc_hd__xnor2_1 _09123_ (.A(_02217_),
    .B(_02218_),
    .Y(_02220_));
 sky130_fd_sc_hd__xnor2_1 _09124_ (.A(_02208_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _09125_ (.A(_02207_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand2_1 _09126_ (.A(_02207_),
    .B(_02221_),
    .Y(_02223_));
 sky130_fd_sc_hd__and2b_1 _09127_ (.A_N(_02222_),
    .B(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__xor2_4 _09128_ (.A(_02158_),
    .B(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__a21bo_2 _09129_ (.A1(_02037_),
    .A2(_02112_),
    .B1_N(_02110_),
    .X(_02226_));
 sky130_fd_sc_hd__a21o_1 _09130_ (.A1(_02032_),
    .A2(_02033_),
    .B1(_02035_),
    .X(_02227_));
 sky130_fd_sc_hd__a21oi_2 _09131_ (.A1(_02043_),
    .A2(_02095_),
    .B1(_02094_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21oi_2 _09132_ (.A1(_02104_),
    .A2(_02106_),
    .B1(_02108_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _09133_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__xor2_2 _09134_ (.A(_02228_),
    .B(_02229_),
    .X(_02231_));
 sky130_fd_sc_hd__xnor2_2 _09135_ (.A(_02227_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_4 _09136_ (.A1(_02115_),
    .A2(_02119_),
    .B1(_02118_),
    .Y(_02233_));
 sky130_fd_sc_hd__xnor2_2 _09137_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2b_1 _09138_ (.A_N(_02234_),
    .B(_02226_),
    .Y(_02235_));
 sky130_fd_sc_hd__xnor2_4 _09139_ (.A(_02226_),
    .B(_02234_),
    .Y(_02236_));
 sky130_fd_sc_hd__and2_1 _09140_ (.A(_02225_),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__xor2_4 _09141_ (.A(_02225_),
    .B(_02236_),
    .X(_02238_));
 sky130_fd_sc_hd__xnor2_4 _09142_ (.A(_02141_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _09143_ (.A(_02140_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__xor2_1 _09144_ (.A(_02140_),
    .B(_02239_),
    .X(_02241_));
 sky130_fd_sc_hd__xnor2_4 _09145_ (.A(_02140_),
    .B(_02239_),
    .Y(_02242_));
 sky130_fd_sc_hd__xnor2_2 _09146_ (.A(_02139_),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__a21oi_1 _09147_ (.A1(net162),
    .A2(_02135_),
    .B1(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_4 _09148_ (.A(_06430_),
    .B(_06436_),
    .Y(_02245_));
 sky130_fd_sc_hd__or2_2 _09149_ (.A(_06430_),
    .B(_06436_),
    .X(_02246_));
 sky130_fd_sc_hd__a311o_1 _09150_ (.A1(net162),
    .A2(_02135_),
    .A3(_02243_),
    .B1(_02244_),
    .C1(net187),
    .X(_02247_));
 sky130_fd_sc_hd__or3b_1 _09151_ (.A(_06415_),
    .B(_06459_),
    .C_N(_06413_),
    .X(_02248_));
 sky130_fd_sc_hd__nor2_1 _09152_ (.A(net284),
    .B(_06453_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_2 _09153_ (.A(net294),
    .B(_06452_),
    .Y(_02250_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(net289),
    .A1(reg1_val[30]),
    .S(net169),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(net293),
    .A1(reg1_val[31]),
    .S(net170),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(_02251_),
    .A1(_02252_),
    .S(net210),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net169),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net169),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(_02254_),
    .A1(_02255_),
    .S(net207),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(_02253_),
    .A1(_02256_),
    .S(net212),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net169),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net169),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(_02258_),
    .A1(_02259_),
    .S(net207),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net169),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net169),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(_02261_),
    .A1(_02262_),
    .S(net207),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(_02260_),
    .A1(_02263_),
    .S(net211),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(_02257_),
    .A1(_02264_),
    .S(net214),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net169),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net169),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(_02266_),
    .A1(_02267_),
    .S(net207),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net169),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net169),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(_02269_),
    .A1(_02270_),
    .S(net205),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(_02268_),
    .A1(_02271_),
    .S(net211),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net169),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net169),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_02273_),
    .A1(_02274_),
    .S(net205),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(net291),
    .A1(reg1_val[17]),
    .S(net169),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(net290),
    .A1(reg1_val[16]),
    .S(net169),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(_02276_),
    .A1(_02277_),
    .S(net205),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(_02275_),
    .A1(_02278_),
    .S(net211),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _09183_ (.A0(_02272_),
    .A1(_02279_),
    .S(net214),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(_02265_),
    .A1(_02280_),
    .S(net217),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net167),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net167),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(_02282_),
    .A1(_02283_),
    .S(net205),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net167),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _09189_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net167),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(_02285_),
    .A1(_02286_),
    .S(net206),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _09191_ (.A0(_02284_),
    .A1(_02287_),
    .S(net212),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net167),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net167),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(_02289_),
    .A1(_02290_),
    .S(net206),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(net289),
    .A1(reg1_val[30]),
    .S(net168),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net293),
    .A1(reg1_val[31]),
    .S(net168),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(_02292_),
    .A1(_02293_),
    .S(net206),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(_02291_),
    .A1(_02294_),
    .S(net212),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(_02288_),
    .A1(_02295_),
    .S(net214),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net290),
    .A1(reg1_val[16]),
    .S(net167),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net291),
    .A1(reg1_val[17]),
    .S(net167),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(_02297_),
    .A1(_02298_),
    .S(net205),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net167),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net167),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(_02300_),
    .A1(_02301_),
    .S(net205),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(_02299_),
    .A1(_02302_),
    .S(net212),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net167),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net167),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(_02304_),
    .A1(_02305_),
    .S(net205),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net167),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net167),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(_02307_),
    .A1(_02308_),
    .S(net205),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(_02306_),
    .A1(_02309_),
    .S(net212),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(_02303_),
    .A1(_02310_),
    .S(net215),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(_02296_),
    .A1(_02311_),
    .S(net219),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(_02281_),
    .A1(_02312_),
    .S(net220),
    .X(_02313_));
 sky130_fd_sc_hd__inv_2 _09217_ (.A(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(net293),
    .B(curr_PC[0]),
    .Y(_02315_));
 sky130_fd_sc_hd__or2_1 _09219_ (.A(net293),
    .B(curr_PC[0]),
    .X(_02316_));
 sky130_fd_sc_hd__a21oi_2 _09220_ (.A1(_02315_),
    .A2(_02316_),
    .B1(net223),
    .Y(_02317_));
 sky130_fd_sc_hd__a211o_1 _09221_ (.A1(net224),
    .A2(_02314_),
    .B1(_02317_),
    .C1(net196),
    .X(_02318_));
 sky130_fd_sc_hd__nor2_4 _09222_ (.A(net294),
    .B(_06453_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_8 _09223_ (.A(net284),
    .B(_06452_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_4 _09224_ (.A(_06451_),
    .B(_06459_),
    .Y(_02321_));
 sky130_fd_sc_hd__or2_2 _09225_ (.A(_06451_),
    .B(_06459_),
    .X(_02322_));
 sky130_fd_sc_hd__nor2_8 _09226_ (.A(_06415_),
    .B(_06450_),
    .Y(_02323_));
 sky130_fd_sc_hd__or2_1 _09227_ (.A(_06415_),
    .B(_06450_),
    .X(_02324_));
 sky130_fd_sc_hd__nor2_4 _09228_ (.A(_06428_),
    .B(_06459_),
    .Y(_02325_));
 sky130_fd_sc_hd__or2_1 _09229_ (.A(_06428_),
    .B(_06459_),
    .X(_02326_));
 sky130_fd_sc_hd__a21o_1 _09230_ (.A1(net236),
    .A2(net235),
    .B1(_06416_),
    .X(_02327_));
 sky130_fd_sc_hd__a21oi_1 _09231_ (.A1(net186),
    .A2(_02327_),
    .B1(_06417_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_2 _09232_ (.A(_06415_),
    .B(_06436_),
    .Y(_02329_));
 sky130_fd_sc_hd__or2_4 _09233_ (.A(_06415_),
    .B(_06436_),
    .X(_02330_));
 sky130_fd_sc_hd__and4bb_4 _09234_ (.A_N(instruction[4]),
    .B_N(instruction[6]),
    .C(instruction[5]),
    .D(instruction[3]),
    .X(_02331_));
 sky130_fd_sc_hd__or3b_4 _09235_ (.A(_06430_),
    .B(instruction[6]),
    .C_N(instruction[5]),
    .X(_02332_));
 sky130_fd_sc_hd__o21a_1 _09236_ (.A1(net233),
    .A2(_02331_),
    .B1(_06416_),
    .X(_02333_));
 sky130_fd_sc_hd__nor2_4 _09237_ (.A(_06436_),
    .B(_06451_),
    .Y(_02334_));
 sky130_fd_sc_hd__or2_1 _09238_ (.A(_06436_),
    .B(_06451_),
    .X(_02335_));
 sky130_fd_sc_hd__nor2_2 _09239_ (.A(_06428_),
    .B(_06436_),
    .Y(_02336_));
 sky130_fd_sc_hd__or2_2 _09240_ (.A(_06428_),
    .B(_06436_),
    .X(_02337_));
 sky130_fd_sc_hd__a221o_1 _09241_ (.A1(\div_res[0] ),
    .A2(_02334_),
    .B1(_02336_),
    .B2(\div_shifter[32] ),
    .C1(_02333_),
    .X(_02338_));
 sky130_fd_sc_hd__nor2_1 _09242_ (.A(_02328_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_2 _09243_ (.A(_04427_),
    .B(net196),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _09244_ (.A(_06318_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__or2_4 _09245_ (.A(_06318_),
    .B(_02340_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _09246_ (.A0(_02293_),
    .A1(_02340_),
    .S(net206),
    .X(_02343_));
 sky130_fd_sc_hd__o21a_1 _09247_ (.A1(_06336_),
    .A2(_02340_),
    .B1(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__or2_1 _09248_ (.A(_06330_),
    .B(_02340_),
    .X(_02345_));
 sky130_fd_sc_hd__and2_1 _09249_ (.A(_02344_),
    .B(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__or2_2 _09250_ (.A(net219),
    .B(_02340_),
    .X(_02347_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(_02346_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__or2_2 _09252_ (.A(_02341_),
    .B(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__o221a_1 _09253_ (.A1(_02314_),
    .A2(_02320_),
    .B1(_02349_),
    .B2(net168),
    .C1(_02339_),
    .X(_02350_));
 sky130_fd_sc_hd__o311a_1 _09254_ (.A1(instruction[5]),
    .A2(_06405_),
    .A3(_06428_),
    .B1(_02318_),
    .C1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__a31o_1 _09255_ (.A1(_02247_),
    .A2(_02248_),
    .A3(_02351_),
    .B1(_06463_),
    .X(_02352_));
 sky130_fd_sc_hd__a21o_1 _09256_ (.A1(_06462_),
    .A2(_02352_),
    .B1(net248),
    .X(_02353_));
 sky130_fd_sc_hd__o21ai_4 _09257_ (.A1(curr_PC[0]),
    .A2(net244),
    .B1(_02353_),
    .Y(dest_val[0]));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02354_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .Y(_02355_));
 sky130_fd_sc_hd__o21a_1 _09260_ (.A1(_02135_),
    .A2(_02243_),
    .B1(net161),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_4 _09261_ (.A1(_02141_),
    .A2(_02238_),
    .B1(_02237_),
    .Y(_02357_));
 sky130_fd_sc_hd__o21ai_4 _09262_ (.A1(_02232_),
    .A2(_02233_),
    .B1(_02235_),
    .Y(_02358_));
 sky130_fd_sc_hd__a32o_1 _09263_ (.A1(_02183_),
    .A2(_02184_),
    .A3(_02195_),
    .B1(_02196_),
    .B2(_02174_),
    .X(_02359_));
 sky130_fd_sc_hd__o22a_1 _09264_ (.A1(net130),
    .A2(net23),
    .B1(net15),
    .B2(net128),
    .X(_02360_));
 sky130_fd_sc_hd__xnor2_1 _09265_ (.A(net70),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__a22o_1 _09266_ (.A1(net37),
    .A2(_00293_),
    .B1(_00315_),
    .B2(net39),
    .X(_02362_));
 sky130_fd_sc_hd__xor2_1 _09267_ (.A(net91),
    .B(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__and2b_1 _09268_ (.A_N(_02361_),
    .B(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__and2b_1 _09269_ (.A_N(_02363_),
    .B(_02361_),
    .X(_02365_));
 sky130_fd_sc_hd__or2_1 _09270_ (.A(_02364_),
    .B(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__a22o_1 _09271_ (.A1(net43),
    .A2(net112),
    .B1(_00360_),
    .B2(net41),
    .X(_02367_));
 sky130_fd_sc_hd__xor2_1 _09272_ (.A(net94),
    .B(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__and2b_1 _09273_ (.A_N(_02366_),
    .B(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__and2b_1 _09274_ (.A_N(_02368_),
    .B(_02366_),
    .X(_02370_));
 sky130_fd_sc_hd__or2_1 _09275_ (.A(_02369_),
    .B(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__a21oi_1 _09276_ (.A1(_02160_),
    .A2(_02163_),
    .B1(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__and3_1 _09277_ (.A(_02160_),
    .B(_02163_),
    .C(_02371_),
    .X(_02373_));
 sky130_fd_sc_hd__nor2_1 _09278_ (.A(_02372_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__xnor2_1 _09279_ (.A(_02359_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__and2b_1 _09280_ (.A_N(_02179_),
    .B(_02183_),
    .X(_02376_));
 sky130_fd_sc_hd__a21o_1 _09281_ (.A1(_02214_),
    .A2(_02216_),
    .B1(_02213_),
    .X(_02377_));
 sky130_fd_sc_hd__a21o_1 _09282_ (.A1(_02170_),
    .A2(_02173_),
    .B1(_02169_),
    .X(_02378_));
 sky130_fd_sc_hd__xor2_1 _09283_ (.A(_02377_),
    .B(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__and2b_1 _09284_ (.A_N(_02376_),
    .B(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__xnor2_1 _09285_ (.A(_02376_),
    .B(_02379_),
    .Y(_02381_));
 sky130_fd_sc_hd__o22a_1 _09286_ (.A1(net55),
    .A2(net147),
    .B1(net145),
    .B2(net67),
    .X(_02382_));
 sky130_fd_sc_hd__xnor2_1 _09287_ (.A(net189),
    .B(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__o22a_1 _09288_ (.A1(net56),
    .A2(net105),
    .B1(net103),
    .B2(net62),
    .X(_02384_));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(net135),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_1 _09290_ (.A(_02383_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__xor2_1 _09291_ (.A(_02383_),
    .B(_02385_),
    .X(_02387_));
 sky130_fd_sc_hd__o22a_1 _09292_ (.A1(net64),
    .A2(net134),
    .B1(net132),
    .B2(net58),
    .X(_02388_));
 sky130_fd_sc_hd__xnor2_1 _09293_ (.A(net172),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__and2b_1 _09294_ (.A_N(_02389_),
    .B(_02387_),
    .X(_02390_));
 sky130_fd_sc_hd__and2b_1 _09295_ (.A_N(_02387_),
    .B(_02389_),
    .X(_02391_));
 sky130_fd_sc_hd__nor2_1 _09296_ (.A(_02390_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__o22a_1 _09297_ (.A1(net149),
    .A2(net11),
    .B1(net7),
    .B2(net151),
    .X(_02393_));
 sky130_fd_sc_hd__xor2_1 _09298_ (.A(net192),
    .B(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__a21o_1 _09299_ (.A1(_00687_),
    .A2(_00688_),
    .B1(net155),
    .X(_02395_));
 sky130_fd_sc_hd__or3_1 _09300_ (.A(net153),
    .B(_00395_),
    .C(_00397_),
    .X(_02396_));
 sky130_fd_sc_hd__nand3_1 _09301_ (.A(_06507_),
    .B(_02395_),
    .C(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__a21o_1 _09302_ (.A1(_02395_),
    .A2(_02396_),
    .B1(_06507_),
    .X(_02398_));
 sky130_fd_sc_hd__a21oi_1 _09303_ (.A1(_02397_),
    .A2(_02398_),
    .B1(net239),
    .Y(_02399_));
 sky130_fd_sc_hd__a21o_1 _09304_ (.A1(_02397_),
    .A2(_02398_),
    .B1(net239),
    .X(_02400_));
 sky130_fd_sc_hd__nand3_1 _09305_ (.A(net239),
    .B(_02397_),
    .C(_02398_),
    .Y(_02401_));
 sky130_fd_sc_hd__and3_1 _09306_ (.A(_02394_),
    .B(_02400_),
    .C(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__a21oi_1 _09307_ (.A1(_02400_),
    .A2(_02401_),
    .B1(_02394_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _09308_ (.A(_02402_),
    .B(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__o22a_1 _09309_ (.A1(net60),
    .A2(net85),
    .B1(net81),
    .B2(net52),
    .X(_02405_));
 sky130_fd_sc_hd__xnor2_1 _09310_ (.A(net137),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__o22a_1 _09311_ (.A1(net99),
    .A2(net34),
    .B1(net32),
    .B2(net84),
    .X(_02407_));
 sky130_fd_sc_hd__xnor2_1 _09312_ (.A(net124),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__or2_1 _09313_ (.A(_02406_),
    .B(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__nand2_1 _09314_ (.A(_02406_),
    .B(_02408_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _09315_ (.A(_02409_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__o22a_1 _09316_ (.A1(net50),
    .A2(net77),
    .B1(net73),
    .B2(net100),
    .X(_02412_));
 sky130_fd_sc_hd__xnor2_1 _09317_ (.A(net121),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__xor2_1 _09318_ (.A(_02411_),
    .B(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__nand2_1 _09319_ (.A(_02404_),
    .B(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__xor2_1 _09320_ (.A(_02404_),
    .B(_02414_),
    .X(_02416_));
 sky130_fd_sc_hd__and2_1 _09321_ (.A(_02392_),
    .B(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__inv_2 _09322_ (.A(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__xnor2_1 _09323_ (.A(_02392_),
    .B(_02416_),
    .Y(_02419_));
 sky130_fd_sc_hd__nor2_1 _09324_ (.A(net143),
    .B(net20),
    .Y(_02420_));
 sky130_fd_sc_hd__o22a_1 _09325_ (.A1(_00242_),
    .A2(net10),
    .B1(net5),
    .B2(_00249_),
    .X(_02421_));
 sky130_fd_sc_hd__xnor2_1 _09326_ (.A(net20),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21oi_1 _09327_ (.A1(_02191_),
    .A2(_02193_),
    .B1(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__a21o_1 _09328_ (.A1(_02191_),
    .A2(_02193_),
    .B1(_02422_),
    .X(_02424_));
 sky130_fd_sc_hd__and3_1 _09329_ (.A(_02191_),
    .B(_02193_),
    .C(_02422_),
    .X(_02425_));
 sky130_fd_sc_hd__nor2_1 _09330_ (.A(_02423_),
    .B(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__xnor2_2 _09331_ (.A(_02420_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__or2_1 _09332_ (.A(_02419_),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__nand2_1 _09333_ (.A(_02419_),
    .B(_02427_),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_1 _09334_ (.A(_02419_),
    .B(_02427_),
    .Y(_02430_));
 sky130_fd_sc_hd__xnor2_1 _09335_ (.A(_02381_),
    .B(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__a21o_1 _09336_ (.A1(_02145_),
    .A2(_02147_),
    .B1(_02151_),
    .X(_02432_));
 sky130_fd_sc_hd__o22a_1 _09337_ (.A1(net47),
    .A2(net117),
    .B1(net111),
    .B2(net45),
    .X(_02433_));
 sky130_fd_sc_hd__xnor2_1 _09338_ (.A(net97),
    .B(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__o22a_1 _09339_ (.A1(net27),
    .A2(net80),
    .B1(net76),
    .B2(net24),
    .X(_02435_));
 sky130_fd_sc_hd__xnor2_1 _09340_ (.A(_00286_),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__and2_1 _09341_ (.A(_02434_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__nor2_1 _09342_ (.A(_02434_),
    .B(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__nor2_1 _09343_ (.A(_02437_),
    .B(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__a22o_1 _09344_ (.A1(net118),
    .A2(net28),
    .B1(_00352_),
    .B2(net30),
    .X(_02440_));
 sky130_fd_sc_hd__xnor2_2 _09345_ (.A(net49),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__xnor2_2 _09346_ (.A(_02439_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21boi_2 _09347_ (.A1(_02198_),
    .A2(_02203_),
    .B1_N(_02202_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _09348_ (.A(_02442_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__xor2_2 _09349_ (.A(_02442_),
    .B(_02443_),
    .X(_02445_));
 sky130_fd_sc_hd__xor2_2 _09350_ (.A(_02432_),
    .B(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__xnor2_1 _09351_ (.A(_02431_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_1 _09352_ (.A(_02375_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__and2_1 _09353_ (.A(_02375_),
    .B(_02447_),
    .X(_02449_));
 sky130_fd_sc_hd__nor2_2 _09354_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__a21o_2 _09355_ (.A1(_02158_),
    .A2(_02223_),
    .B1(_02222_),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_02154_),
    .B(_02157_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21oi_2 _09357_ (.A1(_02164_),
    .A2(_02206_),
    .B1(_02205_),
    .Y(_02453_));
 sky130_fd_sc_hd__a21oi_2 _09358_ (.A1(_02208_),
    .A2(_02220_),
    .B1(_02219_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _09359_ (.A(_02453_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__xor2_2 _09360_ (.A(_02453_),
    .B(_02454_),
    .X(_02456_));
 sky130_fd_sc_hd__xnor2_2 _09361_ (.A(_02452_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__a21oi_2 _09362_ (.A1(_02227_),
    .A2(_02231_),
    .B1(_02230_),
    .Y(_02458_));
 sky130_fd_sc_hd__xnor2_2 _09363_ (.A(_02457_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2b_1 _09364_ (.A_N(_02459_),
    .B(_02451_),
    .Y(_02460_));
 sky130_fd_sc_hd__xnor2_4 _09365_ (.A(_02451_),
    .B(_02459_),
    .Y(_02461_));
 sky130_fd_sc_hd__and2_1 _09366_ (.A(_02450_),
    .B(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__xor2_4 _09367_ (.A(_02450_),
    .B(_02461_),
    .X(_02463_));
 sky130_fd_sc_hd__xnor2_4 _09368_ (.A(_02358_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__or2_1 _09369_ (.A(_02357_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__xnor2_4 _09370_ (.A(_02357_),
    .B(_02464_),
    .Y(_02466_));
 sky130_fd_sc_hd__and4_1 _09371_ (.A(_01800_),
    .B(_02129_),
    .C(_02132_),
    .D(_02241_),
    .X(_02467_));
 sky130_fd_sc_hd__a2bb2o_1 _09372_ (.A1_N(_02239_),
    .A2_N(_02140_),
    .B1(_02127_),
    .B2(_02020_),
    .X(_02468_));
 sky130_fd_sc_hd__a32o_1 _09373_ (.A1(_02129_),
    .A2(_02131_),
    .A3(_02241_),
    .B1(_02468_),
    .B2(_02240_),
    .X(_02469_));
 sky130_fd_sc_hd__or2_2 _09374_ (.A(_02467_),
    .B(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__xnor2_2 _09375_ (.A(_02466_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__o21ai_1 _09376_ (.A1(_02356_),
    .A2(_02471_),
    .B1(_02245_),
    .Y(_02472_));
 sky130_fd_sc_hd__a21oi_1 _09377_ (.A1(_02356_),
    .A2(_02471_),
    .B1(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(_02251_),
    .A1(_02254_),
    .S(net205),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(_02255_),
    .A1(_02258_),
    .S(net207),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _09380_ (.A0(_02474_),
    .A1(_02475_),
    .S(net211),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(_02259_),
    .A1(_02261_),
    .S(net207),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(_02262_),
    .A1(_02266_),
    .S(net207),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(_02477_),
    .A1(_02478_),
    .S(net211),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(_02476_),
    .A1(_02479_),
    .S(net214),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(_02267_),
    .A1(_02269_),
    .S(net207),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(_02270_),
    .A1(_02273_),
    .S(net205),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(_02481_),
    .A1(_02482_),
    .S(net211),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(_02274_),
    .A1(_02276_),
    .S(net205),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(_02277_),
    .A1(_02297_),
    .S(net205),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(_02484_),
    .A1(_02485_),
    .S(net211),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_02483_),
    .A1(_02486_),
    .S(net214),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(_02480_),
    .A1(_02487_),
    .S(net217),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(_02283_),
    .A1(_02285_),
    .S(net205),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _09394_ (.A0(_02286_),
    .A1(_02289_),
    .S(net206),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(_02489_),
    .A1(_02490_),
    .S(net212),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(_02290_),
    .A1(_02292_),
    .S(net206),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _09397_ (.A0(_02343_),
    .A1(_02492_),
    .S(_06336_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(_02491_),
    .A1(_02493_),
    .S(net215),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(_02298_),
    .A1(_02300_),
    .S(net205),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _09400_ (.A0(_02301_),
    .A1(_02304_),
    .S(net205),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(_02495_),
    .A1(_02496_),
    .S(net211),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(_02305_),
    .A1(_02307_),
    .S(net205),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _09403_ (.A0(_02282_),
    .A1(_02308_),
    .S(net209),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(_02498_),
    .A1(_02499_),
    .S(net212),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _09405_ (.A0(_02497_),
    .A1(_02500_),
    .S(net214),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(_02494_),
    .A1(_02501_),
    .S(net219),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_2 _09407_ (.A0(_02488_),
    .A1(_02502_),
    .S(net220),
    .X(_02503_));
 sky130_fd_sc_hd__inv_2 _09408_ (.A(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__and2_1 _09409_ (.A(net289),
    .B(curr_PC[1]),
    .X(_02505_));
 sky130_fd_sc_hd__xor2_1 _09410_ (.A(net289),
    .B(curr_PC[1]),
    .X(_02506_));
 sky130_fd_sc_hd__xnor2_1 _09411_ (.A(_02315_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__o21a_1 _09412_ (.A1(net223),
    .A2(_02507_),
    .B1(net197),
    .X(_02508_));
 sky130_fd_sc_hd__o21a_1 _09413_ (.A1(_02319_),
    .A2(_02508_),
    .B1(_02503_),
    .X(_02509_));
 sky130_fd_sc_hd__a21oi_1 _09414_ (.A1(\div_res[0] ),
    .A2(_06464_),
    .B1(\div_res[1] ),
    .Y(_02510_));
 sky130_fd_sc_hd__a311o_1 _09415_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(_06464_),
    .B1(net183),
    .C1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__xnor2_1 _09416_ (.A(_06339_),
    .B(_06343_),
    .Y(_02512_));
 sky130_fd_sc_hd__o21ai_1 _09417_ (.A1(net294),
    .A2(net210),
    .B1(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__or3_1 _09418_ (.A(net294),
    .B(net210),
    .C(_02512_),
    .X(_02514_));
 sky130_fd_sc_hd__nor2_1 _09419_ (.A(_06339_),
    .B(net234),
    .Y(_02515_));
 sky130_fd_sc_hd__and2_1 _09420_ (.A(divi1_sign),
    .B(instruction[7]),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_1 _09421_ (.A1(\div_shifter[32] ),
    .A2(net230),
    .B1(\div_shifter[33] ),
    .Y(_02517_));
 sky130_fd_sc_hd__a31o_1 _09422_ (.A1(\div_shifter[33] ),
    .A2(\div_shifter[32] ),
    .A3(net230),
    .B1(_02337_),
    .X(_02518_));
 sky130_fd_sc_hd__a2bb2o_1 _09423_ (.A1_N(_02518_),
    .A2_N(_02517_),
    .B1(_06460_),
    .B2(net213),
    .X(_02519_));
 sky130_fd_sc_hd__a31o_1 _09424_ (.A1(reg1_val[1]),
    .A2(net213),
    .A3(_02331_),
    .B1(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a221o_1 _09425_ (.A1(_06338_),
    .A2(_02321_),
    .B1(_02508_),
    .B2(net250),
    .C1(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__a311o_1 _09426_ (.A1(_02323_),
    .A2(_02513_),
    .A3(_02514_),
    .B1(_02515_),
    .C1(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__or3b_1 _09427_ (.A(_02509_),
    .B(_02522_),
    .C_N(_02511_),
    .X(_02523_));
 sky130_fd_sc_hd__o21ai_1 _09428_ (.A1(net156),
    .A2(net239),
    .B1(_06416_),
    .Y(_02524_));
 sky130_fd_sc_hd__a21o_1 _09429_ (.A1(net156),
    .A2(net239),
    .B1(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__xnor2_1 _09430_ (.A(_01751_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__mux2_1 _09431_ (.A0(_02294_),
    .A1(_02340_),
    .S(net212),
    .X(_02527_));
 sky130_fd_sc_hd__o21a_1 _09432_ (.A1(net215),
    .A2(_02527_),
    .B1(_02345_),
    .X(_02528_));
 sky130_fd_sc_hd__o21a_1 _09433_ (.A1(net217),
    .A2(_02528_),
    .B1(_02347_),
    .X(_02529_));
 sky130_fd_sc_hd__o21ai_2 _09434_ (.A1(net221),
    .A2(_02529_),
    .B1(_02342_),
    .Y(_02530_));
 sky130_fd_sc_hd__a2bb2o_1 _09435_ (.A1_N(net167),
    .A2_N(_02530_),
    .B1(_02526_),
    .B2(net233),
    .X(_02531_));
 sky130_fd_sc_hd__o31a_1 _09436_ (.A1(_02473_),
    .A2(_02523_),
    .A3(_02531_),
    .B1(net245),
    .X(_02532_));
 sky130_fd_sc_hd__a31o_4 _09437_ (.A1(net248),
    .A2(_02354_),
    .A3(_02355_),
    .B1(_02532_),
    .X(dest_val[1]));
 sky130_fd_sc_hd__nand3_1 _09438_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .Y(_02533_));
 sky130_fd_sc_hd__a21o_1 _09439_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .X(_02534_));
 sky130_fd_sc_hd__or3_2 _09440_ (.A(_02135_),
    .B(_02243_),
    .C(_02471_),
    .X(_02535_));
 sky130_fd_sc_hd__a21oi_4 _09441_ (.A1(_02358_),
    .A2(_02463_),
    .B1(_02462_),
    .Y(_02536_));
 sky130_fd_sc_hd__o21ai_4 _09442_ (.A1(_02457_),
    .A2(_02458_),
    .B1(_02460_),
    .Y(_02537_));
 sky130_fd_sc_hd__o22a_1 _09443_ (.A1(_00361_),
    .A2(net23),
    .B1(net15),
    .B2(net130),
    .X(_02538_));
 sky130_fd_sc_hd__xnor2_1 _09444_ (.A(net70),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__a22o_1 _09445_ (.A1(net39),
    .A2(_00309_),
    .B1(_00315_),
    .B2(net37),
    .X(_02540_));
 sky130_fd_sc_hd__xor2_1 _09446_ (.A(net91),
    .B(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__and2b_1 _09447_ (.A_N(_02539_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__and2b_1 _09448_ (.A_N(_02541_),
    .B(_02539_),
    .X(_02543_));
 sky130_fd_sc_hd__or2_1 _09449_ (.A(_02542_),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__a22o_1 _09450_ (.A1(net43),
    .A2(_00293_),
    .B1(net112),
    .B2(net41),
    .X(_02545_));
 sky130_fd_sc_hd__xor2_1 _09451_ (.A(net94),
    .B(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__and2b_1 _09452_ (.A_N(_02544_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__and2b_1 _09453_ (.A_N(_02546_),
    .B(_02544_),
    .X(_02548_));
 sky130_fd_sc_hd__or2_2 _09454_ (.A(_02547_),
    .B(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__a21oi_2 _09455_ (.A1(_02377_),
    .A2(_02378_),
    .B1(_02380_),
    .Y(_02550_));
 sky130_fd_sc_hd__xnor2_1 _09456_ (.A(_02549_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__a21o_1 _09457_ (.A1(_02415_),
    .A2(_02418_),
    .B1(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__nand3_1 _09458_ (.A(_02415_),
    .B(_02418_),
    .C(_02551_),
    .Y(_02553_));
 sky130_fd_sc_hd__and2_2 _09459_ (.A(_02552_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__o21a_1 _09460_ (.A1(_02411_),
    .A2(_02413_),
    .B1(_02409_),
    .X(_02555_));
 sky130_fd_sc_hd__a21o_1 _09461_ (.A1(_02439_),
    .A2(_02441_),
    .B1(_02437_),
    .X(_02556_));
 sky130_fd_sc_hd__nor2_1 _09462_ (.A(_02386_),
    .B(_02390_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21ai_1 _09463_ (.A1(_02386_),
    .A2(_02390_),
    .B1(_02556_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_1 _09464_ (.A(_02556_),
    .B(_02557_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2b_1 _09465_ (.A_N(_02555_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__xnor2_1 _09466_ (.A(_02555_),
    .B(_02559_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _09467_ (.A(_00249_),
    .B(net20),
    .Y(_02562_));
 sky130_fd_sc_hd__o22a_1 _09468_ (.A1(net128),
    .A2(net10),
    .B1(net5),
    .B2(net141),
    .X(_02563_));
 sky130_fd_sc_hd__xnor2_1 _09469_ (.A(net21),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__o21a_1 _09470_ (.A1(_02399_),
    .A2(_02402_),
    .B1(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__or3_1 _09471_ (.A(_02399_),
    .B(_02402_),
    .C(_02564_),
    .X(_02566_));
 sky130_fd_sc_hd__and2b_1 _09472_ (.A_N(_02565_),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__xnor2_1 _09473_ (.A(_02562_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o22a_1 _09474_ (.A1(net58),
    .A2(net105),
    .B1(net103),
    .B2(net56),
    .X(_02569_));
 sky130_fd_sc_hd__xnor2_1 _09475_ (.A(net135),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__o22a_1 _09476_ (.A1(net55),
    .A2(net145),
    .B1(net16),
    .B2(net147),
    .X(_02571_));
 sky130_fd_sc_hd__xnor2_1 _09477_ (.A(net189),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__and2_1 _09479_ (.A(_02570_),
    .B(_02572_),
    .X(_02574_));
 sky130_fd_sc_hd__nor2_1 _09480_ (.A(_02573_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__o22a_1 _09481_ (.A1(net67),
    .A2(net134),
    .B1(net132),
    .B2(net64),
    .X(_02576_));
 sky130_fd_sc_hd__xnor2_1 _09482_ (.A(net173),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_1 _09483_ (.A(_02575_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__o22a_1 _09484_ (.A1(net62),
    .A2(net85),
    .B1(net81),
    .B2(net60),
    .X(_02579_));
 sky130_fd_sc_hd__xnor2_1 _09485_ (.A(net137),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__o22a_1 _09486_ (.A1(net100),
    .A2(net34),
    .B1(net32),
    .B2(net98),
    .X(_02581_));
 sky130_fd_sc_hd__xnor2_1 _09487_ (.A(net124),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__or2_1 _09488_ (.A(_02580_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(_02580_),
    .B(_02582_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _09490_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o22a_1 _09491_ (.A1(net52),
    .A2(net77),
    .B1(net73),
    .B2(net50),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_1 _09492_ (.A(net121),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__xnor2_1 _09493_ (.A(_02585_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__o22a_1 _09494_ (.A1(net153),
    .A2(net13),
    .B1(net11),
    .B2(_06513_),
    .X(_02589_));
 sky130_fd_sc_hd__xnor2_2 _09495_ (.A(net194),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nor2_1 _09496_ (.A(net239),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__xnor2_2 _09497_ (.A(_06468_),
    .B(_02590_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _09498_ (.A1(_06540_),
    .A2(net8),
    .B1(net192),
    .Y(_02593_));
 sky130_fd_sc_hd__a31o_2 _09499_ (.A1(net192),
    .A2(_06530_),
    .A3(net8),
    .B1(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__xnor2_2 _09500_ (.A(_02592_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nor2_1 _09501_ (.A(_02588_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__xor2_1 _09502_ (.A(_02588_),
    .B(_02595_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _09503_ (.A(_02578_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__nor2_1 _09504_ (.A(_02568_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__xor2_1 _09505_ (.A(_02568_),
    .B(_02598_),
    .X(_02600_));
 sky130_fd_sc_hd__xor2_1 _09506_ (.A(_02561_),
    .B(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__nor2_1 _09507_ (.A(_02364_),
    .B(_02369_),
    .Y(_02602_));
 sky130_fd_sc_hd__o22a_1 _09508_ (.A1(net26),
    .A2(net84),
    .B1(net80),
    .B2(net24),
    .X(_02603_));
 sky130_fd_sc_hd__xnor2_1 _09509_ (.A(net87),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__o22a_1 _09510_ (.A1(net47),
    .A2(net120),
    .B1(net117),
    .B2(net45),
    .X(_02605_));
 sky130_fd_sc_hd__xnor2_1 _09511_ (.A(net97),
    .B(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__and2_1 _09512_ (.A(_02604_),
    .B(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__nor2_1 _09513_ (.A(_02604_),
    .B(_02606_),
    .Y(_02608_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__a22o_1 _09515_ (.A1(net30),
    .A2(_00347_),
    .B1(_00352_),
    .B2(net28),
    .X(_02610_));
 sky130_fd_sc_hd__xnor2_2 _09516_ (.A(net48),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__xnor2_2 _09517_ (.A(_02609_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__o31a_1 _09518_ (.A1(net143),
    .A2(net20),
    .A3(_02425_),
    .B1(_02424_),
    .X(_02613_));
 sky130_fd_sc_hd__nor2_1 _09519_ (.A(_02612_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__xor2_1 _09520_ (.A(_02612_),
    .B(_02613_),
    .X(_02615_));
 sky130_fd_sc_hd__and2b_1 _09521_ (.A_N(_02602_),
    .B(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__xnor2_1 _09522_ (.A(_02602_),
    .B(_02615_),
    .Y(_02617_));
 sky130_fd_sc_hd__and2_1 _09523_ (.A(_02601_),
    .B(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__nor2_1 _09524_ (.A(_02601_),
    .B(_02617_),
    .Y(_02619_));
 sky130_fd_sc_hd__nor2_2 _09525_ (.A(_02618_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__xor2_4 _09526_ (.A(_02554_),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__a21o_2 _09527_ (.A1(_02431_),
    .A2(_02446_),
    .B1(_02448_),
    .X(_02622_));
 sky130_fd_sc_hd__a21o_1 _09528_ (.A1(_02452_),
    .A2(_02456_),
    .B1(_02455_),
    .X(_02623_));
 sky130_fd_sc_hd__a21o_1 _09529_ (.A1(_02359_),
    .A2(_02374_),
    .B1(_02372_),
    .X(_02624_));
 sky130_fd_sc_hd__a21bo_1 _09530_ (.A1(_02381_),
    .A2(_02429_),
    .B1_N(_02428_),
    .X(_02625_));
 sky130_fd_sc_hd__a21o_1 _09531_ (.A1(_02432_),
    .A2(_02445_),
    .B1(_02444_),
    .X(_02626_));
 sky130_fd_sc_hd__and2_1 _09532_ (.A(_02625_),
    .B(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__xor2_2 _09533_ (.A(_02625_),
    .B(_02626_),
    .X(_02628_));
 sky130_fd_sc_hd__xor2_2 _09534_ (.A(_02624_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__xnor2_2 _09535_ (.A(_02623_),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2b_1 _09536_ (.A_N(_02630_),
    .B(_02622_),
    .Y(_02631_));
 sky130_fd_sc_hd__xnor2_4 _09537_ (.A(_02622_),
    .B(_02630_),
    .Y(_02632_));
 sky130_fd_sc_hd__and2_1 _09538_ (.A(_02621_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__xor2_4 _09539_ (.A(_02621_),
    .B(_02632_),
    .X(_02634_));
 sky130_fd_sc_hd__xnor2_4 _09540_ (.A(_02537_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__or2_1 _09541_ (.A(_02536_),
    .B(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__and2_1 _09542_ (.A(_02536_),
    .B(_02635_),
    .X(_02637_));
 sky130_fd_sc_hd__xnor2_4 _09543_ (.A(_02536_),
    .B(_02635_),
    .Y(_02638_));
 sky130_fd_sc_hd__or4_1 _09544_ (.A(_02012_),
    .B(_02130_),
    .C(_02242_),
    .D(_02466_),
    .X(_02639_));
 sky130_fd_sc_hd__o22a_1 _09545_ (.A1(_02140_),
    .A2(_02239_),
    .B1(_02357_),
    .B2(_02464_),
    .X(_02640_));
 sky130_fd_sc_hd__a21o_1 _09546_ (.A1(_02357_),
    .A2(_02464_),
    .B1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__or4_1 _09547_ (.A(_02128_),
    .B(_02137_),
    .C(_02242_),
    .D(_02466_),
    .X(_02642_));
 sky130_fd_sc_hd__o211a_2 _09548_ (.A1(_02017_),
    .A2(_02639_),
    .B1(_02641_),
    .C1(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__xor2_4 _09549_ (.A(_02638_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__a21oi_1 _09550_ (.A1(net162),
    .A2(_02535_),
    .B1(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__a31o_1 _09551_ (.A1(net162),
    .A2(_02535_),
    .A3(_02644_),
    .B1(net187),
    .X(_02646_));
 sky130_fd_sc_hd__nor2_1 _09552_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _09553_ (.A(net161),
    .B(_01752_),
    .Y(_02648_));
 sky130_fd_sc_hd__mux2_1 _09554_ (.A0(_01750_),
    .A1(_01804_),
    .S(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__o21ai_1 _09555_ (.A1(net216),
    .A2(_02493_),
    .B1(_02345_),
    .Y(_02650_));
 sky130_fd_sc_hd__inv_2 _09556_ (.A(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__o21a_1 _09557_ (.A1(net218),
    .A2(_02651_),
    .B1(_02347_),
    .X(_02652_));
 sky130_fd_sc_hd__o21ai_2 _09558_ (.A1(net221),
    .A2(_02652_),
    .B1(_02342_),
    .Y(_02653_));
 sky130_fd_sc_hd__inv_2 _09559_ (.A(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__nor2_1 _09560_ (.A(net167),
    .B(_02653_),
    .Y(_02655_));
 sky130_fd_sc_hd__mux2_1 _09561_ (.A0(_02256_),
    .A1(_02260_),
    .S(net212),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _09562_ (.A0(_02263_),
    .A1(_02268_),
    .S(net211),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(_02656_),
    .A1(_02657_),
    .S(net215),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_02271_),
    .A1(_02275_),
    .S(net211),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(_02278_),
    .A1(_02299_),
    .S(net211),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _09566_ (.A0(_02659_),
    .A1(_02660_),
    .S(net215),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(_02658_),
    .A1(_02661_),
    .S(net217),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(_02287_),
    .A1(_02291_),
    .S(net212),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(_02527_),
    .A1(_02663_),
    .S(_06330_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(_02302_),
    .A1(_02306_),
    .S(net212),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(_02284_),
    .A1(_02309_),
    .S(_06336_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(_02665_),
    .A1(_02666_),
    .S(net214),
    .X(_02667_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(_02664_),
    .A1(_02667_),
    .S(net219),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(_02662_),
    .A1(_02668_),
    .S(net220),
    .X(_02669_));
 sky130_fd_sc_hd__a31oi_2 _09575_ (.A1(net293),
    .A2(curr_PC[0]),
    .A3(_02506_),
    .B1(_02505_),
    .Y(_02670_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02671_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2b_1 _09578_ (.A_N(_02671_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__xnor2_1 _09579_ (.A(_02670_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21o_1 _09580_ (.A1(net251),
    .A2(_02674_),
    .B1(net196),
    .X(_02675_));
 sky130_fd_sc_hd__a21boi_1 _09581_ (.A1(_02320_),
    .A2(_02675_),
    .B1_N(_02669_),
    .Y(_02676_));
 sky130_fd_sc_hd__or2_1 _09582_ (.A(\div_res[1] ),
    .B(\div_res[0] ),
    .X(_02677_));
 sky130_fd_sc_hd__a21oi_1 _09583_ (.A1(net160),
    .A2(_02677_),
    .B1(\div_res[2] ),
    .Y(_02678_));
 sky130_fd_sc_hd__a31o_1 _09584_ (.A1(\div_res[2] ),
    .A2(net160),
    .A3(_02677_),
    .B1(net183),
    .X(_02679_));
 sky130_fd_sc_hd__a22o_1 _09585_ (.A1(net289),
    .A2(net212),
    .B1(net206),
    .B2(net293),
    .X(_02680_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_06338_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(_06345_),
    .A1(_02681_),
    .S(net285),
    .X(_02682_));
 sky130_fd_sc_hd__a21oi_1 _09588_ (.A1(_06334_),
    .A2(_02682_),
    .B1(net236),
    .Y(_02683_));
 sky130_fd_sc_hd__o21ai_1 _09589_ (.A1(_06334_),
    .A2(_02682_),
    .B1(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__or2_1 _09590_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .X(_02685_));
 sky130_fd_sc_hd__a21oi_1 _09591_ (.A1(net230),
    .A2(_02685_),
    .B1(\div_shifter[34] ),
    .Y(_02686_));
 sky130_fd_sc_hd__a31o_1 _09592_ (.A1(\div_shifter[34] ),
    .A2(net230),
    .A3(_02685_),
    .B1(_02337_),
    .X(_02687_));
 sky130_fd_sc_hd__or2_1 _09593_ (.A(_02686_),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o221a_1 _09594_ (.A1(_06330_),
    .A2(net241),
    .B1(net185),
    .B2(_06332_),
    .C1(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__nand2_1 _09595_ (.A(_06333_),
    .B(_02321_),
    .Y(_02690_));
 sky130_fd_sc_hd__or2_1 _09596_ (.A(net224),
    .B(_02675_),
    .X(_02691_));
 sky130_fd_sc_hd__o2111a_1 _09597_ (.A1(_06334_),
    .A2(net234),
    .B1(_02689_),
    .C1(_02690_),
    .D1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__o211a_1 _09598_ (.A1(_02678_),
    .A2(_02679_),
    .B1(_02684_),
    .C1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__or3b_1 _09599_ (.A(_02655_),
    .B(_02676_),
    .C_N(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__a21o_1 _09600_ (.A1(net233),
    .A2(_02649_),
    .B1(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__o21a_1 _09601_ (.A1(_02647_),
    .A2(_02695_),
    .B1(net245),
    .X(_02696_));
 sky130_fd_sc_hd__a31o_4 _09602_ (.A1(net248),
    .A2(_02533_),
    .A3(_02534_),
    .B1(_02696_),
    .X(dest_val[2]));
 sky130_fd_sc_hd__o21ai_1 _09603_ (.A1(_02535_),
    .A2(_02644_),
    .B1(net161),
    .Y(_02697_));
 sky130_fd_sc_hd__a21oi_4 _09604_ (.A1(_02537_),
    .A2(_02634_),
    .B1(_02633_),
    .Y(_02698_));
 sky130_fd_sc_hd__a21bo_2 _09605_ (.A1(_02623_),
    .A2(_02629_),
    .B1_N(_02631_),
    .X(_02699_));
 sky130_fd_sc_hd__a21o_2 _09606_ (.A1(_02578_),
    .A2(_02597_),
    .B1(_02596_),
    .X(_02700_));
 sky130_fd_sc_hd__o22a_1 _09607_ (.A1(_00298_),
    .A2(net23),
    .B1(net15),
    .B2(_00361_),
    .X(_02701_));
 sky130_fd_sc_hd__xnor2_1 _09608_ (.A(net70),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__inv_2 _09609_ (.A(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__a22o_1 _09610_ (.A1(net39),
    .A2(net115),
    .B1(_00309_),
    .B2(net37),
    .X(_02704_));
 sky130_fd_sc_hd__xor2_1 _09611_ (.A(net91),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__xor2_1 _09612_ (.A(_02702_),
    .B(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _09613_ (.A1(net41),
    .A2(_00293_),
    .B1(_00315_),
    .B2(net43),
    .X(_02707_));
 sky130_fd_sc_hd__xor2_1 _09614_ (.A(net94),
    .B(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__and2b_1 _09615_ (.A_N(_02706_),
    .B(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__and2b_1 _09616_ (.A_N(_02708_),
    .B(_02706_),
    .X(_02710_));
 sky130_fd_sc_hd__or2_1 _09617_ (.A(_02709_),
    .B(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__a21oi_1 _09618_ (.A1(_02558_),
    .A2(_02560_),
    .B1(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__and3_1 _09619_ (.A(_02558_),
    .B(_02560_),
    .C(_02711_),
    .X(_02713_));
 sky130_fd_sc_hd__nor2_2 _09620_ (.A(_02712_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__xor2_4 _09621_ (.A(_02700_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__or2_1 _09622_ (.A(_02542_),
    .B(_02547_),
    .X(_02716_));
 sky130_fd_sc_hd__o22a_1 _09623_ (.A1(net99),
    .A2(net27),
    .B1(net25),
    .B2(net83),
    .X(_02717_));
 sky130_fd_sc_hd__xnor2_1 _09624_ (.A(_00286_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__o22a_1 _09625_ (.A1(net45),
    .A2(net120),
    .B1(net71),
    .B2(net47),
    .X(_02719_));
 sky130_fd_sc_hd__xnor2_1 _09626_ (.A(net97),
    .B(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__and2_1 _09627_ (.A(_02718_),
    .B(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__xor2_1 _09628_ (.A(_02718_),
    .B(_02720_),
    .X(_02722_));
 sky130_fd_sc_hd__a22o_1 _09629_ (.A1(net30),
    .A2(_00340_),
    .B1(_00347_),
    .B2(net28),
    .X(_02723_));
 sky130_fd_sc_hd__xnor2_1 _09630_ (.A(net48),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__xnor2_1 _09631_ (.A(_02722_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__a21o_1 _09632_ (.A1(_02562_),
    .A2(_02566_),
    .B1(_02565_),
    .X(_02726_));
 sky130_fd_sc_hd__nand2b_1 _09633_ (.A_N(_02725_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__xnor2_1 _09634_ (.A(_02725_),
    .B(_02726_),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_02716_),
    .B(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__or2_1 _09636_ (.A(_02716_),
    .B(_02728_),
    .X(_02730_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_02729_),
    .B(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__o21a_1 _09638_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02583_),
    .X(_02732_));
 sky130_fd_sc_hd__o21bai_2 _09639_ (.A1(_02574_),
    .A2(_02577_),
    .B1_N(_02573_),
    .Y(_02733_));
 sky130_fd_sc_hd__a21o_1 _09640_ (.A1(_02609_),
    .A2(_02611_),
    .B1(_02607_),
    .X(_02734_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__xor2_2 _09642_ (.A(_02733_),
    .B(_02734_),
    .X(_02736_));
 sky130_fd_sc_hd__nand2b_1 _09643_ (.A_N(_02732_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__xnor2_2 _09644_ (.A(_02732_),
    .B(_02736_),
    .Y(_02738_));
 sky130_fd_sc_hd__o22a_1 _09645_ (.A1(net64),
    .A2(net105),
    .B1(net103),
    .B2(net58),
    .X(_02739_));
 sky130_fd_sc_hd__xnor2_1 _09646_ (.A(_00328_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__a21o_1 _09647_ (.A1(_00687_),
    .A2(_00688_),
    .B1(net147),
    .X(_02741_));
 sky130_fd_sc_hd__or3_1 _09648_ (.A(net145),
    .B(_00395_),
    .C(_00397_),
    .X(_02742_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(_02741_),
    .A2(_02742_),
    .B1(net189),
    .X(_02743_));
 sky130_fd_sc_hd__nand3_1 _09650_ (.A(net189),
    .B(_02741_),
    .C(_02742_),
    .Y(_02744_));
 sky130_fd_sc_hd__and3_1 _09651_ (.A(_02740_),
    .B(_02743_),
    .C(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__a21oi_1 _09652_ (.A1(_02743_),
    .A2(_02744_),
    .B1(_02740_),
    .Y(_02746_));
 sky130_fd_sc_hd__nor2_1 _09653_ (.A(_02745_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__o22a_1 _09654_ (.A1(net55),
    .A2(net134),
    .B1(net132),
    .B2(net67),
    .X(_02748_));
 sky130_fd_sc_hd__xnor2_2 _09655_ (.A(net172),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__xnor2_2 _09656_ (.A(_02747_),
    .B(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__o22a_1 _09657_ (.A1(net57),
    .A2(net85),
    .B1(net81),
    .B2(net62),
    .X(_02751_));
 sky130_fd_sc_hd__xnor2_1 _09658_ (.A(_00323_),
    .B(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__o22a_1 _09659_ (.A1(net50),
    .A2(net34),
    .B1(net33),
    .B2(net100),
    .X(_02753_));
 sky130_fd_sc_hd__xnor2_1 _09660_ (.A(net124),
    .B(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__or2_1 _09661_ (.A(_02752_),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__nand2_1 _09662_ (.A(_02752_),
    .B(_02754_),
    .Y(_02756_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_02755_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__o22a_1 _09664_ (.A1(net60),
    .A2(net77),
    .B1(net73),
    .B2(net52),
    .X(_02758_));
 sky130_fd_sc_hd__xnor2_2 _09665_ (.A(net122),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__xnor2_2 _09666_ (.A(_02757_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__o22a_1 _09667_ (.A1(net153),
    .A2(net11),
    .B1(net7),
    .B2(net155),
    .X(_02761_));
 sky130_fd_sc_hd__xnor2_2 _09668_ (.A(net194),
    .B(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__nor2_1 _09669_ (.A(_06468_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__xnor2_2 _09670_ (.A(net239),
    .B(_02762_),
    .Y(_02764_));
 sky130_fd_sc_hd__xnor2_2 _09671_ (.A(net192),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _09672_ (.A(_02760_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__xor2_2 _09673_ (.A(_02760_),
    .B(_02765_),
    .X(_02767_));
 sky130_fd_sc_hd__xnor2_2 _09674_ (.A(_02750_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__nor2_1 _09675_ (.A(_00242_),
    .B(net20),
    .Y(_02769_));
 sky130_fd_sc_hd__a21oi_2 _09676_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02591_),
    .Y(_02770_));
 sky130_fd_sc_hd__o22a_1 _09677_ (.A1(net130),
    .A2(net10),
    .B1(net5),
    .B2(net128),
    .X(_02771_));
 sky130_fd_sc_hd__xnor2_2 _09678_ (.A(net21),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2b_1 _09679_ (.A_N(_02770_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__xnor2_2 _09680_ (.A(_02770_),
    .B(_02772_),
    .Y(_02774_));
 sky130_fd_sc_hd__xnor2_2 _09681_ (.A(_02769_),
    .B(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_1 _09682_ (.A(_02768_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__xor2_2 _09683_ (.A(_02768_),
    .B(_02775_),
    .X(_02777_));
 sky130_fd_sc_hd__xnor2_1 _09684_ (.A(_02738_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nor2_1 _09685_ (.A(_02731_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_1 _09686_ (.A(_02731_),
    .B(_02778_),
    .Y(_02780_));
 sky130_fd_sc_hd__and2b_1 _09687_ (.A_N(_02779_),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__xor2_4 _09688_ (.A(_02715_),
    .B(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__a21o_1 _09689_ (.A1(_02554_),
    .A2(_02620_),
    .B1(_02618_),
    .X(_02783_));
 sky130_fd_sc_hd__o21ai_4 _09690_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02552_),
    .Y(_02784_));
 sky130_fd_sc_hd__a21o_2 _09691_ (.A1(_02561_),
    .A2(_02600_),
    .B1(_02599_),
    .X(_02785_));
 sky130_fd_sc_hd__nor2_2 _09692_ (.A(_02614_),
    .B(_02616_),
    .Y(_02786_));
 sky130_fd_sc_hd__o21ai_1 _09693_ (.A1(_02614_),
    .A2(_02616_),
    .B1(_02785_),
    .Y(_02787_));
 sky130_fd_sc_hd__xnor2_4 _09694_ (.A(_02785_),
    .B(_02786_),
    .Y(_02788_));
 sky130_fd_sc_hd__xnor2_4 _09695_ (.A(_02784_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__a21oi_2 _09696_ (.A1(_02624_),
    .A2(_02628_),
    .B1(_02627_),
    .Y(_02790_));
 sky130_fd_sc_hd__xnor2_2 _09697_ (.A(_02789_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2b_1 _09698_ (.A_N(_02791_),
    .B(_02783_),
    .Y(_02792_));
 sky130_fd_sc_hd__xnor2_2 _09699_ (.A(_02783_),
    .B(_02791_),
    .Y(_02793_));
 sky130_fd_sc_hd__and2_1 _09700_ (.A(_02782_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__xor2_4 _09701_ (.A(_02782_),
    .B(_02793_),
    .X(_02795_));
 sky130_fd_sc_hd__xnor2_4 _09702_ (.A(_02699_),
    .B(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__or2_1 _09703_ (.A(_02698_),
    .B(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__and2_1 _09704_ (.A(_02698_),
    .B(_02796_),
    .X(_02798_));
 sky130_fd_sc_hd__xnor2_4 _09705_ (.A(_02698_),
    .B(_02796_),
    .Y(_02799_));
 sky130_fd_sc_hd__or4_1 _09706_ (.A(_02130_),
    .B(_02242_),
    .C(_02466_),
    .D(_02638_),
    .X(_02800_));
 sky130_fd_sc_hd__a21o_1 _09707_ (.A1(_02465_),
    .A2(_02636_),
    .B1(_02637_),
    .X(_02801_));
 sky130_fd_sc_hd__or4bb_1 _09708_ (.A(_02466_),
    .B(_02638_),
    .C_N(_02468_),
    .D_N(_02240_),
    .X(_02802_));
 sky130_fd_sc_hd__o211a_2 _09709_ (.A1(_02133_),
    .A2(_02800_),
    .B1(_02801_),
    .C1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__xnor2_2 _09710_ (.A(_02799_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__a21oi_1 _09711_ (.A1(_02697_),
    .A2(_02804_),
    .B1(net187),
    .Y(_02805_));
 sky130_fd_sc_hd__o21a_1 _09712_ (.A1(_02697_),
    .A2(_02804_),
    .B1(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__o21ai_1 _09713_ (.A1(net156),
    .A2(_01805_),
    .B1(_01807_),
    .Y(_02807_));
 sky130_fd_sc_hd__or3_1 _09714_ (.A(net156),
    .B(_01805_),
    .C(_01807_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(_02475_),
    .A1(_02477_),
    .S(net211),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _09716_ (.A0(_02478_),
    .A1(_02481_),
    .S(net211),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(_02809_),
    .A1(_02810_),
    .S(net214),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(_02482_),
    .A1(_02484_),
    .S(net211),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(_02485_),
    .A1(_02495_),
    .S(net211),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(_02812_),
    .A1(_02813_),
    .S(net214),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(_02811_),
    .A1(_02814_),
    .S(net217),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(_02490_),
    .A1(_02492_),
    .S(net212),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(_02344_),
    .A1(_02816_),
    .S(_06330_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(_02496_),
    .A1(_02498_),
    .S(net211),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(_02489_),
    .A1(_02499_),
    .S(_06336_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _09726_ (.A0(_02818_),
    .A1(_02819_),
    .S(net214),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(_02817_),
    .A1(_02820_),
    .S(net219),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_2 _09728_ (.A0(_02815_),
    .A1(_02821_),
    .S(net220),
    .X(_02822_));
 sky130_fd_sc_hd__o21a_1 _09729_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_02672_),
    .X(_02823_));
 sky130_fd_sc_hd__nor2_1 _09730_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02824_));
 sky130_fd_sc_hd__or2_1 _09731_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02826_));
 sky130_fd_sc_hd__a21oi_1 _09733_ (.A1(_02825_),
    .A2(_02826_),
    .B1(_02823_),
    .Y(_02827_));
 sky130_fd_sc_hd__a31o_1 _09734_ (.A1(_02823_),
    .A2(_02825_),
    .A3(_02826_),
    .B1(net223),
    .X(_02828_));
 sky130_fd_sc_hd__o221a_1 _09735_ (.A1(net250),
    .A2(_02822_),
    .B1(_02827_),
    .B2(_02828_),
    .C1(net197),
    .X(_02829_));
 sky130_fd_sc_hd__o21a_1 _09736_ (.A1(net215),
    .A2(_02295_),
    .B1(_02345_),
    .X(_02830_));
 sky130_fd_sc_hd__o21a_1 _09737_ (.A1(net217),
    .A2(_02830_),
    .B1(_02347_),
    .X(_02831_));
 sky130_fd_sc_hd__o21a_1 _09738_ (.A1(net221),
    .A2(_02831_),
    .B1(_02342_),
    .X(_02832_));
 sky130_fd_sc_hd__and2_1 _09739_ (.A(net294),
    .B(_06347_),
    .X(_02833_));
 sky130_fd_sc_hd__a21bo_1 _09740_ (.A1(_06338_),
    .A2(_02680_),
    .B1_N(_06332_),
    .X(_02834_));
 sky130_fd_sc_hd__a31o_1 _09741_ (.A1(net285),
    .A2(_06333_),
    .A3(_02834_),
    .B1(_02833_),
    .X(_02835_));
 sky130_fd_sc_hd__or2_1 _09742_ (.A(_06328_),
    .B(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(_06328_),
    .B(_02835_),
    .Y(_02837_));
 sky130_fd_sc_hd__o31a_1 _09744_ (.A1(\div_res[2] ),
    .A2(\div_res[1] ),
    .A3(\div_res[0] ),
    .B1(net160),
    .X(_02838_));
 sky130_fd_sc_hd__xor2_1 _09745_ (.A(\div_res[3] ),
    .B(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__o31a_1 _09746_ (.A1(\div_shifter[34] ),
    .A2(\div_shifter[33] ),
    .A3(\div_shifter[32] ),
    .B1(net230),
    .X(_02840_));
 sky130_fd_sc_hd__xor2_1 _09747_ (.A(\div_shifter[35] ),
    .B(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__a22o_1 _09748_ (.A1(_06324_),
    .A2(net242),
    .B1(_02336_),
    .B2(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__a221o_1 _09749_ (.A1(_06326_),
    .A2(_02321_),
    .B1(_02331_),
    .B2(_06327_),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a221o_1 _09750_ (.A1(_06328_),
    .A2(_02325_),
    .B1(_02334_),
    .B2(_02839_),
    .C1(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__a311o_1 _09751_ (.A1(_02323_),
    .A2(_02836_),
    .A3(_02837_),
    .B1(_02844_),
    .C1(_02829_),
    .X(_02845_));
 sky130_fd_sc_hd__a221o_1 _09752_ (.A1(_02319_),
    .A2(_02822_),
    .B1(_02832_),
    .B2(net170),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__a311o_2 _09753_ (.A1(_02329_),
    .A2(_02807_),
    .A3(_02808_),
    .B1(_02846_),
    .C1(_02806_),
    .X(_02847_));
 sky130_fd_sc_hd__a31o_1 _09754_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .A3(curr_PC[2]),
    .B1(curr_PC[3]),
    .X(_02848_));
 sky130_fd_sc_hd__and4_1 _09755_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .D(curr_PC[3]),
    .X(_02849_));
 sky130_fd_sc_hd__nor2_1 _09756_ (.A(net243),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__a22o_4 _09757_ (.A1(net243),
    .A2(_02847_),
    .B1(_02848_),
    .B2(_02850_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__nor3b_1 _09758_ (.A(_02535_),
    .B(_02644_),
    .C_N(_02804_),
    .Y(_02851_));
 sky130_fd_sc_hd__or2_1 _09759_ (.A(net156),
    .B(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a21oi_4 _09760_ (.A1(_02699_),
    .A2(_02795_),
    .B1(_02794_),
    .Y(_02853_));
 sky130_fd_sc_hd__o21ai_4 _09761_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02792_),
    .Y(_02854_));
 sky130_fd_sc_hd__a21o_2 _09762_ (.A1(_02750_),
    .A2(_02767_),
    .B1(_02766_),
    .X(_02855_));
 sky130_fd_sc_hd__a32o_1 _09763_ (.A1(_00299_),
    .A2(_00676_),
    .A3(_00677_),
    .B1(_00442_),
    .B2(_00293_),
    .X(_02856_));
 sky130_fd_sc_hd__xnor2_1 _09764_ (.A(_00668_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__a22o_1 _09765_ (.A1(net39),
    .A2(net118),
    .B1(net115),
    .B2(net37),
    .X(_02858_));
 sky130_fd_sc_hd__xor2_1 _09766_ (.A(net91),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__and2b_1 _09767_ (.A_N(_02857_),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__and2b_1 _09768_ (.A_N(_02859_),
    .B(_02857_),
    .X(_02861_));
 sky130_fd_sc_hd__or2_1 _09769_ (.A(_02860_),
    .B(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__inv_2 _09770_ (.A(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__a22o_1 _09771_ (.A1(net43),
    .A2(_00309_),
    .B1(_00315_),
    .B2(net41),
    .X(_02864_));
 sky130_fd_sc_hd__xor2_1 _09772_ (.A(net93),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__xor2_1 _09773_ (.A(_02862_),
    .B(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__a21oi_1 _09774_ (.A1(_02735_),
    .A2(_02737_),
    .B1(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__and3_1 _09775_ (.A(_02735_),
    .B(_02737_),
    .C(_02866_),
    .X(_02868_));
 sky130_fd_sc_hd__nor2_2 _09776_ (.A(_02867_),
    .B(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__xor2_4 _09777_ (.A(_02855_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__o21a_1 _09778_ (.A1(_02757_),
    .A2(_02759_),
    .B1(_02755_),
    .X(_02871_));
 sky130_fd_sc_hd__a21oi_1 _09779_ (.A1(_02722_),
    .A2(_02724_),
    .B1(_02721_),
    .Y(_02872_));
 sky130_fd_sc_hd__o21ba_1 _09780_ (.A1(_02746_),
    .A2(_02749_),
    .B1_N(_02745_),
    .X(_02873_));
 sky130_fd_sc_hd__xor2_1 _09781_ (.A(_02872_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__and2b_1 _09782_ (.A_N(_02871_),
    .B(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__xnor2_1 _09783_ (.A(_02871_),
    .B(_02874_),
    .Y(_02876_));
 sky130_fd_sc_hd__o22a_1 _09784_ (.A1(net66),
    .A2(net105),
    .B1(net103),
    .B2(net64),
    .X(_02877_));
 sky130_fd_sc_hd__xnor2_1 _09785_ (.A(net135),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__o22a_1 _09786_ (.A1(net58),
    .A2(net85),
    .B1(net81),
    .B2(net57),
    .X(_02879_));
 sky130_fd_sc_hd__xnor2_1 _09787_ (.A(net137),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__o32a_1 _09788_ (.A1(net134),
    .A2(_00395_),
    .A3(_00397_),
    .B1(net132),
    .B2(net55),
    .X(_02881_));
 sky130_fd_sc_hd__xnor2_1 _09789_ (.A(net172),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__or2_1 _09790_ (.A(_02880_),
    .B(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_02880_),
    .B(_02882_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _09792_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__xor2_1 _09793_ (.A(_02878_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__o22a_1 _09794_ (.A1(net101),
    .A2(net27),
    .B1(net25),
    .B2(net98),
    .X(_02887_));
 sky130_fd_sc_hd__xnor2_2 _09795_ (.A(net87),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__inv_2 _09796_ (.A(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__o22a_1 _09797_ (.A1(net63),
    .A2(net77),
    .B1(net73),
    .B2(net61),
    .X(_02890_));
 sky130_fd_sc_hd__xnor2_1 _09798_ (.A(net122),
    .B(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__nor2_1 _09799_ (.A(_02889_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__xnor2_1 _09800_ (.A(_02888_),
    .B(_02891_),
    .Y(_02893_));
 sky130_fd_sc_hd__o22a_1 _09801_ (.A1(net52),
    .A2(net34),
    .B1(net32),
    .B2(net50),
    .X(_02894_));
 sky130_fd_sc_hd__xnor2_1 _09802_ (.A(net125),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__and2_1 _09803_ (.A(_02893_),
    .B(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__xor2_1 _09804_ (.A(_02893_),
    .B(_02895_),
    .X(_02897_));
 sky130_fd_sc_hd__o22a_1 _09805_ (.A1(net145),
    .A2(net13),
    .B1(net11),
    .B2(net147),
    .X(_02898_));
 sky130_fd_sc_hd__xnor2_1 _09806_ (.A(net190),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__o21ai_1 _09807_ (.A1(_06512_),
    .A2(net7),
    .B1(_06507_),
    .Y(_02900_));
 sky130_fd_sc_hd__o31ai_2 _09808_ (.A1(_06507_),
    .A2(_06511_),
    .A3(net7),
    .B1(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__and2b_1 _09809_ (.A_N(_02901_),
    .B(_02899_),
    .X(_02902_));
 sky130_fd_sc_hd__xor2_1 _09810_ (.A(_02899_),
    .B(_02901_),
    .X(_02903_));
 sky130_fd_sc_hd__and2_1 _09811_ (.A(_02897_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__nor2_1 _09812_ (.A(_02897_),
    .B(_02903_),
    .Y(_02905_));
 sky130_fd_sc_hd__nor2_1 _09813_ (.A(_02904_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__xnor2_1 _09814_ (.A(_02886_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__nor2_1 _09815_ (.A(net128),
    .B(net20),
    .Y(_02908_));
 sky130_fd_sc_hd__a21oi_2 _09816_ (.A1(net193),
    .A2(_02764_),
    .B1(_02763_),
    .Y(_02909_));
 sky130_fd_sc_hd__o22a_1 _09817_ (.A1(_00361_),
    .A2(net10),
    .B1(net5),
    .B2(net130),
    .X(_02910_));
 sky130_fd_sc_hd__xnor2_2 _09818_ (.A(net20),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__nor2_1 _09819_ (.A(_02909_),
    .B(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__xor2_2 _09820_ (.A(_02909_),
    .B(_02911_),
    .X(_02913_));
 sky130_fd_sc_hd__xnor2_2 _09821_ (.A(_02908_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_02907_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__xor2_1 _09823_ (.A(_02907_),
    .B(_02914_),
    .X(_02916_));
 sky130_fd_sc_hd__xnor2_1 _09824_ (.A(_02876_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21o_1 _09825_ (.A1(_02703_),
    .A2(_02705_),
    .B1(_02709_),
    .X(_02918_));
 sky130_fd_sc_hd__o22a_1 _09826_ (.A1(net47),
    .A2(net76),
    .B1(net72),
    .B2(net45),
    .X(_02919_));
 sky130_fd_sc_hd__xnor2_2 _09827_ (.A(net97),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__a22o_1 _09828_ (.A1(net31),
    .A2(_00334_),
    .B1(_00340_),
    .B2(net28),
    .X(_02921_));
 sky130_fd_sc_hd__xnor2_2 _09829_ (.A(net49),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_2 _09830_ (.A(_02920_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__or2_1 _09831_ (.A(_02920_),
    .B(_02922_),
    .X(_02924_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(_02923_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__a21bo_1 _09833_ (.A1(_02769_),
    .A2(_02774_),
    .B1_N(_02773_),
    .X(_02926_));
 sky130_fd_sc_hd__and3_1 _09834_ (.A(_02923_),
    .B(_02924_),
    .C(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__xnor2_1 _09835_ (.A(_02925_),
    .B(_02926_),
    .Y(_02928_));
 sky130_fd_sc_hd__xnor2_1 _09836_ (.A(_02918_),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__nor2_1 _09837_ (.A(_02917_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand2_1 _09838_ (.A(_02917_),
    .B(_02929_),
    .Y(_02931_));
 sky130_fd_sc_hd__and2b_1 _09839_ (.A_N(_02930_),
    .B(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__xor2_4 _09840_ (.A(_02870_),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a21o_1 _09841_ (.A1(_02715_),
    .A2(_02780_),
    .B1(_02779_),
    .X(_02934_));
 sky130_fd_sc_hd__a21o_2 _09842_ (.A1(_02700_),
    .A2(_02714_),
    .B1(_02712_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_2 _09843_ (.A(_02727_),
    .B(_02729_),
    .Y(_02936_));
 sky130_fd_sc_hd__a21oi_4 _09844_ (.A1(_02738_),
    .A2(_02777_),
    .B1(_02776_),
    .Y(_02937_));
 sky130_fd_sc_hd__a21oi_1 _09845_ (.A1(_02727_),
    .A2(_02729_),
    .B1(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__xnor2_4 _09846_ (.A(_02936_),
    .B(_02937_),
    .Y(_02939_));
 sky130_fd_sc_hd__xnor2_4 _09847_ (.A(_02935_),
    .B(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__a21boi_4 _09848_ (.A1(_02784_),
    .A2(_02788_),
    .B1_N(_02787_),
    .Y(_02941_));
 sky130_fd_sc_hd__xnor2_2 _09849_ (.A(_02940_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2b_1 _09850_ (.A_N(_02942_),
    .B(_02934_),
    .Y(_02943_));
 sky130_fd_sc_hd__xnor2_2 _09851_ (.A(_02934_),
    .B(_02942_),
    .Y(_02944_));
 sky130_fd_sc_hd__and2_1 _09852_ (.A(_02933_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__xor2_4 _09853_ (.A(_02933_),
    .B(_02944_),
    .X(_02946_));
 sky130_fd_sc_hd__xnor2_4 _09854_ (.A(_02854_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__or2_1 _09855_ (.A(_02853_),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__and2_1 _09856_ (.A(_02853_),
    .B(_02947_),
    .X(_02949_));
 sky130_fd_sc_hd__xnor2_4 _09857_ (.A(_02853_),
    .B(_02947_),
    .Y(_02950_));
 sky130_fd_sc_hd__or4_1 _09858_ (.A(_02242_),
    .B(_02466_),
    .C(_02638_),
    .D(_02799_),
    .X(_02951_));
 sky130_fd_sc_hd__a21o_1 _09859_ (.A1(_02136_),
    .A2(_02138_),
    .B1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__a21o_1 _09860_ (.A1(_02636_),
    .A2(_02797_),
    .B1(_02798_),
    .X(_02953_));
 sky130_fd_sc_hd__o31a_2 _09861_ (.A1(_02638_),
    .A2(_02641_),
    .A3(_02799_),
    .B1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_1 _09862_ (.A1(_02952_),
    .A2(_02954_),
    .B1(_02950_),
    .Y(_02955_));
 sky130_fd_sc_hd__and3_1 _09863_ (.A(_02950_),
    .B(_02952_),
    .C(_02954_),
    .X(_02956_));
 sky130_fd_sc_hd__or2_2 _09864_ (.A(_02955_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_1 _09865_ (.A1(_02852_),
    .A2(_02957_),
    .B1(_02245_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21oi_1 _09866_ (.A1(_02852_),
    .A2(_02957_),
    .B1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__a21oi_1 _09867_ (.A1(net161),
    .A2(_01808_),
    .B1(_01809_),
    .Y(_02960_));
 sky130_fd_sc_hd__a311oi_1 _09868_ (.A1(net161),
    .A2(_01808_),
    .A3(_01809_),
    .B1(_02330_),
    .C1(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__a31o_1 _09869_ (.A1(_06326_),
    .A2(_06333_),
    .A3(_02834_),
    .B1(_06327_),
    .X(_02962_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(net285),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21a_1 _09871_ (.A1(net285),
    .A2(_06349_),
    .B1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__a21oi_1 _09872_ (.A1(_06321_),
    .A2(_02964_),
    .B1(net236),
    .Y(_02965_));
 sky130_fd_sc_hd__o21a_1 _09873_ (.A1(_06321_),
    .A2(_02964_),
    .B1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__o21ai_2 _09874_ (.A1(net218),
    .A2(_02817_),
    .B1(_02347_),
    .Y(_02967_));
 sky130_fd_sc_hd__a21oi_2 _09875_ (.A1(_06318_),
    .A2(_02967_),
    .B1(_02341_),
    .Y(_02968_));
 sky130_fd_sc_hd__mux2_1 _09876_ (.A0(_02264_),
    .A1(_02272_),
    .S(net214),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(_02279_),
    .A1(_02303_),
    .S(net214),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(_02969_),
    .A1(_02970_),
    .S(net217),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(_02288_),
    .A1(_02310_),
    .S(_06330_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(_02830_),
    .A1(_02972_),
    .S(net219),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(_02971_),
    .A1(_02973_),
    .S(net220),
    .X(_02974_));
 sky130_fd_sc_hd__a21o_1 _09882_ (.A1(net224),
    .A2(_06448_),
    .B1(_02319_),
    .X(_02975_));
 sky130_fd_sc_hd__or4_2 _09883_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_02976_));
 sky130_fd_sc_hd__a21oi_1 _09884_ (.A1(net160),
    .A2(_02976_),
    .B1(\div_res[4] ),
    .Y(_02977_));
 sky130_fd_sc_hd__a311o_1 _09885_ (.A1(\div_res[4] ),
    .A2(net160),
    .A3(_02976_),
    .B1(_02977_),
    .C1(net183),
    .X(_02978_));
 sky130_fd_sc_hd__nor2_1 _09886_ (.A(_06321_),
    .B(net234),
    .Y(_02979_));
 sky130_fd_sc_hd__or4_2 _09887_ (.A(\div_shifter[35] ),
    .B(\div_shifter[34] ),
    .C(\div_shifter[33] ),
    .D(\div_shifter[32] ),
    .X(_02980_));
 sky130_fd_sc_hd__a21oi_1 _09888_ (.A1(net230),
    .A2(_02980_),
    .B1(\div_shifter[36] ),
    .Y(_02981_));
 sky130_fd_sc_hd__a31o_1 _09889_ (.A1(\div_shifter[36] ),
    .A2(net230),
    .A3(_02980_),
    .B1(_02337_),
    .X(_02982_));
 sky130_fd_sc_hd__a2bb2o_1 _09890_ (.A1_N(_02981_),
    .A2_N(_02982_),
    .B1(net222),
    .B2(net242),
    .X(_02983_));
 sky130_fd_sc_hd__o21a_1 _09891_ (.A1(_02823_),
    .A2(_02824_),
    .B1(_02826_),
    .X(_02984_));
 sky130_fd_sc_hd__nor2_1 _09892_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _09893_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02986_));
 sky130_fd_sc_hd__nand2b_1 _09894_ (.A_N(_02985_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__xor2_1 _09895_ (.A(_02984_),
    .B(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__a32o_1 _09896_ (.A1(net250),
    .A2(_06448_),
    .A3(_02988_),
    .B1(_02321_),
    .B2(_06319_),
    .X(_02989_));
 sky130_fd_sc_hd__a311o_1 _09897_ (.A1(reg1_val[4]),
    .A2(net222),
    .A3(_02331_),
    .B1(_02983_),
    .C1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__or3b_1 _09898_ (.A(_02990_),
    .B(_02979_),
    .C_N(_02978_),
    .X(_02991_));
 sky130_fd_sc_hd__a221o_1 _09899_ (.A1(net170),
    .A2(_02968_),
    .B1(_02974_),
    .B2(_02975_),
    .C1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o41a_2 _09900_ (.A1(_02959_),
    .A2(_02961_),
    .A3(_02966_),
    .A4(_02992_),
    .B1(net245),
    .X(_02993_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(curr_PC[4]),
    .B(_02849_),
    .Y(_02994_));
 sky130_fd_sc_hd__or2_1 _09902_ (.A(curr_PC[4]),
    .B(_02849_),
    .X(_02995_));
 sky130_fd_sc_hd__a31o_4 _09903_ (.A1(net248),
    .A2(_02994_),
    .A3(_02995_),
    .B1(_02993_),
    .X(dest_val[4]));
 sky130_fd_sc_hd__nand2_1 _09904_ (.A(_02851_),
    .B(_02957_),
    .Y(_02996_));
 sky130_fd_sc_hd__a21oi_4 _09905_ (.A1(_02854_),
    .A2(_02946_),
    .B1(_02945_),
    .Y(_02997_));
 sky130_fd_sc_hd__o21ai_4 _09906_ (.A1(_02940_),
    .A2(_02941_),
    .B1(_02943_),
    .Y(_02998_));
 sky130_fd_sc_hd__a21o_1 _09907_ (.A1(_02886_),
    .A2(_02906_),
    .B1(_02904_),
    .X(_02999_));
 sky130_fd_sc_hd__a22o_1 _09908_ (.A1(net42),
    .A2(net115),
    .B1(_00309_),
    .B2(net40),
    .X(_03000_));
 sky130_fd_sc_hd__xor2_1 _09909_ (.A(net93),
    .B(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__o22a_1 _09910_ (.A1(net46),
    .A2(net80),
    .B1(net76),
    .B2(net44),
    .X(_03002_));
 sky130_fd_sc_hd__xnor2_1 _09911_ (.A(net96),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__and2_1 _09912_ (.A(_03001_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nor2_1 _09913_ (.A(_03001_),
    .B(_03003_),
    .Y(_03005_));
 sky130_fd_sc_hd__nor2_1 _09914_ (.A(_03004_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__a22o_1 _09915_ (.A1(net36),
    .A2(net118),
    .B1(_00352_),
    .B2(net38),
    .X(_03007_));
 sky130_fd_sc_hd__xor2_1 _09916_ (.A(net90),
    .B(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__xor2_1 _09917_ (.A(_03006_),
    .B(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__o21bai_2 _09918_ (.A1(_02872_),
    .A2(_02873_),
    .B1_N(_02875_),
    .Y(_03010_));
 sky130_fd_sc_hd__xnor2_1 _09919_ (.A(_03009_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__and2b_1 _09920_ (.A_N(_03011_),
    .B(_02999_),
    .X(_03012_));
 sky130_fd_sc_hd__and2b_1 _09921_ (.A_N(_02999_),
    .B(_03011_),
    .X(_03013_));
 sky130_fd_sc_hd__nor2_2 _09922_ (.A(_03012_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__o21ai_1 _09923_ (.A1(_02878_),
    .A2(_02885_),
    .B1(_02883_),
    .Y(_03015_));
 sky130_fd_sc_hd__o21ba_1 _09924_ (.A1(_02892_),
    .A2(_02896_),
    .B1_N(_02902_),
    .X(_03016_));
 sky130_fd_sc_hd__or3b_1 _09925_ (.A(_02892_),
    .B(_02896_),
    .C_N(_02902_),
    .X(_03017_));
 sky130_fd_sc_hd__nand2b_1 _09926_ (.A_N(_03016_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__xor2_1 _09927_ (.A(_03015_),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(net130),
    .B(net20),
    .Y(_03020_));
 sky130_fd_sc_hd__a32o_1 _09929_ (.A1(_00293_),
    .A2(_00676_),
    .A3(_00677_),
    .B1(_00315_),
    .B2(_00442_),
    .X(_03021_));
 sky130_fd_sc_hd__xnor2_1 _09930_ (.A(net70),
    .B(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2_1 _09931_ (.A(_03020_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__or2_1 _09932_ (.A(_03020_),
    .B(_03022_),
    .X(_03024_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__o22a_1 _09934_ (.A1(_00298_),
    .A2(net10),
    .B1(net5),
    .B2(_00361_),
    .X(_03026_));
 sky130_fd_sc_hd__xnor2_2 _09935_ (.A(net20),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__xor2_2 _09936_ (.A(_03025_),
    .B(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__o22a_2 _09937_ (.A1(net145),
    .A2(net11),
    .B1(net7),
    .B2(net147),
    .X(_03029_));
 sky130_fd_sc_hd__xnor2_4 _09938_ (.A(net190),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__o22a_2 _09939_ (.A1(net132),
    .A2(net16),
    .B1(net13),
    .B2(_00169_),
    .X(_03031_));
 sky130_fd_sc_hd__xnor2_4 _09940_ (.A(net172),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__xnor2_4 _09941_ (.A(net195),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2b_1 _09942_ (.A_N(_03030_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__xnor2_4 _09943_ (.A(_03030_),
    .B(_03033_),
    .Y(_03035_));
 sky130_fd_sc_hd__o22a_2 _09944_ (.A1(net65),
    .A2(net85),
    .B1(net81),
    .B2(net58),
    .X(_03036_));
 sky130_fd_sc_hd__xnor2_4 _09945_ (.A(_00323_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__o22a_2 _09946_ (.A1(net55),
    .A2(net105),
    .B1(net103),
    .B2(net66),
    .X(_03038_));
 sky130_fd_sc_hd__xnor2_4 _09947_ (.A(_00327_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__o22a_2 _09948_ (.A1(net57),
    .A2(net77),
    .B1(net73),
    .B2(net63),
    .X(_03040_));
 sky130_fd_sc_hd__xnor2_4 _09949_ (.A(net122),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nor2_1 _09950_ (.A(_03039_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__xnor2_4 _09951_ (.A(_03039_),
    .B(_03041_),
    .Y(_03043_));
 sky130_fd_sc_hd__nor2_1 _09952_ (.A(_03037_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__xor2_4 _09953_ (.A(_03037_),
    .B(_03043_),
    .X(_03045_));
 sky130_fd_sc_hd__xnor2_2 _09954_ (.A(_02923_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__xor2_1 _09955_ (.A(_03035_),
    .B(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__and2_1 _09956_ (.A(_03028_),
    .B(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__xnor2_1 _09957_ (.A(_03028_),
    .B(_03047_),
    .Y(_03049_));
 sky130_fd_sc_hd__nor2_1 _09958_ (.A(_03019_),
    .B(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__and2_1 _09959_ (.A(_03019_),
    .B(_03049_),
    .X(_03051_));
 sky130_fd_sc_hd__or2_1 _09960_ (.A(_03050_),
    .B(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__a21o_1 _09961_ (.A1(_02863_),
    .A2(_02865_),
    .B1(_02860_),
    .X(_03053_));
 sky130_fd_sc_hd__o22a_1 _09962_ (.A1(net60),
    .A2(net34),
    .B1(net32),
    .B2(net52),
    .X(_03054_));
 sky130_fd_sc_hd__xnor2_2 _09963_ (.A(net125),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__a22o_1 _09964_ (.A1(_00174_),
    .A2(net31),
    .B1(net29),
    .B2(_00334_),
    .X(_03056_));
 sky130_fd_sc_hd__xnor2_2 _09965_ (.A(net49),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__and2_1 _09966_ (.A(_03055_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__xor2_2 _09967_ (.A(_03055_),
    .B(_03057_),
    .X(_03059_));
 sky130_fd_sc_hd__o22a_1 _09968_ (.A1(net51),
    .A2(net27),
    .B1(net25),
    .B2(net101),
    .X(_03060_));
 sky130_fd_sc_hd__xnor2_2 _09969_ (.A(net88),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__xnor2_2 _09970_ (.A(_03059_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21oi_2 _09971_ (.A1(_02908_),
    .A2(_02913_),
    .B1(_02912_),
    .Y(_03063_));
 sky130_fd_sc_hd__nor2_1 _09972_ (.A(_03062_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__xor2_2 _09973_ (.A(_03062_),
    .B(_03063_),
    .X(_03065_));
 sky130_fd_sc_hd__xnor2_1 _09974_ (.A(_03053_),
    .B(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__nor2_1 _09975_ (.A(_03052_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _09976_ (.A(_03052_),
    .B(_03066_),
    .Y(_03068_));
 sky130_fd_sc_hd__and2b_1 _09977_ (.A_N(_03067_),
    .B(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__xor2_4 _09978_ (.A(_03014_),
    .B(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__a21o_1 _09979_ (.A1(_02870_),
    .A2(_02931_),
    .B1(_02930_),
    .X(_03071_));
 sky130_fd_sc_hd__a21o_1 _09980_ (.A1(_02935_),
    .A2(_02939_),
    .B1(_02938_),
    .X(_03072_));
 sky130_fd_sc_hd__a21o_1 _09981_ (.A1(_02855_),
    .A2(_02869_),
    .B1(_02867_),
    .X(_03073_));
 sky130_fd_sc_hd__a21oi_1 _09982_ (.A1(_02876_),
    .A2(_02916_),
    .B1(_02915_),
    .Y(_03074_));
 sky130_fd_sc_hd__a21oi_1 _09983_ (.A1(_02918_),
    .A2(_02928_),
    .B1(_02927_),
    .Y(_03075_));
 sky130_fd_sc_hd__nor2_1 _09984_ (.A(_03074_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__xor2_1 _09985_ (.A(_03074_),
    .B(_03075_),
    .X(_03077_));
 sky130_fd_sc_hd__xor2_1 _09986_ (.A(_03073_),
    .B(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__xnor2_1 _09987_ (.A(_03072_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2b_1 _09988_ (.A_N(_03079_),
    .B(_03071_),
    .Y(_03080_));
 sky130_fd_sc_hd__xnor2_2 _09989_ (.A(_03071_),
    .B(_03079_),
    .Y(_03081_));
 sky130_fd_sc_hd__and2_1 _09990_ (.A(_03070_),
    .B(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__xor2_4 _09991_ (.A(_03070_),
    .B(_03081_),
    .X(_03083_));
 sky130_fd_sc_hd__xnor2_4 _09992_ (.A(_02998_),
    .B(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__or2_1 _09993_ (.A(_02997_),
    .B(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__and2_1 _09994_ (.A(_02997_),
    .B(_03084_),
    .X(_03086_));
 sky130_fd_sc_hd__xnor2_4 _09995_ (.A(_02997_),
    .B(_03084_),
    .Y(_03087_));
 sky130_fd_sc_hd__nor4_1 _09996_ (.A(_02466_),
    .B(_02638_),
    .C(_02799_),
    .D(_02950_),
    .Y(_03088_));
 sky130_fd_sc_hd__a21o_1 _09997_ (.A1(_02797_),
    .A2(_02948_),
    .B1(_02949_),
    .X(_03089_));
 sky130_fd_sc_hd__o31a_1 _09998_ (.A1(_02799_),
    .A2(_02801_),
    .A3(_02950_),
    .B1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__a21boi_2 _09999_ (.A1(_02470_),
    .A2(_03088_),
    .B1_N(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__xor2_2 _10000_ (.A(_03087_),
    .B(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__a21o_1 _10001_ (.A1(net161),
    .A2(_02996_),
    .B1(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__a31oi_1 _10002_ (.A1(net162),
    .A2(_02996_),
    .A3(_03092_),
    .B1(net187),
    .Y(_03094_));
 sky130_fd_sc_hd__o21ai_1 _10003_ (.A1(net156),
    .A2(_01810_),
    .B1(_01811_),
    .Y(_03095_));
 sky130_fd_sc_hd__o31a_1 _10004_ (.A1(net156),
    .A2(_01810_),
    .A3(_01811_),
    .B1(net233),
    .X(_03096_));
 sky130_fd_sc_hd__a21boi_1 _10005_ (.A1(_06319_),
    .A2(_02962_),
    .B1_N(_06320_),
    .Y(_03097_));
 sky130_fd_sc_hd__nor2_1 _10006_ (.A(net294),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__a21oi_1 _10007_ (.A1(net294),
    .A2(_06351_),
    .B1(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__xnor2_1 _10008_ (.A(_06314_),
    .B(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__o21ai_1 _10009_ (.A1(net218),
    .A2(_02664_),
    .B1(_02347_),
    .Y(_03101_));
 sky130_fd_sc_hd__a21oi_2 _10010_ (.A1(_06318_),
    .A2(_03101_),
    .B1(_02341_),
    .Y(_03102_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(_02479_),
    .A1(_02483_),
    .S(net214),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(_02486_),
    .A1(_02497_),
    .S(net214),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(_03103_),
    .A1(_03104_),
    .S(net217),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(_02491_),
    .A1(_02500_),
    .S(_06330_),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_02651_),
    .A1(_03106_),
    .S(net219),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(_03105_),
    .A1(_03107_),
    .S(net221),
    .X(_03108_));
 sky130_fd_sc_hd__o21ai_1 _10017_ (.A1(\div_res[4] ),
    .A2(_02976_),
    .B1(net160),
    .Y(_03109_));
 sky130_fd_sc_hd__xnor2_1 _10018_ (.A(\div_res[5] ),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__o21a_1 _10019_ (.A1(\div_shifter[36] ),
    .A2(_02980_),
    .B1(net230),
    .X(_03111_));
 sky130_fd_sc_hd__and2_1 _10020_ (.A(\div_shifter[37] ),
    .B(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__nor2_1 _10021_ (.A(\div_shifter[37] ),
    .B(_03111_),
    .Y(_03113_));
 sky130_fd_sc_hd__o32a_1 _10022_ (.A1(_02337_),
    .A2(_03112_),
    .A3(_03113_),
    .B1(net241),
    .B2(_06309_),
    .X(_03114_));
 sky130_fd_sc_hd__o221a_1 _10023_ (.A1(_06311_),
    .A2(net186),
    .B1(net185),
    .B2(_06313_),
    .C1(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__o21ai_1 _10024_ (.A1(_06315_),
    .A2(net234),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__o21a_1 _10025_ (.A1(_02984_),
    .A2(_02985_),
    .B1(_02986_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_1 _10026_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03118_));
 sky130_fd_sc_hd__nand2_1 _10027_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03119_));
 sky130_fd_sc_hd__and2b_1 _10028_ (.A_N(_03118_),
    .B(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__xnor2_1 _10029_ (.A(_03117_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__a31o_1 _10030_ (.A1(net250),
    .A2(_06448_),
    .A3(_03121_),
    .B1(_03116_),
    .X(_03122_));
 sky130_fd_sc_hd__a221o_1 _10031_ (.A1(_02975_),
    .A2(_03108_),
    .B1(_03110_),
    .B2(_02334_),
    .C1(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__a221o_1 _10032_ (.A1(_02323_),
    .A2(_03100_),
    .B1(_03102_),
    .B2(net169),
    .C1(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__a221o_2 _10033_ (.A1(_03093_),
    .A2(_03094_),
    .B1(_03095_),
    .B2(_03096_),
    .C1(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__a21o_1 _10034_ (.A1(curr_PC[4]),
    .A2(_02849_),
    .B1(curr_PC[5]),
    .X(_03126_));
 sky130_fd_sc_hd__and3_1 _10035_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02849_),
    .X(_03127_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(net243),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__a22o_4 _10037_ (.A1(net243),
    .A2(_03125_),
    .B1(_03126_),
    .B2(_03128_),
    .X(dest_val[5]));
 sky130_fd_sc_hd__or2_1 _10038_ (.A(_02996_),
    .B(_03092_),
    .X(_03129_));
 sky130_fd_sc_hd__a21oi_4 _10039_ (.A1(_02998_),
    .A2(_03083_),
    .B1(_03082_),
    .Y(_03130_));
 sky130_fd_sc_hd__a21bo_2 _10040_ (.A1(_03072_),
    .A2(_03078_),
    .B1_N(_03080_),
    .X(_03131_));
 sky130_fd_sc_hd__o21ai_2 _10041_ (.A1(_06507_),
    .A2(_03032_),
    .B1(_03034_),
    .Y(_03132_));
 sky130_fd_sc_hd__o211a_1 _10042_ (.A1(_03042_),
    .A2(_03044_),
    .B1(_00360_),
    .C1(net21),
    .X(_03133_));
 sky130_fd_sc_hd__a211o_1 _10043_ (.A1(_00360_),
    .A2(net21),
    .B1(_03042_),
    .C1(_03044_),
    .X(_03134_));
 sky130_fd_sc_hd__and2b_1 _10044_ (.A_N(_03133_),
    .B(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__xnor2_2 _10045_ (.A(_03132_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__o22a_1 _10046_ (.A1(net66),
    .A2(net85),
    .B1(net81),
    .B2(net65),
    .X(_03137_));
 sky130_fd_sc_hd__xnor2_2 _10047_ (.A(_00324_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__o32a_1 _10048_ (.A1(net105),
    .A2(_00395_),
    .A3(_00397_),
    .B1(net103),
    .B2(net54),
    .X(_03139_));
 sky130_fd_sc_hd__xnor2_1 _10049_ (.A(_00327_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__o22a_1 _10050_ (.A1(net59),
    .A2(net77),
    .B1(net73),
    .B2(net57),
    .X(_03141_));
 sky130_fd_sc_hd__xnor2_2 _10051_ (.A(net122),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__nor2_1 _10052_ (.A(_03140_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(_03140_),
    .B(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__xnor2_1 _10054_ (.A(_03140_),
    .B(_03142_),
    .Y(_03145_));
 sky130_fd_sc_hd__xnor2_2 _10055_ (.A(_03138_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__a21o_1 _10056_ (.A1(_03059_),
    .A2(_03061_),
    .B1(_03058_),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_1 _10057_ (.A(_03146_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__xor2_2 _10058_ (.A(_03146_),
    .B(_03147_),
    .X(_03149_));
 sky130_fd_sc_hd__o22a_1 _10059_ (.A1(net132),
    .A2(net13),
    .B1(net11),
    .B2(net134),
    .X(_03150_));
 sky130_fd_sc_hd__xnor2_1 _10060_ (.A(net172),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_00143_),
    .B(net7),
    .Y(_03152_));
 sky130_fd_sc_hd__o22a_1 _10062_ (.A1(_00150_),
    .A2(net7),
    .B1(_03152_),
    .B2(net190),
    .X(_03153_));
 sky130_fd_sc_hd__and2_1 _10063_ (.A(_03151_),
    .B(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__nor2_1 _10064_ (.A(_03151_),
    .B(_03153_),
    .Y(_03155_));
 sky130_fd_sc_hd__or2_1 _10065_ (.A(_03154_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__xor2_2 _10066_ (.A(_03149_),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__o22a_1 _10067_ (.A1(net110),
    .A2(net22),
    .B1(net15),
    .B2(_00314_),
    .X(_03158_));
 sky130_fd_sc_hd__xnor2_2 _10068_ (.A(net69),
    .B(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__a22o_1 _10069_ (.A1(_00293_),
    .A2(_01970_),
    .B1(_02085_),
    .B2(_00299_),
    .X(_03160_));
 sky130_fd_sc_hd__xnor2_2 _10070_ (.A(net19),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__a22o_1 _10071_ (.A1(net43),
    .A2(net118),
    .B1(net115),
    .B2(net40),
    .X(_03162_));
 sky130_fd_sc_hd__xor2_2 _10072_ (.A(net93),
    .B(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__nand2_1 _10073_ (.A(_03161_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__xnor2_2 _10074_ (.A(_03161_),
    .B(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__xor2_2 _10075_ (.A(_03159_),
    .B(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__nand2_1 _10076_ (.A(_03157_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__xnor2_2 _10077_ (.A(_03157_),
    .B(_03166_),
    .Y(_03168_));
 sky130_fd_sc_hd__xor2_1 _10078_ (.A(_03136_),
    .B(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__a21o_1 _10079_ (.A1(_03006_),
    .A2(_03008_),
    .B1(_03004_),
    .X(_03170_));
 sky130_fd_sc_hd__o22a_1 _10080_ (.A1(net63),
    .A2(net35),
    .B1(net32),
    .B2(net60),
    .X(_03171_));
 sky130_fd_sc_hd__xnor2_1 _10081_ (.A(net125),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__o22a_1 _10082_ (.A1(net53),
    .A2(net27),
    .B1(net25),
    .B2(net51),
    .X(_03173_));
 sky130_fd_sc_hd__xnor2_1 _10083_ (.A(net88),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand2_1 _10084_ (.A(_03172_),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__or2_1 _10085_ (.A(_03172_),
    .B(_03174_),
    .X(_03176_));
 sky130_fd_sc_hd__and2_1 _10086_ (.A(_03175_),
    .B(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__o21ai_2 _10087_ (.A1(_03025_),
    .A2(_03027_),
    .B1(_03023_),
    .Y(_03178_));
 sky130_fd_sc_hd__and2_1 _10088_ (.A(_03177_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_1 _10089_ (.A(_03177_),
    .B(_03178_),
    .Y(_03180_));
 sky130_fd_sc_hd__and2b_1 _10090_ (.A_N(_03180_),
    .B(_03170_),
    .X(_03181_));
 sky130_fd_sc_hd__xnor2_1 _10091_ (.A(_03170_),
    .B(_03180_),
    .Y(_03182_));
 sky130_fd_sc_hd__and2_1 _10092_ (.A(_03169_),
    .B(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_1 _10093_ (.A(_03169_),
    .B(_03182_),
    .Y(_03184_));
 sky130_fd_sc_hd__nor2_2 _10094_ (.A(_03183_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__a32oi_4 _10095_ (.A1(_02920_),
    .A2(_02922_),
    .A3(_03045_),
    .B1(_03046_),
    .B2(_03035_),
    .Y(_03186_));
 sky130_fd_sc_hd__a22o_1 _10096_ (.A1(net38),
    .A2(_00347_),
    .B1(_00352_),
    .B2(net36),
    .X(_03187_));
 sky130_fd_sc_hd__xor2_1 _10097_ (.A(net90),
    .B(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__a22o_1 _10098_ (.A1(net102),
    .A2(net31),
    .B1(net29),
    .B2(_00174_),
    .X(_03189_));
 sky130_fd_sc_hd__xnor2_1 _10099_ (.A(net49),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__and2_1 _10100_ (.A(_03188_),
    .B(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__nor2_1 _10101_ (.A(_03188_),
    .B(_03190_),
    .Y(_03192_));
 sky130_fd_sc_hd__nor2_2 _10102_ (.A(_03191_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__o22a_2 _10103_ (.A1(_00208_),
    .A2(net84),
    .B1(net80),
    .B2(net44),
    .X(_03194_));
 sky130_fd_sc_hd__xnor2_4 _10104_ (.A(net96),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__xor2_4 _10105_ (.A(_03193_),
    .B(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__a21o_1 _10106_ (.A1(_03015_),
    .A2(_03017_),
    .B1(_03016_),
    .X(_03197_));
 sky130_fd_sc_hd__xor2_4 _10107_ (.A(_03196_),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__nand2b_1 _10108_ (.A_N(_03186_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_4 _10109_ (.A(_03186_),
    .B(_03198_),
    .Y(_03200_));
 sky130_fd_sc_hd__xor2_4 _10110_ (.A(_03185_),
    .B(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__a21o_1 _10111_ (.A1(_03014_),
    .A2(_03068_),
    .B1(_03067_),
    .X(_03202_));
 sky130_fd_sc_hd__a21o_2 _10112_ (.A1(_03009_),
    .A2(_03010_),
    .B1(_03012_),
    .X(_03203_));
 sky130_fd_sc_hd__or2_2 _10113_ (.A(_03048_),
    .B(_03050_),
    .X(_03204_));
 sky130_fd_sc_hd__a21oi_4 _10114_ (.A1(_03053_),
    .A2(_03065_),
    .B1(_03064_),
    .Y(_03205_));
 sky130_fd_sc_hd__o21ba_1 _10115_ (.A1(_03048_),
    .A2(_03050_),
    .B1_N(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__xnor2_4 _10116_ (.A(_03204_),
    .B(_03205_),
    .Y(_03207_));
 sky130_fd_sc_hd__xnor2_2 _10117_ (.A(_03203_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__a21oi_2 _10118_ (.A1(_03073_),
    .A2(_03077_),
    .B1(_03076_),
    .Y(_03209_));
 sky130_fd_sc_hd__xnor2_1 _10119_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__and2b_1 _10120_ (.A_N(_03210_),
    .B(_03202_),
    .X(_03211_));
 sky130_fd_sc_hd__xnor2_2 _10121_ (.A(_03202_),
    .B(_03210_),
    .Y(_03212_));
 sky130_fd_sc_hd__and2_1 _10122_ (.A(_03201_),
    .B(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__xor2_4 _10123_ (.A(_03201_),
    .B(_03212_),
    .X(_03214_));
 sky130_fd_sc_hd__xnor2_4 _10124_ (.A(_03131_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__or2_1 _10125_ (.A(_03130_),
    .B(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__and2_1 _10126_ (.A(_03130_),
    .B(_03215_),
    .X(_03217_));
 sky130_fd_sc_hd__xnor2_4 _10127_ (.A(_03130_),
    .B(_03215_),
    .Y(_03218_));
 sky130_fd_sc_hd__or4_2 _10128_ (.A(_02638_),
    .B(_02799_),
    .C(_02950_),
    .D(_03087_),
    .X(_03219_));
 sky130_fd_sc_hd__or3_1 _10129_ (.A(_02017_),
    .B(_02639_),
    .C(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__a21o_1 _10130_ (.A1(_02641_),
    .A2(_02642_),
    .B1(_03219_),
    .X(_03221_));
 sky130_fd_sc_hd__a21oi_2 _10131_ (.A1(_02948_),
    .A2(_03085_),
    .B1(_03086_),
    .Y(_03222_));
 sky130_fd_sc_hd__a2111oi_1 _10132_ (.A1(_02636_),
    .A2(_02797_),
    .B1(_02798_),
    .C1(_02950_),
    .D1(_03087_),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_1 _10133_ (.A(_03222_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a31oi_2 _10134_ (.A1(_03220_),
    .A2(_03221_),
    .A3(_03224_),
    .B1(_03218_),
    .Y(_03225_));
 sky130_fd_sc_hd__o211a_1 _10135_ (.A1(_02643_),
    .A2(_03219_),
    .B1(_03224_),
    .C1(_03218_),
    .X(_03226_));
 sky130_fd_sc_hd__nor2_1 _10136_ (.A(_03225_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand3_1 _10137_ (.A(net161),
    .B(_03129_),
    .C(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__a21o_1 _10138_ (.A1(net161),
    .A2(_03129_),
    .B1(_03227_),
    .X(_03229_));
 sky130_fd_sc_hd__o21ai_1 _10139_ (.A1(net156),
    .A2(_01812_),
    .B1(_01813_),
    .Y(_03230_));
 sky130_fd_sc_hd__or3_1 _10140_ (.A(net156),
    .B(_01812_),
    .C(_01813_),
    .X(_03231_));
 sky130_fd_sc_hd__o21ai_1 _10141_ (.A1(_06311_),
    .A2(_03097_),
    .B1(_06313_),
    .Y(_03232_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_06353_),
    .A1(_03232_),
    .S(net285),
    .X(_03233_));
 sky130_fd_sc_hd__nand2_1 _10143_ (.A(_06306_),
    .B(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__o21a_1 _10144_ (.A1(_06306_),
    .A2(_03233_),
    .B1(_02323_),
    .X(_03235_));
 sky130_fd_sc_hd__o21a_1 _10145_ (.A1(net218),
    .A2(_02494_),
    .B1(_02347_),
    .X(_03236_));
 sky130_fd_sc_hd__o21a_1 _10146_ (.A1(net220),
    .A2(_03236_),
    .B1(_02342_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _10147_ (.A0(_02657_),
    .A1(_02659_),
    .S(net215),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(_02660_),
    .A1(_02665_),
    .S(net215),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(_03238_),
    .A1(_03239_),
    .S(net217),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(_02663_),
    .A1(_02666_),
    .S(_06330_),
    .X(_03241_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(_02528_),
    .A1(_03241_),
    .S(net219),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(_03240_),
    .A1(_03242_),
    .S(net220),
    .X(_03243_));
 sky130_fd_sc_hd__or3_1 _10153_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_02976_),
    .X(_03244_));
 sky130_fd_sc_hd__a21oi_1 _10154_ (.A1(net160),
    .A2(_03244_),
    .B1(\div_res[6] ),
    .Y(_03245_));
 sky130_fd_sc_hd__a311oi_1 _10155_ (.A1(\div_res[6] ),
    .A2(net160),
    .A3(_03244_),
    .B1(_03245_),
    .C1(net183),
    .Y(_03246_));
 sky130_fd_sc_hd__or3_2 _10156_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_02980_),
    .X(_03247_));
 sky130_fd_sc_hd__a21oi_1 _10157_ (.A1(net230),
    .A2(_03247_),
    .B1(\div_shifter[38] ),
    .Y(_03248_));
 sky130_fd_sc_hd__a31o_1 _10158_ (.A1(\div_shifter[38] ),
    .A2(net230),
    .A3(_03247_),
    .B1(_02337_),
    .X(_03249_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_03248_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a221o_1 _10160_ (.A1(_06302_),
    .A2(net242),
    .B1(_02321_),
    .B2(_06303_),
    .C1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__a221o_1 _10161_ (.A1(_06306_),
    .A2(_02325_),
    .B1(_02331_),
    .B2(_06305_),
    .C1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__o21a_1 _10162_ (.A1(_03117_),
    .A2(_03118_),
    .B1(_03119_),
    .X(_03253_));
 sky130_fd_sc_hd__nor2_1 _10163_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _10164_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03255_));
 sky130_fd_sc_hd__and2b_1 _10165_ (.A_N(_03254_),
    .B(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__xnor2_1 _10166_ (.A(_03253_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a311o_1 _10167_ (.A1(net250),
    .A2(net197),
    .A3(_03257_),
    .B1(_03252_),
    .C1(_03246_),
    .X(_03258_));
 sky130_fd_sc_hd__a221o_1 _10168_ (.A1(net170),
    .A2(_03237_),
    .B1(_03243_),
    .B2(_02975_),
    .C1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__a21o_1 _10169_ (.A1(_03234_),
    .A2(_03235_),
    .B1(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__a31o_1 _10170_ (.A1(net233),
    .A2(_03230_),
    .A3(_03231_),
    .B1(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__a31o_1 _10171_ (.A1(_02245_),
    .A2(_03228_),
    .A3(_03229_),
    .B1(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__and2_1 _10172_ (.A(curr_PC[6]),
    .B(_03127_),
    .X(_03263_));
 sky130_fd_sc_hd__o21ai_1 _10173_ (.A1(curr_PC[6]),
    .A2(_03127_),
    .B1(net248),
    .Y(_03264_));
 sky130_fd_sc_hd__a2bb2o_4 _10174_ (.A1_N(_03263_),
    .A2_N(_03264_),
    .B1(net243),
    .B2(_03262_),
    .X(dest_val[6]));
 sky130_fd_sc_hd__o21a_1 _10175_ (.A1(_03129_),
    .A2(_03227_),
    .B1(net161),
    .X(_03265_));
 sky130_fd_sc_hd__a21oi_4 _10176_ (.A1(_03131_),
    .A2(_03214_),
    .B1(_03213_),
    .Y(_03266_));
 sky130_fd_sc_hd__o21bai_4 _10177_ (.A1(_03208_),
    .A2(_03209_),
    .B1_N(_03211_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21bo_2 _10178_ (.A1(_03149_),
    .A2(_03156_),
    .B1_N(_03148_),
    .X(_03268_));
 sky130_fd_sc_hd__a21o_2 _10179_ (.A1(_03132_),
    .A2(_03134_),
    .B1(_03133_),
    .X(_03269_));
 sky130_fd_sc_hd__o22a_1 _10180_ (.A1(net99),
    .A2(net46),
    .B1(net44),
    .B2(net84),
    .X(_03270_));
 sky130_fd_sc_hd__xnor2_1 _10181_ (.A(net96),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__o22a_1 _10182_ (.A1(net61),
    .A2(net27),
    .B1(net25),
    .B2(net53),
    .X(_03272_));
 sky130_fd_sc_hd__xnor2_1 _10183_ (.A(net88),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__and2_1 _10184_ (.A(_03271_),
    .B(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__nor2_1 _10185_ (.A(_03271_),
    .B(_03273_),
    .Y(_03275_));
 sky130_fd_sc_hd__nor2_2 _10186_ (.A(_03274_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_2 _10187_ (.A1(_00157_),
    .A2(net31),
    .B1(net29),
    .B2(net102),
    .X(_03277_));
 sky130_fd_sc_hd__xnor2_4 _10188_ (.A(net49),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__xnor2_4 _10189_ (.A(_03276_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__and2b_1 _10190_ (.A_N(_03279_),
    .B(_03269_),
    .X(_03280_));
 sky130_fd_sc_hd__xnor2_4 _10191_ (.A(_03269_),
    .B(_03279_),
    .Y(_03281_));
 sky130_fd_sc_hd__xnor2_4 _10192_ (.A(_03268_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__a21oi_1 _10193_ (.A1(_03193_),
    .A2(_03195_),
    .B1(_03191_),
    .Y(_03283_));
 sky130_fd_sc_hd__o22a_1 _10194_ (.A1(net54),
    .A2(net86),
    .B1(net82),
    .B2(net66),
    .X(_03284_));
 sky130_fd_sc_hd__xnor2_1 _10195_ (.A(net138),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__o22a_1 _10196_ (.A1(net57),
    .A2(net35),
    .B1(net32),
    .B2(net63),
    .X(_03286_));
 sky130_fd_sc_hd__xnor2_1 _10197_ (.A(net124),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nor2_1 _10198_ (.A(_03285_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__and2_1 _10199_ (.A(_03285_),
    .B(_03287_),
    .X(_03289_));
 sky130_fd_sc_hd__or2_1 _10200_ (.A(_03288_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__o22a_1 _10201_ (.A1(net65),
    .A2(net77),
    .B1(net73),
    .B2(net59),
    .X(_03291_));
 sky130_fd_sc_hd__xnor2_1 _10202_ (.A(net122),
    .B(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_1 _10203_ (.A(_03290_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__o21a_1 _10204_ (.A1(_03159_),
    .A2(_03165_),
    .B1(_03164_),
    .X(_03294_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(_03293_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__xor2_1 _10206_ (.A(_03293_),
    .B(_03294_),
    .X(_03296_));
 sky130_fd_sc_hd__and2b_1 _10207_ (.A_N(_03283_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__xnor2_1 _10208_ (.A(_03283_),
    .B(_03296_),
    .Y(_03298_));
 sky130_fd_sc_hd__a22o_1 _10209_ (.A1(_00315_),
    .A2(_01970_),
    .B1(_02085_),
    .B2(_00293_),
    .X(_03299_));
 sky130_fd_sc_hd__xnor2_1 _10210_ (.A(net21),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__nor2_1 _10211_ (.A(_03154_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__xor2_1 _10212_ (.A(_03154_),
    .B(_03300_),
    .X(_03302_));
 sky130_fd_sc_hd__and3_1 _10213_ (.A(_00299_),
    .B(net21),
    .C(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__a21oi_1 _10214_ (.A1(_00299_),
    .A2(net21),
    .B1(_03302_),
    .Y(_03304_));
 sky130_fd_sc_hd__or2_1 _10215_ (.A(_03303_),
    .B(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__a32o_1 _10216_ (.A1(_00309_),
    .A2(_00676_),
    .A3(_00677_),
    .B1(_00442_),
    .B2(net115),
    .X(_03306_));
 sky130_fd_sc_hd__xnor2_1 _10217_ (.A(_00668_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a22o_1 _10218_ (.A1(_00247_),
    .A2(_00340_),
    .B1(_00347_),
    .B2(net36),
    .X(_03308_));
 sky130_fd_sc_hd__xor2_1 _10219_ (.A(net90),
    .B(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__nand2b_1 _10220_ (.A_N(_03307_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__xor2_1 _10221_ (.A(_03307_),
    .B(_03309_),
    .X(_03311_));
 sky130_fd_sc_hd__a22o_1 _10222_ (.A1(net40),
    .A2(net118),
    .B1(_00352_),
    .B2(_00234_),
    .X(_03312_));
 sky130_fd_sc_hd__xor2_1 _10223_ (.A(net93),
    .B(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__nand2b_1 _10224_ (.A_N(_03311_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__xnor2_1 _10225_ (.A(_03311_),
    .B(_03313_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21o_1 _10226_ (.A1(_03138_),
    .A2(_03144_),
    .B1(_03143_),
    .X(_03316_));
 sky130_fd_sc_hd__a21o_1 _10227_ (.A1(_00687_),
    .A2(_00688_),
    .B1(net106),
    .X(_03317_));
 sky130_fd_sc_hd__or3_1 _10228_ (.A(net103),
    .B(_00395_),
    .C(_00397_),
    .X(_03318_));
 sky130_fd_sc_hd__a21o_1 _10229_ (.A1(_03317_),
    .A2(_03318_),
    .B1(_00327_),
    .X(_03319_));
 sky130_fd_sc_hd__nand3_1 _10230_ (.A(net135),
    .B(_03317_),
    .C(_03318_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand3_1 _10231_ (.A(net189),
    .B(_03319_),
    .C(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__a21o_1 _10232_ (.A1(_03319_),
    .A2(_03320_),
    .B1(net189),
    .X(_03322_));
 sky130_fd_sc_hd__o22a_1 _10233_ (.A1(net132),
    .A2(net11),
    .B1(net7),
    .B2(net134),
    .X(_03323_));
 sky130_fd_sc_hd__xor2_2 _10234_ (.A(net172),
    .B(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__nand3_1 _10235_ (.A(_03321_),
    .B(_03322_),
    .C(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__a21o_1 _10236_ (.A1(_03321_),
    .A2(_03322_),
    .B1(_03324_),
    .X(_03326_));
 sky130_fd_sc_hd__nand3_1 _10237_ (.A(_03316_),
    .B(_03325_),
    .C(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__a21o_1 _10238_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03316_),
    .X(_03328_));
 sky130_fd_sc_hd__nand3b_1 _10239_ (.A_N(_03175_),
    .B(_03327_),
    .C(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__a21bo_1 _10240_ (.A1(_03327_),
    .A2(_03328_),
    .B1_N(_03175_),
    .X(_03330_));
 sky130_fd_sc_hd__and3_1 _10241_ (.A(_03315_),
    .B(_03329_),
    .C(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__a21oi_1 _10242_ (.A1(_03329_),
    .A2(_03330_),
    .B1(_03315_),
    .Y(_03332_));
 sky130_fd_sc_hd__or3_1 _10243_ (.A(_03305_),
    .B(_03331_),
    .C(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__o21ai_1 _10244_ (.A1(_03331_),
    .A2(_03332_),
    .B1(_03305_),
    .Y(_03334_));
 sky130_fd_sc_hd__and3_1 _10245_ (.A(_03298_),
    .B(_03333_),
    .C(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__a21oi_1 _10246_ (.A1(_03333_),
    .A2(_03334_),
    .B1(_03298_),
    .Y(_03336_));
 sky130_fd_sc_hd__nor2_2 _10247_ (.A(_03335_),
    .B(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__xnor2_4 _10248_ (.A(_03282_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__a21o_1 _10249_ (.A1(_03185_),
    .A2(_03200_),
    .B1(_03183_),
    .X(_03339_));
 sky130_fd_sc_hd__a21oi_4 _10250_ (.A1(_03203_),
    .A2(_03207_),
    .B1(_03206_),
    .Y(_03340_));
 sky130_fd_sc_hd__a21bo_2 _10251_ (.A1(_03196_),
    .A2(_03197_),
    .B1_N(_03199_),
    .X(_03341_));
 sky130_fd_sc_hd__o21ai_4 _10252_ (.A1(_03136_),
    .A2(_03168_),
    .B1(_03167_),
    .Y(_03342_));
 sky130_fd_sc_hd__nor2_2 _10253_ (.A(_03179_),
    .B(_03181_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21ai_1 _10254_ (.A1(_03179_),
    .A2(_03181_),
    .B1(_03342_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_4 _10255_ (.A(_03342_),
    .B(_03343_),
    .Y(_03345_));
 sky130_fd_sc_hd__xor2_4 _10256_ (.A(_03341_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__and2b_1 _10257_ (.A_N(_03340_),
    .B(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__xnor2_4 _10258_ (.A(_03340_),
    .B(_03346_),
    .Y(_03348_));
 sky130_fd_sc_hd__xor2_2 _10259_ (.A(_03339_),
    .B(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__and2_1 _10260_ (.A(_03338_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__xor2_4 _10261_ (.A(_03338_),
    .B(_03349_),
    .X(_03351_));
 sky130_fd_sc_hd__xnor2_4 _10262_ (.A(_03267_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__or2_1 _10263_ (.A(_03266_),
    .B(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__and2_1 _10264_ (.A(_03266_),
    .B(_03352_),
    .X(_03354_));
 sky130_fd_sc_hd__xnor2_4 _10265_ (.A(_03266_),
    .B(_03352_),
    .Y(_03355_));
 sky130_fd_sc_hd__nor2_1 _10266_ (.A(_03087_),
    .B(_03218_),
    .Y(_03356_));
 sky130_fd_sc_hd__or4_1 _10267_ (.A(_02799_),
    .B(_02950_),
    .C(_03087_),
    .D(_03218_),
    .X(_03357_));
 sky130_fd_sc_hd__a21oi_2 _10268_ (.A1(_03085_),
    .A2(_03216_),
    .B1(_03217_),
    .Y(_03358_));
 sky130_fd_sc_hd__a2111oi_1 _10269_ (.A1(_02797_),
    .A2(_02948_),
    .B1(_02949_),
    .C1(_03087_),
    .D1(_03218_),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_1 _10270_ (.A(_03358_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__o21a_1 _10271_ (.A1(_02803_),
    .A2(_03357_),
    .B1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__xor2_4 _10272_ (.A(_03355_),
    .B(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__o21ai_1 _10273_ (.A1(_03265_),
    .A2(_03362_),
    .B1(_02245_),
    .Y(_03363_));
 sky130_fd_sc_hd__a21oi_1 _10274_ (.A1(_03265_),
    .A2(_03362_),
    .B1(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__o21ai_1 _10275_ (.A1(net156),
    .A2(_01814_),
    .B1(_01815_),
    .Y(_03365_));
 sky130_fd_sc_hd__or3_1 _10276_ (.A(net156),
    .B(_01814_),
    .C(_01815_),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_1 _10277_ (.A1(_06303_),
    .A2(_03232_),
    .B1(_06305_),
    .Y(_03367_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(_06355_),
    .A1(_03367_),
    .S(net285),
    .X(_03368_));
 sky130_fd_sc_hd__or2_1 _10279_ (.A(_06300_),
    .B(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_1 _10280_ (.A(_06300_),
    .B(_03368_),
    .Y(_03370_));
 sky130_fd_sc_hd__o21a_1 _10281_ (.A1(net218),
    .A2(_02296_),
    .B1(_02347_),
    .X(_03371_));
 sky130_fd_sc_hd__o21a_1 _10282_ (.A1(net221),
    .A2(_03371_),
    .B1(_02342_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(_02810_),
    .A1(_02812_),
    .S(net214),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(_02813_),
    .A1(_02818_),
    .S(net214),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _10285_ (.A0(_03373_),
    .A1(_03374_),
    .S(net217),
    .X(_03375_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(_02816_),
    .A1(_02819_),
    .S(_06330_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _10287_ (.A0(_02346_),
    .A1(_03376_),
    .S(net219),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(_03375_),
    .A1(_03377_),
    .S(net221),
    .X(_03378_));
 sky130_fd_sc_hd__or2_1 _10289_ (.A(\div_res[6] ),
    .B(_03244_),
    .X(_03379_));
 sky130_fd_sc_hd__a21oi_1 _10290_ (.A1(net160),
    .A2(_03379_),
    .B1(\div_res[7] ),
    .Y(_03380_));
 sky130_fd_sc_hd__a31o_1 _10291_ (.A1(\div_res[7] ),
    .A2(net160),
    .A3(_03379_),
    .B1(net183),
    .X(_03381_));
 sky130_fd_sc_hd__or2_1 _10292_ (.A(\div_shifter[38] ),
    .B(_03247_),
    .X(_03382_));
 sky130_fd_sc_hd__a21oi_1 _10293_ (.A1(net229),
    .A2(_03382_),
    .B1(\div_shifter[39] ),
    .Y(_03383_));
 sky130_fd_sc_hd__a31o_1 _10294_ (.A1(\div_shifter[39] ),
    .A2(net229),
    .A3(_03382_),
    .B1(net232),
    .X(_03384_));
 sky130_fd_sc_hd__o2bb2a_1 _10295_ (.A1_N(_06285_),
    .A2_N(net242),
    .B1(_03383_),
    .B2(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__o221a_1 _10296_ (.A1(_06292_),
    .A2(net186),
    .B1(net185),
    .B2(_06299_),
    .C1(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__o221a_1 _10297_ (.A1(_06300_),
    .A2(net234),
    .B1(_03380_),
    .B2(_03381_),
    .C1(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__o21a_1 _10298_ (.A1(_03253_),
    .A2(_03254_),
    .B1(_03255_),
    .X(_03388_));
 sky130_fd_sc_hd__nor2_1 _10299_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _10300_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03390_));
 sky130_fd_sc_hd__nand2b_1 _10301_ (.A_N(_03389_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__xnor2_1 _10302_ (.A(_03388_),
    .B(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__o31ai_1 _10303_ (.A1(net224),
    .A2(net196),
    .A3(_03392_),
    .B1(_03387_),
    .Y(_03393_));
 sky130_fd_sc_hd__a221o_1 _10304_ (.A1(_02249_),
    .A2(_03372_),
    .B1(_03378_),
    .B2(_02975_),
    .C1(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__a31o_1 _10305_ (.A1(_02323_),
    .A2(_03369_),
    .A3(_03370_),
    .B1(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__a311o_1 _10306_ (.A1(net233),
    .A2(_03365_),
    .A3(_03366_),
    .B1(_03395_),
    .C1(_03364_),
    .X(_03396_));
 sky130_fd_sc_hd__or2_1 _10307_ (.A(curr_PC[7]),
    .B(_03263_),
    .X(_03397_));
 sky130_fd_sc_hd__a21oi_1 _10308_ (.A1(curr_PC[7]),
    .A2(_03263_),
    .B1(net243),
    .Y(_03398_));
 sky130_fd_sc_hd__a22o_4 _10309_ (.A1(net243),
    .A2(_03396_),
    .B1(_03397_),
    .B2(_03398_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__or3_1 _10310_ (.A(_02135_),
    .B(_02243_),
    .C(_02644_),
    .X(_03399_));
 sky130_fd_sc_hd__o21bai_1 _10311_ (.A1(_02955_),
    .A2(_02956_),
    .B1_N(_02471_),
    .Y(_03400_));
 sky130_fd_sc_hd__o21ai_1 _10312_ (.A1(_03225_),
    .A2(_03226_),
    .B1(_02804_),
    .Y(_03401_));
 sky130_fd_sc_hd__or4_1 _10313_ (.A(_03092_),
    .B(_03399_),
    .C(_03400_),
    .D(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__nor2_1 _10314_ (.A(_03362_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__or2_1 _10315_ (.A(net156),
    .B(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__a21oi_1 _10316_ (.A1(_03216_),
    .A2(_03353_),
    .B1(_03354_),
    .Y(_03405_));
 sky130_fd_sc_hd__nor2_1 _10317_ (.A(_03218_),
    .B(_03355_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21oi_2 _10318_ (.A1(_03222_),
    .A2(_03406_),
    .B1(_03405_),
    .Y(_03407_));
 sky130_fd_sc_hd__or4_2 _10319_ (.A(_02950_),
    .B(_03087_),
    .C(_03218_),
    .D(_03355_),
    .X(_03408_));
 sky130_fd_sc_hd__a211o_1 _10320_ (.A1(_02136_),
    .A2(_02138_),
    .B1(_02951_),
    .C1(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__o211ai_4 _10321_ (.A1(_02954_),
    .A2(_03408_),
    .B1(_03409_),
    .C1(_03407_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21oi_4 _10322_ (.A1(_03267_),
    .A2(_03351_),
    .B1(_03350_),
    .Y(_03411_));
 sky130_fd_sc_hd__a21oi_4 _10323_ (.A1(_03339_),
    .A2(_03348_),
    .B1(_03347_),
    .Y(_03412_));
 sky130_fd_sc_hd__o22a_1 _10324_ (.A1(net111),
    .A2(net10),
    .B1(net5),
    .B2(_00314_),
    .X(_03413_));
 sky130_fd_sc_hd__xnor2_1 _10325_ (.A(net19),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _10326_ (.A(_00293_),
    .B(net21),
    .Y(_03415_));
 sky130_fd_sc_hd__o22a_1 _10327_ (.A1(net120),
    .A2(net23),
    .B1(net14),
    .B2(net117),
    .X(_03416_));
 sky130_fd_sc_hd__xnor2_1 _10328_ (.A(net69),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__or2_1 _10329_ (.A(_03415_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__xnor2_1 _10330_ (.A(_03415_),
    .B(_03417_),
    .Y(_03419_));
 sky130_fd_sc_hd__or2_1 _10331_ (.A(_03414_),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(_03414_),
    .B(_03419_),
    .Y(_03421_));
 sky130_fd_sc_hd__and2_1 _10333_ (.A(_03420_),
    .B(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__o21bai_1 _10334_ (.A1(_03290_),
    .A2(_03292_),
    .B1_N(_03288_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21bo_1 _10335_ (.A1(_03322_),
    .A2(_03324_),
    .B1_N(_03321_),
    .X(_03424_));
 sky130_fd_sc_hd__o22a_1 _10336_ (.A1(net103),
    .A2(net13),
    .B1(net11),
    .B2(net105),
    .X(_03425_));
 sky130_fd_sc_hd__xnor2_1 _10337_ (.A(_00328_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__o21ba_1 _10338_ (.A1(_00168_),
    .A2(net7),
    .B1_N(net172),
    .X(_03427_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(_00167_),
    .B(net7),
    .Y(_03428_));
 sky130_fd_sc_hd__a21o_1 _10340_ (.A1(net173),
    .A2(_03428_),
    .B1(_03427_),
    .X(_03429_));
 sky130_fd_sc_hd__nor2_2 _10341_ (.A(_03426_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__xor2_1 _10342_ (.A(_03426_),
    .B(_03429_),
    .X(_03431_));
 sky130_fd_sc_hd__a21oi_1 _10343_ (.A1(_03321_),
    .A2(_03325_),
    .B1(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__xnor2_1 _10344_ (.A(_03424_),
    .B(_03431_),
    .Y(_03433_));
 sky130_fd_sc_hd__xor2_1 _10345_ (.A(_03423_),
    .B(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__o22a_1 _10346_ (.A1(net101),
    .A2(net46),
    .B1(net44),
    .B2(net99),
    .X(_03435_));
 sky130_fd_sc_hd__xnor2_1 _10347_ (.A(net95),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a22o_1 _10348_ (.A1(net43),
    .A2(_00347_),
    .B1(_00352_),
    .B2(net40),
    .X(_03437_));
 sky130_fd_sc_hd__xor2_1 _10349_ (.A(net92),
    .B(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__and2_1 _10350_ (.A(_03436_),
    .B(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__nor2_1 _10351_ (.A(_03436_),
    .B(_03438_),
    .Y(_03440_));
 sky130_fd_sc_hd__nor2_1 _10352_ (.A(_03439_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__a22o_1 _10353_ (.A1(net38),
    .A2(_00334_),
    .B1(_00340_),
    .B2(net36),
    .X(_03442_));
 sky130_fd_sc_hd__xor2_1 _10354_ (.A(net90),
    .B(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__xor2_1 _10355_ (.A(_03441_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__xor2_1 _10356_ (.A(_03434_),
    .B(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__xnor2_1 _10357_ (.A(_03422_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__a21o_1 _10358_ (.A1(_03276_),
    .A2(_03278_),
    .B1(_03274_),
    .X(_03447_));
 sky130_fd_sc_hd__o32a_1 _10359_ (.A1(net86),
    .A2(_00395_),
    .A3(_00397_),
    .B1(net82),
    .B2(net54),
    .X(_03448_));
 sky130_fd_sc_hd__xnor2_2 _10360_ (.A(_00324_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__o22a_1 _10361_ (.A1(net66),
    .A2(net78),
    .B1(net74),
    .B2(net65),
    .X(_03450_));
 sky130_fd_sc_hd__xor2_2 _10362_ (.A(net122),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_1 _10363_ (.A(_03449_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21oi_1 _10364_ (.A1(_03310_),
    .A2(_03314_),
    .B1(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__and3_1 _10365_ (.A(_03310_),
    .B(_03314_),
    .C(_03452_),
    .X(_03454_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(_03453_),
    .B(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__and2b_1 _10367_ (.A_N(_03455_),
    .B(_03447_),
    .X(_03456_));
 sky130_fd_sc_hd__xor2_1 _10368_ (.A(_03447_),
    .B(_03455_),
    .X(_03457_));
 sky130_fd_sc_hd__nor2_1 _10369_ (.A(_03446_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_1 _10370_ (.A(_03446_),
    .B(_03457_),
    .Y(_03459_));
 sky130_fd_sc_hd__and2b_1 _10371_ (.A_N(_03458_),
    .B(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__nand2_1 _10372_ (.A(_03327_),
    .B(_03329_),
    .Y(_03461_));
 sky130_fd_sc_hd__o22a_1 _10373_ (.A1(net58),
    .A2(net35),
    .B1(net33),
    .B2(net56),
    .X(_03462_));
 sky130_fd_sc_hd__xnor2_1 _10374_ (.A(net126),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__a22o_1 _10375_ (.A1(_00148_),
    .A2(net31),
    .B1(net29),
    .B2(_00157_),
    .X(_03464_));
 sky130_fd_sc_hd__xnor2_1 _10376_ (.A(net49),
    .B(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__and2_1 _10377_ (.A(_03463_),
    .B(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__nor2_1 _10378_ (.A(_03463_),
    .B(_03465_),
    .Y(_03467_));
 sky130_fd_sc_hd__nor2_1 _10379_ (.A(_03466_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__o22a_1 _10380_ (.A1(net62),
    .A2(net27),
    .B1(net25),
    .B2(net61),
    .X(_03469_));
 sky130_fd_sc_hd__xnor2_2 _10381_ (.A(net88),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__xor2_1 _10382_ (.A(_03468_),
    .B(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__o21a_1 _10383_ (.A1(_03301_),
    .A2(_03303_),
    .B1(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__or3_1 _10384_ (.A(_03301_),
    .B(_03303_),
    .C(_03471_),
    .X(_03473_));
 sky130_fd_sc_hd__and2b_1 _10385_ (.A_N(_03472_),
    .B(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__xor2_1 _10386_ (.A(_03461_),
    .B(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__xnor2_1 _10387_ (.A(_03460_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__o21bai_1 _10388_ (.A1(_03282_),
    .A2(_03336_),
    .B1_N(_03335_),
    .Y(_03477_));
 sky130_fd_sc_hd__a21o_1 _10389_ (.A1(_03268_),
    .A2(_03281_),
    .B1(_03280_),
    .X(_03478_));
 sky130_fd_sc_hd__or2_1 _10390_ (.A(_03295_),
    .B(_03297_),
    .X(_03479_));
 sky130_fd_sc_hd__o21ba_1 _10391_ (.A1(_03305_),
    .A2(_03332_),
    .B1_N(_03331_),
    .X(_03480_));
 sky130_fd_sc_hd__o21ba_1 _10392_ (.A1(_03295_),
    .A2(_03297_),
    .B1_N(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__xnor2_1 _10393_ (.A(_03479_),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor2_1 _10394_ (.A(_03478_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__a21boi_1 _10395_ (.A1(_03341_),
    .A2(_03345_),
    .B1_N(_03344_),
    .Y(_03484_));
 sky130_fd_sc_hd__nor2_1 _10396_ (.A(_03483_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__xor2_1 _10397_ (.A(_03483_),
    .B(_03484_),
    .X(_03486_));
 sky130_fd_sc_hd__xnor2_1 _10398_ (.A(_03477_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__nor2_1 _10399_ (.A(_03476_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__and2_1 _10400_ (.A(_03476_),
    .B(_03487_),
    .X(_03489_));
 sky130_fd_sc_hd__nor2_2 _10401_ (.A(_03488_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__xor2_4 _10402_ (.A(_03412_),
    .B(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__or2_1 _10403_ (.A(_03411_),
    .B(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__and2_1 _10404_ (.A(_03411_),
    .B(_03491_),
    .X(_03493_));
 sky130_fd_sc_hd__xnor2_4 _10405_ (.A(_03411_),
    .B(_03491_),
    .Y(_03494_));
 sky130_fd_sc_hd__xor2_2 _10406_ (.A(_03410_),
    .B(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__o21ai_1 _10407_ (.A1(_03404_),
    .A2(_03495_),
    .B1(_02245_),
    .Y(_03496_));
 sky130_fd_sc_hd__a21o_1 _10408_ (.A1(_03404_),
    .A2(_03495_),
    .B1(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__o21ai_1 _10409_ (.A1(net157),
    .A2(_01816_),
    .B1(_01817_),
    .Y(_03498_));
 sky130_fd_sc_hd__o31a_1 _10410_ (.A1(net157),
    .A2(_01816_),
    .A3(_01817_),
    .B1(net233),
    .X(_03499_));
 sky130_fd_sc_hd__nand2_1 _10411_ (.A(_03498_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__o21a_1 _10412_ (.A1(_06292_),
    .A2(_03367_),
    .B1(_06299_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _10413_ (.A0(_06357_),
    .A1(_03501_),
    .S(net285),
    .X(_03502_));
 sky130_fd_sc_hd__nor2_1 _10414_ (.A(_06267_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__a211o_1 _10415_ (.A1(_06267_),
    .A2(_03502_),
    .B1(_03503_),
    .C1(net236),
    .X(_03504_));
 sky130_fd_sc_hd__o21a_1 _10416_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03390_),
    .X(_03505_));
 sky130_fd_sc_hd__nor2_1 _10417_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2b_1 _10419_ (.A_N(_03506_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__xnor2_1 _10420_ (.A(_03505_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__or2_1 _10421_ (.A(net218),
    .B(_02280_),
    .X(_03510_));
 sky130_fd_sc_hd__o211a_1 _10422_ (.A1(net219),
    .A2(_02311_),
    .B1(_03510_),
    .C1(_06318_),
    .X(_03511_));
 sky130_fd_sc_hd__a21oi_2 _10423_ (.A1(net220),
    .A2(_03371_),
    .B1(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(_03509_),
    .A1(_03512_),
    .S(net223),
    .X(_03513_));
 sky130_fd_sc_hd__or2_1 _10425_ (.A(\div_res[7] ),
    .B(_03379_),
    .X(_03514_));
 sky130_fd_sc_hd__a21oi_1 _10426_ (.A1(net160),
    .A2(_03514_),
    .B1(\div_res[8] ),
    .Y(_03515_));
 sky130_fd_sc_hd__a31o_1 _10427_ (.A1(\div_res[8] ),
    .A2(net160),
    .A3(_03514_),
    .B1(net183),
    .X(_03516_));
 sky130_fd_sc_hd__a21oi_1 _10428_ (.A1(_06258_),
    .A2(_02325_),
    .B1(_02321_),
    .Y(_03517_));
 sky130_fd_sc_hd__or2_1 _10429_ (.A(\div_shifter[39] ),
    .B(_03382_),
    .X(_03518_));
 sky130_fd_sc_hd__a21oi_1 _10430_ (.A1(net229),
    .A2(_03518_),
    .B1(\div_shifter[40] ),
    .Y(_03519_));
 sky130_fd_sc_hd__a31o_1 _10431_ (.A1(\div_shifter[40] ),
    .A2(net229),
    .A3(_03518_),
    .B1(net232),
    .X(_03520_));
 sky130_fd_sc_hd__o2bb2a_1 _10432_ (.A1_N(_06241_),
    .A2_N(net242),
    .B1(_03519_),
    .B2(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__o221a_1 _10433_ (.A1(_06258_),
    .A2(net185),
    .B1(_03517_),
    .B2(_06249_),
    .C1(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__o21ai_2 _10434_ (.A1(net221),
    .A2(_03377_),
    .B1(_02342_),
    .Y(_03523_));
 sky130_fd_sc_hd__o221a_1 _10435_ (.A1(_03515_),
    .A2(_03516_),
    .B1(_03523_),
    .B2(net168),
    .C1(_03522_),
    .X(_03524_));
 sky130_fd_sc_hd__o221a_1 _10436_ (.A1(_02320_),
    .A2(_03512_),
    .B1(_03513_),
    .B2(net196),
    .C1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__a41o_1 _10437_ (.A1(_03497_),
    .A2(_03500_),
    .A3(_03504_),
    .A4(_03525_),
    .B1(net248),
    .X(_03526_));
 sky130_fd_sc_hd__and3_2 _10438_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03263_),
    .X(_03527_));
 sky130_fd_sc_hd__a21oi_1 _10439_ (.A1(curr_PC[7]),
    .A2(_03263_),
    .B1(curr_PC[8]),
    .Y(_03528_));
 sky130_fd_sc_hd__o31ai_4 _10440_ (.A1(net243),
    .A2(_03527_),
    .A3(_03528_),
    .B1(_03526_),
    .Y(dest_val[8]));
 sky130_fd_sc_hd__xor2_1 _10441_ (.A(curr_PC[9]),
    .B(_03527_),
    .X(_03529_));
 sky130_fd_sc_hd__a21o_1 _10442_ (.A1(_03403_),
    .A2(_03495_),
    .B1(net156),
    .X(_03530_));
 sky130_fd_sc_hd__o21ba_2 _10443_ (.A1(_03412_),
    .A2(_03489_),
    .B1_N(_03488_),
    .X(_03531_));
 sky130_fd_sc_hd__a21o_2 _10444_ (.A1(_03477_),
    .A2(_03486_),
    .B1(_03485_),
    .X(_03532_));
 sky130_fd_sc_hd__a21o_1 _10445_ (.A1(_03423_),
    .A2(_03433_),
    .B1(_03432_),
    .X(_03533_));
 sky130_fd_sc_hd__o22a_1 _10446_ (.A1(net54),
    .A2(net78),
    .B1(net74),
    .B2(net66),
    .X(_03534_));
 sky130_fd_sc_hd__xnor2_1 _10447_ (.A(net122),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__o22a_1 _10448_ (.A1(net56),
    .A2(net27),
    .B1(net25),
    .B2(net62),
    .X(_03536_));
 sky130_fd_sc_hd__xnor2_1 _10449_ (.A(net88),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2b_1 _10450_ (.A_N(_03535_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__xor2_1 _10451_ (.A(_03535_),
    .B(_03537_),
    .X(_03539_));
 sky130_fd_sc_hd__o22a_1 _10452_ (.A1(net64),
    .A2(net35),
    .B1(net33),
    .B2(net58),
    .X(_03540_));
 sky130_fd_sc_hd__xnor2_1 _10453_ (.A(net126),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2b_1 _10454_ (.A_N(_03539_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2b_1 _10455_ (.A_N(_03541_),
    .B(_03539_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_03542_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_1 _10457_ (.A1(_03418_),
    .A2(_03420_),
    .B1(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__and3_1 _10458_ (.A(_03418_),
    .B(_03420_),
    .C(_03544_),
    .X(_03546_));
 sky130_fd_sc_hd__or2_1 _10459_ (.A(_03545_),
    .B(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__and2b_1 _10460_ (.A_N(_03547_),
    .B(_03533_),
    .X(_03548_));
 sky130_fd_sc_hd__xnor2_1 _10461_ (.A(_03533_),
    .B(_03547_),
    .Y(_03549_));
 sky130_fd_sc_hd__a21oi_2 _10462_ (.A1(_03468_),
    .A2(_03470_),
    .B1(_03466_),
    .Y(_03550_));
 sky130_fd_sc_hd__o22a_2 _10463_ (.A1(net104),
    .A2(net11),
    .B1(net7),
    .B2(net105),
    .X(_03551_));
 sky130_fd_sc_hd__xnor2_4 _10464_ (.A(_00328_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__a21o_1 _10465_ (.A1(_00687_),
    .A2(_00688_),
    .B1(net85),
    .X(_03553_));
 sky130_fd_sc_hd__or3_1 _10466_ (.A(net81),
    .B(_00395_),
    .C(_00397_),
    .X(_03554_));
 sky130_fd_sc_hd__a21o_1 _10467_ (.A1(_03553_),
    .A2(_03554_),
    .B1(net138),
    .X(_03555_));
 sky130_fd_sc_hd__nand3_1 _10468_ (.A(net138),
    .B(_03553_),
    .C(_03554_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand3_1 _10469_ (.A(net173),
    .B(_03555_),
    .C(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__a21o_1 _10470_ (.A1(_03555_),
    .A2(_03556_),
    .B1(net173),
    .X(_03558_));
 sky130_fd_sc_hd__nand2_2 _10471_ (.A(_03557_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__xnor2_4 _10472_ (.A(_03552_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__a21o_1 _10473_ (.A1(_03441_),
    .A2(_03443_),
    .B1(_03439_),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _10474_ (.A(_03560_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__xnor2_2 _10475_ (.A(_03560_),
    .B(_03561_),
    .Y(_03563_));
 sky130_fd_sc_hd__nor2_1 _10476_ (.A(_03550_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__and2_1 _10477_ (.A(_03550_),
    .B(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__o22a_1 _10478_ (.A1(net72),
    .A2(net22),
    .B1(net14),
    .B2(net120),
    .X(_03566_));
 sky130_fd_sc_hd__xnor2_1 _10479_ (.A(net69),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__o22a_1 _10480_ (.A1(net116),
    .A2(net10),
    .B1(net5),
    .B2(net111),
    .X(_03568_));
 sky130_fd_sc_hd__xnor2_1 _10481_ (.A(net19),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__a22o_1 _10482_ (.A1(net42),
    .A2(_00340_),
    .B1(_00347_),
    .B2(net40),
    .X(_03570_));
 sky130_fd_sc_hd__xor2_1 _10483_ (.A(net92),
    .B(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__nand2b_1 _10484_ (.A_N(_03569_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2b_1 _10485_ (.A_N(_03571_),
    .B(_03569_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _10486_ (.A(_03572_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__or2_1 _10487_ (.A(_03567_),
    .B(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__nand2_1 _10488_ (.A(_03567_),
    .B(_03574_),
    .Y(_03576_));
 sky130_fd_sc_hd__and2_1 _10489_ (.A(_03575_),
    .B(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__nor2_1 _10490_ (.A(_00314_),
    .B(net19),
    .Y(_03578_));
 sky130_fd_sc_hd__and3_1 _10491_ (.A(_03449_),
    .B(_03451_),
    .C(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__a21oi_1 _10492_ (.A1(_03449_),
    .A2(_03451_),
    .B1(_03578_),
    .Y(_03580_));
 sky130_fd_sc_hd__or2_1 _10493_ (.A(_03579_),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__xor2_2 _10494_ (.A(_03430_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__a22o_1 _10495_ (.A1(_00174_),
    .A2(net38),
    .B1(net36),
    .B2(_00334_),
    .X(_03583_));
 sky130_fd_sc_hd__xor2_1 _10496_ (.A(net90),
    .B(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_1 _10497_ (.A1(_06522_),
    .A2(net31),
    .B1(net29),
    .B2(_00148_),
    .X(_03585_));
 sky130_fd_sc_hd__xnor2_1 _10498_ (.A(net49),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(_03584_),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__nor2_1 _10500_ (.A(_03584_),
    .B(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__nor2_1 _10501_ (.A(_03587_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__o22a_1 _10502_ (.A1(net51),
    .A2(net46),
    .B1(net44),
    .B2(net101),
    .X(_03590_));
 sky130_fd_sc_hd__xnor2_2 _10503_ (.A(net95),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__xor2_2 _10504_ (.A(_03589_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__xor2_1 _10505_ (.A(_03582_),
    .B(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__xnor2_1 _10506_ (.A(_03577_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__or3_1 _10507_ (.A(_03564_),
    .B(_03565_),
    .C(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__o21ai_1 _10508_ (.A1(_03564_),
    .A2(_03565_),
    .B1(_03594_),
    .Y(_03596_));
 sky130_fd_sc_hd__and3_1 _10509_ (.A(_03549_),
    .B(_03595_),
    .C(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a21oi_1 _10510_ (.A1(_03595_),
    .A2(_03596_),
    .B1(_03549_),
    .Y(_03598_));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_03597_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__a21o_1 _10512_ (.A1(_03459_),
    .A2(_03475_),
    .B1(_03458_),
    .X(_03600_));
 sky130_fd_sc_hd__a21o_1 _10513_ (.A1(_03461_),
    .A2(_03473_),
    .B1(_03472_),
    .X(_03601_));
 sky130_fd_sc_hd__a32o_1 _10514_ (.A1(_03420_),
    .A2(_03421_),
    .A3(_03445_),
    .B1(_03444_),
    .B2(_03434_),
    .X(_03602_));
 sky130_fd_sc_hd__nor2_1 _10515_ (.A(_03453_),
    .B(_03456_),
    .Y(_03603_));
 sky130_fd_sc_hd__o21a_1 _10516_ (.A1(_03453_),
    .A2(_03456_),
    .B1(_03602_),
    .X(_03604_));
 sky130_fd_sc_hd__xnor2_1 _10517_ (.A(_03602_),
    .B(_03603_),
    .Y(_03605_));
 sky130_fd_sc_hd__xnor2_1 _10518_ (.A(_03601_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__a21oi_2 _10519_ (.A1(_03478_),
    .A2(_03482_),
    .B1(_03481_),
    .Y(_03607_));
 sky130_fd_sc_hd__xnor2_1 _10520_ (.A(_03606_),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__nand2b_1 _10521_ (.A_N(_03608_),
    .B(_03600_),
    .Y(_03609_));
 sky130_fd_sc_hd__xnor2_1 _10522_ (.A(_03600_),
    .B(_03608_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand2_1 _10523_ (.A(_03599_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__or2_1 _10524_ (.A(_03599_),
    .B(_03610_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_2 _10525_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__xor2_4 _10526_ (.A(_03532_),
    .B(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__or2_1 _10527_ (.A(_03531_),
    .B(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__and2_1 _10528_ (.A(_03531_),
    .B(_03614_),
    .X(_03616_));
 sky130_fd_sc_hd__xnor2_4 _10529_ (.A(_03531_),
    .B(_03614_),
    .Y(_03617_));
 sky130_fd_sc_hd__a21oi_2 _10530_ (.A1(_03353_),
    .A2(_03492_),
    .B1(_03493_),
    .Y(_03618_));
 sky130_fd_sc_hd__nor2_2 _10531_ (.A(_03355_),
    .B(_03494_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21oi_1 _10532_ (.A1(_03358_),
    .A2(_03619_),
    .B1(_03618_),
    .Y(_03620_));
 sky130_fd_sc_hd__a21o_1 _10533_ (.A1(_03358_),
    .A2(_03619_),
    .B1(_03618_),
    .X(_03621_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_03356_),
    .B(_03619_),
    .Y(_03622_));
 sky130_fd_sc_hd__o2111ai_1 _10535_ (.A1(_02467_),
    .A2(_02469_),
    .B1(_03088_),
    .C1(_03356_),
    .D1(_03619_),
    .Y(_03623_));
 sky130_fd_sc_hd__o211a_2 _10536_ (.A1(_03090_),
    .A2(_03622_),
    .B1(_03623_),
    .C1(_03620_),
    .X(_03624_));
 sky130_fd_sc_hd__xnor2_2 _10537_ (.A(_03617_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__a21oi_1 _10538_ (.A1(_03530_),
    .A2(_03625_),
    .B1(net187),
    .Y(_03626_));
 sky130_fd_sc_hd__o21a_1 _10539_ (.A1(_03530_),
    .A2(_03625_),
    .B1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__o21ai_1 _10540_ (.A1(net157),
    .A2(_01818_),
    .B1(_01820_),
    .Y(_03628_));
 sky130_fd_sc_hd__or3_1 _10541_ (.A(net157),
    .B(_01818_),
    .C(_01820_),
    .X(_03629_));
 sky130_fd_sc_hd__o21a_1 _10542_ (.A1(_06249_),
    .A2(_03501_),
    .B1(_06258_),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(_06359_),
    .A1(_03630_),
    .S(net285),
    .X(_03631_));
 sky130_fd_sc_hd__a21oi_1 _10544_ (.A1(_06223_),
    .A2(_03631_),
    .B1(net236),
    .Y(_03632_));
 sky130_fd_sc_hd__o21a_1 _10545_ (.A1(_06223_),
    .A2(_03631_),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__o21a_1 _10546_ (.A1(_03505_),
    .A2(_03506_),
    .B1(_03507_),
    .X(_03634_));
 sky130_fd_sc_hd__nor2_1 _10547_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03635_));
 sky130_fd_sc_hd__nand2_1 _10548_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2b_1 _10549_ (.A_N(_03635_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__xor2_1 _10550_ (.A(_03634_),
    .B(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(_02487_),
    .A1(_02501_),
    .S(net217),
    .X(_03639_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(_03236_),
    .A1(_03639_),
    .S(_06318_),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(_03638_),
    .A1(_03640_),
    .S(net223),
    .X(_03641_));
 sky130_fd_sc_hd__or3_1 _10554_ (.A(\div_res[8] ),
    .B(\div_res[7] ),
    .C(_03379_),
    .X(_03642_));
 sky130_fd_sc_hd__a21oi_1 _10555_ (.A1(net159),
    .A2(_03642_),
    .B1(\div_res[9] ),
    .Y(_03643_));
 sky130_fd_sc_hd__a31o_1 _10556_ (.A1(\div_res[9] ),
    .A2(net159),
    .A3(_03642_),
    .B1(net183),
    .X(_03644_));
 sky130_fd_sc_hd__a21oi_1 _10557_ (.A1(_06214_),
    .A2(_02325_),
    .B1(_02321_),
    .Y(_03645_));
 sky130_fd_sc_hd__or3_1 _10558_ (.A(\div_shifter[40] ),
    .B(\div_shifter[39] ),
    .C(_03382_),
    .X(_03646_));
 sky130_fd_sc_hd__a21oi_1 _10559_ (.A1(net229),
    .A2(_03646_),
    .B1(\div_shifter[41] ),
    .Y(_03647_));
 sky130_fd_sc_hd__a31o_1 _10560_ (.A1(\div_shifter[41] ),
    .A2(net229),
    .A3(_03646_),
    .B1(net232),
    .X(_03648_));
 sky130_fd_sc_hd__o221a_1 _10561_ (.A1(_06196_),
    .A2(net241),
    .B1(_02332_),
    .B2(_06214_),
    .C1(net245),
    .X(_03649_));
 sky130_fd_sc_hd__o221a_1 _10562_ (.A1(_06205_),
    .A2(_03645_),
    .B1(_03647_),
    .B2(_03648_),
    .C1(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__o21ai_1 _10563_ (.A1(_03643_),
    .A2(_03644_),
    .B1(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__o21ai_2 _10564_ (.A1(net220),
    .A2(_03242_),
    .B1(_02342_),
    .Y(_03652_));
 sky130_fd_sc_hd__inv_2 _10565_ (.A(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__a221o_1 _10566_ (.A1(_02319_),
    .A2(_03640_),
    .B1(_03653_),
    .B2(net170),
    .C1(_03651_),
    .X(_03654_));
 sky130_fd_sc_hd__a211o_1 _10567_ (.A1(net197),
    .A2(_03641_),
    .B1(_03654_),
    .C1(_03633_),
    .X(_03655_));
 sky130_fd_sc_hd__a31o_1 _10568_ (.A1(net233),
    .A2(_03628_),
    .A3(_03629_),
    .B1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__o22a_4 _10569_ (.A1(net244),
    .A2(_03529_),
    .B1(_03627_),
    .B2(_03656_),
    .X(dest_val[9]));
 sky130_fd_sc_hd__or4bb_4 _10570_ (.A(_03362_),
    .B(_03402_),
    .C_N(_03495_),
    .D_N(_03625_),
    .X(_03657_));
 sky130_fd_sc_hd__a21boi_2 _10571_ (.A1(_03532_),
    .A2(_03612_),
    .B1_N(_03611_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_2 _10572_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03609_),
    .Y(_03659_));
 sky130_fd_sc_hd__o22a_1 _10573_ (.A1(net76),
    .A2(net23),
    .B1(net15),
    .B2(net72),
    .X(_03660_));
 sky130_fd_sc_hd__xnor2_2 _10574_ (.A(net68),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__a22o_1 _10575_ (.A1(net102),
    .A2(net38),
    .B1(net36),
    .B2(_00174_),
    .X(_03662_));
 sky130_fd_sc_hd__xor2_1 _10576_ (.A(net90),
    .B(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__inv_2 _10577_ (.A(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__xnor2_1 _10578_ (.A(_03661_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__a22o_1 _10579_ (.A1(net42),
    .A2(_00334_),
    .B1(_00340_),
    .B2(net41),
    .X(_03666_));
 sky130_fd_sc_hd__xor2_1 _10580_ (.A(net92),
    .B(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__nand2b_1 _10581_ (.A_N(_03665_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand2b_1 _10582_ (.A_N(_03667_),
    .B(_03665_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _10583_ (.A(_03668_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__a21boi_2 _10584_ (.A1(_03552_),
    .A2(_03558_),
    .B1_N(_03557_),
    .Y(_03671_));
 sky130_fd_sc_hd__o22a_1 _10585_ (.A1(net120),
    .A2(net10),
    .B1(net5),
    .B2(net116),
    .X(_03672_));
 sky130_fd_sc_hd__xnor2_2 _10586_ (.A(net19),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__xnor2_2 _10587_ (.A(_03671_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__nor2_1 _10588_ (.A(net111),
    .B(net19),
    .Y(_03675_));
 sky130_fd_sc_hd__or3_1 _10589_ (.A(net111),
    .B(net19),
    .C(_03674_),
    .X(_03676_));
 sky130_fd_sc_hd__xnor2_2 _10590_ (.A(_03674_),
    .B(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__o22a_1 _10591_ (.A1(net53),
    .A2(net46),
    .B1(net44),
    .B2(net51),
    .X(_03678_));
 sky130_fd_sc_hd__xnor2_2 _10592_ (.A(net96),
    .B(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__o22a_1 _10593_ (.A1(net59),
    .A2(net27),
    .B1(net25),
    .B2(net56),
    .X(_03680_));
 sky130_fd_sc_hd__xnor2_2 _10594_ (.A(net88),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__and2_1 _10595_ (.A(_03679_),
    .B(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__xor2_2 _10596_ (.A(_03679_),
    .B(_03681_),
    .X(_03683_));
 sky130_fd_sc_hd__a22o_1 _10597_ (.A1(_06515_),
    .A2(net31),
    .B1(net29),
    .B2(_06522_),
    .X(_03684_));
 sky130_fd_sc_hd__xnor2_2 _10598_ (.A(net49),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__xor2_2 _10599_ (.A(_03683_),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__nand2_1 _10600_ (.A(_03677_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__xnor2_2 _10601_ (.A(_03677_),
    .B(_03686_),
    .Y(_03688_));
 sky130_fd_sc_hd__xor2_2 _10602_ (.A(_03670_),
    .B(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__a21o_1 _10603_ (.A1(_03589_),
    .A2(_03591_),
    .B1(_03587_),
    .X(_03690_));
 sky130_fd_sc_hd__a21o_1 _10604_ (.A1(_00381_),
    .A2(net8),
    .B1(_00327_),
    .X(_03691_));
 sky130_fd_sc_hd__o31a_2 _10605_ (.A1(_00328_),
    .A2(_00377_),
    .A3(net7),
    .B1(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__xnor2_1 _10606_ (.A(_03690_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__a21oi_1 _10607_ (.A1(_03538_),
    .A2(_03542_),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__and3_1 _10608_ (.A(_03538_),
    .B(_03542_),
    .C(_03693_),
    .X(_03695_));
 sky130_fd_sc_hd__nor2_1 _10609_ (.A(_03694_),
    .B(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__xnor2_2 _10610_ (.A(_03689_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__o21ba_1 _10611_ (.A1(_03430_),
    .A2(_03580_),
    .B1_N(_03579_),
    .X(_03698_));
 sky130_fd_sc_hd__o22a_1 _10612_ (.A1(net82),
    .A2(net13),
    .B1(net12),
    .B2(_00333_),
    .X(_03699_));
 sky130_fd_sc_hd__xnor2_2 _10613_ (.A(_00323_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__o22a_1 _10614_ (.A1(net66),
    .A2(net35),
    .B1(net33),
    .B2(net64),
    .X(_03701_));
 sky130_fd_sc_hd__xnor2_1 _10615_ (.A(net124),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__nor2_1 _10616_ (.A(_03700_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__xnor2_1 _10617_ (.A(_03700_),
    .B(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__o22a_1 _10618_ (.A1(net54),
    .A2(net74),
    .B1(net16),
    .B2(net78),
    .X(_03705_));
 sky130_fd_sc_hd__xnor2_1 _10619_ (.A(net122),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__nor2_1 _10620_ (.A(_03704_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__and2_1 _10621_ (.A(_03704_),
    .B(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__or2_1 _10622_ (.A(_03707_),
    .B(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__a21oi_1 _10623_ (.A1(_03572_),
    .A2(_03575_),
    .B1(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__and3_1 _10624_ (.A(_03572_),
    .B(_03575_),
    .C(_03709_),
    .X(_03711_));
 sky130_fd_sc_hd__nor2_1 _10625_ (.A(_03710_),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__xnor2_2 _10626_ (.A(_03698_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__and2b_1 _10627_ (.A_N(_03697_),
    .B(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__xnor2_2 _10628_ (.A(_03697_),
    .B(_03713_),
    .Y(_03715_));
 sky130_fd_sc_hd__a21bo_1 _10629_ (.A1(_03549_),
    .A2(_03596_),
    .B1_N(_03595_),
    .X(_03716_));
 sky130_fd_sc_hd__a21o_1 _10630_ (.A1(_03601_),
    .A2(_03605_),
    .B1(_03604_),
    .X(_03717_));
 sky130_fd_sc_hd__o21ai_2 _10631_ (.A1(_03550_),
    .A2(_03563_),
    .B1(_03562_),
    .Y(_03718_));
 sky130_fd_sc_hd__a32o_1 _10632_ (.A1(_03575_),
    .A2(_03576_),
    .A3(_03593_),
    .B1(_03592_),
    .B2(_03582_),
    .X(_03719_));
 sky130_fd_sc_hd__xor2_1 _10633_ (.A(_03718_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__o21ai_1 _10634_ (.A1(_03545_),
    .A2(_03548_),
    .B1(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__or3_1 _10635_ (.A(_03545_),
    .B(_03548_),
    .C(_03720_),
    .X(_03722_));
 sky130_fd_sc_hd__and2_1 _10636_ (.A(_03721_),
    .B(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__xnor2_2 _10637_ (.A(_03717_),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2b_1 _10638_ (.A_N(_03724_),
    .B(_03716_),
    .Y(_03725_));
 sky130_fd_sc_hd__xnor2_2 _10639_ (.A(_03716_),
    .B(_03724_),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2_1 _10640_ (.A(_03715_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__xnor2_2 _10641_ (.A(_03715_),
    .B(_03726_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand2b_1 _10642_ (.A_N(_03728_),
    .B(_03659_),
    .Y(_03729_));
 sky130_fd_sc_hd__xor2_2 _10643_ (.A(_03659_),
    .B(_03728_),
    .X(_03730_));
 sky130_fd_sc_hd__or2_2 _10644_ (.A(_03658_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__nand2_1 _10645_ (.A(_03658_),
    .B(_03730_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_4 _10646_ (.A(_03731_),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__a21oi_1 _10647_ (.A1(_03492_),
    .A2(_03615_),
    .B1(_03616_),
    .Y(_03734_));
 sky130_fd_sc_hd__nor2_1 _10648_ (.A(_03494_),
    .B(_03617_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21oi_1 _10649_ (.A1(_03405_),
    .A2(_03735_),
    .B1(_03734_),
    .Y(_03736_));
 sky130_fd_sc_hd__or4_1 _10650_ (.A(_03218_),
    .B(_03355_),
    .C(_03494_),
    .D(_03617_),
    .X(_03737_));
 sky130_fd_sc_hd__o21bai_1 _10651_ (.A1(_03222_),
    .A2(_03223_),
    .B1_N(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__o311a_4 _10652_ (.A1(_02643_),
    .A2(_03219_),
    .A3(_03737_),
    .B1(_03738_),
    .C1(_03736_),
    .X(_03739_));
 sky130_fd_sc_hd__xor2_4 _10653_ (.A(_03733_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__a21oi_1 _10654_ (.A1(net159),
    .A2(_03657_),
    .B1(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__a31o_1 _10655_ (.A1(net159),
    .A2(_03657_),
    .A3(_03740_),
    .B1(net187),
    .X(_03742_));
 sky130_fd_sc_hd__nand2_1 _10656_ (.A(net159),
    .B(_01821_),
    .Y(_03743_));
 sky130_fd_sc_hd__xnor2_1 _10657_ (.A(_01825_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__o21ai_1 _10658_ (.A1(_06205_),
    .A2(_03630_),
    .B1(_06214_),
    .Y(_03745_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(_06361_),
    .A1(_03745_),
    .S(net285),
    .X(_03746_));
 sky130_fd_sc_hd__nor2_1 _10660_ (.A(_06169_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__a21o_1 _10661_ (.A1(_06169_),
    .A2(_03746_),
    .B1(net236),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _10662_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03749_));
 sky130_fd_sc_hd__or2_1 _10663_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03750_));
 sky130_fd_sc_hd__o21ai_2 _10664_ (.A1(_03634_),
    .A2(_03635_),
    .B1(_03636_),
    .Y(_03751_));
 sky130_fd_sc_hd__a21oi_1 _10665_ (.A1(_03749_),
    .A2(_03750_),
    .B1(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__and3_1 _10666_ (.A(_03749_),
    .B(_03750_),
    .C(_03751_),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(_02661_),
    .A1(_02667_),
    .S(net217),
    .X(_03754_));
 sky130_fd_sc_hd__inv_2 _10668_ (.A(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(_03101_),
    .A1(_03755_),
    .S(_06318_),
    .X(_03756_));
 sky130_fd_sc_hd__o21a_1 _10670_ (.A1(_03752_),
    .A2(_03753_),
    .B1(net250),
    .X(_03757_));
 sky130_fd_sc_hd__a211o_1 _10671_ (.A1(net224),
    .A2(_03756_),
    .B1(_03757_),
    .C1(net196),
    .X(_03758_));
 sky130_fd_sc_hd__or2_1 _10672_ (.A(\div_res[9] ),
    .B(_03642_),
    .X(_03759_));
 sky130_fd_sc_hd__a21oi_1 _10673_ (.A1(net165),
    .A2(_03759_),
    .B1(\div_res[10] ),
    .Y(_03760_));
 sky130_fd_sc_hd__a31o_1 _10674_ (.A1(\div_res[10] ),
    .A2(net165),
    .A3(_03759_),
    .B1(net183),
    .X(_03761_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(net234),
    .A1(net185),
    .S(_06160_),
    .X(_03762_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(net186),
    .A2(_03762_),
    .B1(_06154_),
    .X(_03763_));
 sky130_fd_sc_hd__or2_1 _10677_ (.A(\div_shifter[41] ),
    .B(_03646_),
    .X(_03764_));
 sky130_fd_sc_hd__a21oi_1 _10678_ (.A1(net228),
    .A2(_03764_),
    .B1(\div_shifter[42] ),
    .Y(_03765_));
 sky130_fd_sc_hd__a31o_1 _10679_ (.A1(\div_shifter[42] ),
    .A2(net228),
    .A3(_03764_),
    .B1(net231),
    .X(_03766_));
 sky130_fd_sc_hd__o2bb2a_1 _10680_ (.A1_N(_06148_),
    .A2_N(net242),
    .B1(_03765_),
    .B2(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__o211a_1 _10681_ (.A1(_03760_),
    .A2(_03761_),
    .B1(_03763_),
    .C1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__o21ai_2 _10682_ (.A1(net221),
    .A2(_03107_),
    .B1(_02342_),
    .Y(_03769_));
 sky130_fd_sc_hd__o221a_1 _10683_ (.A1(_02320_),
    .A2(_03756_),
    .B1(_03769_),
    .B2(net168),
    .C1(_03768_),
    .X(_03770_));
 sky130_fd_sc_hd__o211a_1 _10684_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03758_),
    .C1(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__o221a_1 _10685_ (.A1(_03741_),
    .A2(_03742_),
    .B1(_03744_),
    .B2(_02330_),
    .C1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__and3_1 _10686_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(_03527_),
    .X(_03773_));
 sky130_fd_sc_hd__a21oi_1 _10687_ (.A1(curr_PC[9]),
    .A2(_03527_),
    .B1(curr_PC[10]),
    .Y(_03774_));
 sky130_fd_sc_hd__or3_2 _10688_ (.A(net243),
    .B(_03773_),
    .C(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__o21ai_4 _10689_ (.A1(net248),
    .A2(_03772_),
    .B1(_03775_),
    .Y(dest_val[10]));
 sky130_fd_sc_hd__o21a_1 _10690_ (.A1(_03657_),
    .A2(_03740_),
    .B1(net159),
    .X(_03776_));
 sky130_fd_sc_hd__a21bo_1 _10691_ (.A1(_03717_),
    .A2(_03723_),
    .B1_N(_03725_),
    .X(_03777_));
 sky130_fd_sc_hd__a21oi_1 _10692_ (.A1(_03683_),
    .A2(_03685_),
    .B1(_03682_),
    .Y(_03778_));
 sky130_fd_sc_hd__or2_1 _10693_ (.A(_03692_),
    .B(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__xor2_1 _10694_ (.A(_03692_),
    .B(_03778_),
    .X(_03780_));
 sky130_fd_sc_hd__o21ai_1 _10695_ (.A1(_03703_),
    .A2(_03707_),
    .B1(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__or3_1 _10696_ (.A(_03703_),
    .B(_03707_),
    .C(_03780_),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_03781_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__o22a_1 _10698_ (.A1(net61),
    .A2(net46),
    .B1(net44),
    .B2(net53),
    .X(_03784_));
 sky130_fd_sc_hd__xnor2_1 _10699_ (.A(net96),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__a22o_1 _10700_ (.A1(_00174_),
    .A2(net42),
    .B1(net41),
    .B2(_00334_),
    .X(_03786_));
 sky130_fd_sc_hd__xor2_1 _10701_ (.A(net92),
    .B(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__xor2_1 _10702_ (.A(_03785_),
    .B(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a22o_1 _10703_ (.A1(_00157_),
    .A2(net38),
    .B1(net36),
    .B2(net102),
    .X(_03789_));
 sky130_fd_sc_hd__xor2_1 _10704_ (.A(net90),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__and2_1 _10705_ (.A(_03788_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_1 _10706_ (.A(_03788_),
    .B(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__or2_1 _10707_ (.A(_03791_),
    .B(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__o22a_1 _10708_ (.A1(net72),
    .A2(net9),
    .B1(net4),
    .B2(net120),
    .X(_03794_));
 sky130_fd_sc_hd__xnor2_1 _10709_ (.A(net19),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__a32o_1 _10710_ (.A1(_00347_),
    .A2(_00676_),
    .A3(_00677_),
    .B1(_00442_),
    .B2(_00340_),
    .X(_03796_));
 sky130_fd_sc_hd__xnor2_2 _10711_ (.A(_00668_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _10712_ (.A(net115),
    .B(net21),
    .Y(_03798_));
 sky130_fd_sc_hd__xor2_1 _10713_ (.A(_03797_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2b_1 _10714_ (.A_N(_03795_),
    .B(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__xnor2_1 _10715_ (.A(_03795_),
    .B(_03799_),
    .Y(_03801_));
 sky130_fd_sc_hd__o22a_1 _10716_ (.A1(net54),
    .A2(net35),
    .B1(net33),
    .B2(net66),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _10717_ (.A(net126),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__a22o_1 _10718_ (.A1(_06538_),
    .A2(net31),
    .B1(net29),
    .B2(_06515_),
    .X(_03804_));
 sky130_fd_sc_hd__xnor2_1 _10719_ (.A(net49),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__and2_1 _10720_ (.A(_03803_),
    .B(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__xor2_1 _10721_ (.A(_03803_),
    .B(_03805_),
    .X(_03807_));
 sky130_fd_sc_hd__o22a_1 _10722_ (.A1(net64),
    .A2(net27),
    .B1(net25),
    .B2(net59),
    .X(_03808_));
 sky130_fd_sc_hd__xnor2_1 _10723_ (.A(net88),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__xor2_1 _10724_ (.A(_03807_),
    .B(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__nand2_1 _10725_ (.A(_03801_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__or2_1 _10726_ (.A(_03801_),
    .B(_03810_),
    .X(_03812_));
 sky130_fd_sc_hd__nand2_1 _10727_ (.A(_03811_),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__xnor2_1 _10728_ (.A(_03793_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__xnor2_1 _10729_ (.A(_03783_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__o21ai_1 _10730_ (.A1(_03671_),
    .A2(_03673_),
    .B1(_03676_),
    .Y(_03816_));
 sky130_fd_sc_hd__o22a_1 _10731_ (.A1(net82),
    .A2(net12),
    .B1(net6),
    .B2(net86),
    .X(_03817_));
 sky130_fd_sc_hd__xnor2_1 _10732_ (.A(_00324_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__o22a_1 _10733_ (.A1(net74),
    .A2(_00399_),
    .B1(net13),
    .B2(net78),
    .X(_03819_));
 sky130_fd_sc_hd__xnor2_1 _10734_ (.A(net122),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__nor2_1 _10735_ (.A(_00328_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__xnor2_1 _10736_ (.A(_00327_),
    .B(_03820_),
    .Y(_03822_));
 sky130_fd_sc_hd__and2_1 _10737_ (.A(_03818_),
    .B(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__nor2_1 _10738_ (.A(_03818_),
    .B(_03822_),
    .Y(_03824_));
 sky130_fd_sc_hd__nor2_1 _10739_ (.A(_03823_),
    .B(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__o21ai_2 _10740_ (.A1(_03661_),
    .A2(_03664_),
    .B1(_03668_),
    .Y(_03826_));
 sky130_fd_sc_hd__and2_1 _10741_ (.A(_03825_),
    .B(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__xor2_1 _10742_ (.A(_03825_),
    .B(_03826_),
    .X(_03828_));
 sky130_fd_sc_hd__xnor2_1 _10743_ (.A(_03816_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__or2_1 _10744_ (.A(_03815_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_03815_),
    .B(_03829_),
    .Y(_03831_));
 sky130_fd_sc_hd__and2_1 _10746_ (.A(_03830_),
    .B(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__a21o_1 _10747_ (.A1(_03689_),
    .A2(_03696_),
    .B1(_03714_),
    .X(_03833_));
 sky130_fd_sc_hd__o21bai_2 _10748_ (.A1(_03698_),
    .A2(_03711_),
    .B1_N(_03710_),
    .Y(_03834_));
 sky130_fd_sc_hd__o21a_1 _10749_ (.A1(_03670_),
    .A2(_03688_),
    .B1(_03687_),
    .X(_03835_));
 sky130_fd_sc_hd__a21o_1 _10750_ (.A1(_03690_),
    .A2(_03692_),
    .B1(_03694_),
    .X(_03836_));
 sky130_fd_sc_hd__nand2b_1 _10751_ (.A_N(_03835_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__xnor2_2 _10752_ (.A(_03835_),
    .B(_03836_),
    .Y(_03838_));
 sky130_fd_sc_hd__xnor2_2 _10753_ (.A(_03834_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__a21boi_2 _10754_ (.A1(_03718_),
    .A2(_03719_),
    .B1_N(_03721_),
    .Y(_03840_));
 sky130_fd_sc_hd__xnor2_2 _10755_ (.A(_03839_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2b_1 _10756_ (.A_N(_03841_),
    .B(_03833_),
    .Y(_03842_));
 sky130_fd_sc_hd__xnor2_2 _10757_ (.A(_03833_),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _10758_ (.A(_03832_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__xnor2_1 _10759_ (.A(_03832_),
    .B(_03843_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2b_1 _10760_ (.A_N(_03845_),
    .B(_03777_),
    .Y(_03846_));
 sky130_fd_sc_hd__xor2_1 _10761_ (.A(_03777_),
    .B(_03845_),
    .X(_03847_));
 sky130_fd_sc_hd__a21oi_1 _10762_ (.A1(_03727_),
    .A2(_03729_),
    .B1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__a21o_1 _10763_ (.A1(_03727_),
    .A2(_03729_),
    .B1(_03847_),
    .X(_03849_));
 sky130_fd_sc_hd__and3_1 _10764_ (.A(_03727_),
    .B(_03729_),
    .C(_03847_),
    .X(_03850_));
 sky130_fd_sc_hd__or2_2 _10765_ (.A(_03848_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__a21boi_2 _10766_ (.A1(_03615_),
    .A2(_03731_),
    .B1_N(_03732_),
    .Y(_03852_));
 sky130_fd_sc_hd__nor2_2 _10767_ (.A(_03617_),
    .B(_03733_),
    .Y(_03853_));
 sky130_fd_sc_hd__a21oi_1 _10768_ (.A1(_03618_),
    .A2(_03853_),
    .B1(_03852_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand2_1 _10769_ (.A(_03619_),
    .B(_03853_),
    .Y(_03855_));
 sky130_fd_sc_hd__o211ai_1 _10770_ (.A1(_03358_),
    .A2(_03359_),
    .B1(_03619_),
    .C1(_03853_),
    .Y(_03856_));
 sky130_fd_sc_hd__o311a_4 _10771_ (.A1(_02803_),
    .A2(_03357_),
    .A3(_03855_),
    .B1(_03856_),
    .C1(_03854_),
    .X(_03857_));
 sky130_fd_sc_hd__xor2_4 _10772_ (.A(_03851_),
    .B(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_1 _10773_ (.A(_03776_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__or2_1 _10774_ (.A(_03776_),
    .B(_03858_),
    .X(_03860_));
 sky130_fd_sc_hd__a31o_1 _10775_ (.A1(_01818_),
    .A2(_01820_),
    .A3(_01825_),
    .B1(net157),
    .X(_03861_));
 sky130_fd_sc_hd__xor2_1 _10776_ (.A(_01827_),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__a21o_1 _10777_ (.A1(_06169_),
    .A2(_03745_),
    .B1(_06160_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(_06363_),
    .A1(_03863_),
    .S(net285),
    .X(_03864_));
 sky130_fd_sc_hd__nand2_1 _10779_ (.A(_06136_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__o211a_1 _10780_ (.A1(_06136_),
    .A2(_03864_),
    .B1(_03865_),
    .C1(_02323_),
    .X(_03866_));
 sky130_fd_sc_hd__nand2_1 _10781_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .Y(_03867_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03868_));
 sky130_fd_sc_hd__a21bo_1 _10783_ (.A1(_03750_),
    .A2(_03751_),
    .B1_N(_03749_),
    .X(_03869_));
 sky130_fd_sc_hd__a21o_1 _10784_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__and3_1 _10785_ (.A(_03867_),
    .B(_03868_),
    .C(_03869_),
    .X(_03871_));
 sky130_fd_sc_hd__or3b_1 _10786_ (.A(_03871_),
    .B(net223),
    .C_N(_03870_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(_02814_),
    .A1(_02820_),
    .S(net217),
    .X(_03873_));
 sky130_fd_sc_hd__inv_2 _10788_ (.A(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(_02967_),
    .A1(_03874_),
    .S(_06318_),
    .X(_03875_));
 sky130_fd_sc_hd__o21a_1 _10790_ (.A1(net250),
    .A2(_03875_),
    .B1(_03872_),
    .X(_03876_));
 sky130_fd_sc_hd__or2_1 _10791_ (.A(\div_res[10] ),
    .B(_03759_),
    .X(_03877_));
 sky130_fd_sc_hd__a21oi_1 _10792_ (.A1(net165),
    .A2(_03877_),
    .B1(\div_res[11] ),
    .Y(_03878_));
 sky130_fd_sc_hd__a311o_1 _10793_ (.A1(\div_res[11] ),
    .A2(net165),
    .A3(_03877_),
    .B1(_03878_),
    .C1(net183),
    .X(_03879_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(net234),
    .A1(net185),
    .S(_06124_),
    .X(_03880_));
 sky130_fd_sc_hd__a21o_1 _10795_ (.A1(net186),
    .A2(_03880_),
    .B1(_06130_),
    .X(_03881_));
 sky130_fd_sc_hd__or2_1 _10796_ (.A(\div_shifter[42] ),
    .B(_03764_),
    .X(_03882_));
 sky130_fd_sc_hd__a21oi_1 _10797_ (.A1(net228),
    .A2(_03882_),
    .B1(\div_shifter[43] ),
    .Y(_03883_));
 sky130_fd_sc_hd__a31o_1 _10798_ (.A1(\div_shifter[43] ),
    .A2(net228),
    .A3(_03882_),
    .B1(net231),
    .X(_03884_));
 sky130_fd_sc_hd__o2bb2a_1 _10799_ (.A1_N(_06118_),
    .A2_N(net242),
    .B1(_03883_),
    .B2(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__and3_1 _10800_ (.A(_03879_),
    .B(_03881_),
    .C(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__o21ai_2 _10801_ (.A1(net220),
    .A2(_02973_),
    .B1(_02342_),
    .Y(_03887_));
 sky130_fd_sc_hd__o221a_1 _10802_ (.A1(_02320_),
    .A2(_03875_),
    .B1(_03887_),
    .B2(_02250_),
    .C1(_03886_),
    .X(_03888_));
 sky130_fd_sc_hd__o21ai_1 _10803_ (.A1(net196),
    .A2(_03876_),
    .B1(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__a211o_1 _10804_ (.A1(net233),
    .A2(_03862_),
    .B1(_03866_),
    .C1(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__a31o_1 _10805_ (.A1(_02245_),
    .A2(_03859_),
    .A3(_03860_),
    .B1(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__or2_1 _10806_ (.A(curr_PC[11]),
    .B(_03773_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _10807_ (.A(curr_PC[11]),
    .B(_03773_),
    .X(_03893_));
 sky130_fd_sc_hd__nor2_1 _10808_ (.A(net243),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__a22o_4 _10809_ (.A1(net243),
    .A2(_03891_),
    .B1(_03892_),
    .B2(_03894_),
    .X(dest_val[11]));
 sky130_fd_sc_hd__nor2_1 _10810_ (.A(_03740_),
    .B(_03858_),
    .Y(_03895_));
 sky130_fd_sc_hd__and2b_1 _10811_ (.A_N(_03657_),
    .B(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__or2_1 _10812_ (.A(net157),
    .B(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__o21ai_2 _10813_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03842_),
    .Y(_03898_));
 sky130_fd_sc_hd__o21ai_1 _10814_ (.A1(_03797_),
    .A2(_03798_),
    .B1(_03800_),
    .Y(_03899_));
 sky130_fd_sc_hd__a21o_1 _10815_ (.A1(_03785_),
    .A2(_03787_),
    .B1(_03791_),
    .X(_03900_));
 sky130_fd_sc_hd__o22a_1 _10816_ (.A1(net74),
    .A2(net13),
    .B1(net12),
    .B2(net78),
    .X(_03901_));
 sky130_fd_sc_hd__xnor2_2 _10817_ (.A(net122),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__inv_2 _10818_ (.A(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_1 _10819_ (.A1(_00331_),
    .A2(net6),
    .B1(_00324_),
    .Y(_03904_));
 sky130_fd_sc_hd__o31ai_2 _10820_ (.A1(_00324_),
    .A2(_00332_),
    .A3(net6),
    .B1(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__nor2_1 _10821_ (.A(_03903_),
    .B(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__xnor2_1 _10822_ (.A(_03902_),
    .B(_03905_),
    .Y(_03907_));
 sky130_fd_sc_hd__inv_2 _10823_ (.A(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__xnor2_1 _10824_ (.A(_03900_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand2b_1 _10825_ (.A_N(_03909_),
    .B(_03899_),
    .Y(_03910_));
 sky130_fd_sc_hd__xnor2_1 _10826_ (.A(_03899_),
    .B(_03909_),
    .Y(_03911_));
 sky130_fd_sc_hd__a22o_1 _10827_ (.A1(net102),
    .A2(net43),
    .B1(net41),
    .B2(_00174_),
    .X(_03912_));
 sky130_fd_sc_hd__xor2_1 _10828_ (.A(net92),
    .B(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__o22a_1 _10829_ (.A1(net63),
    .A2(net46),
    .B1(net44),
    .B2(net61),
    .X(_03914_));
 sky130_fd_sc_hd__xnor2_1 _10830_ (.A(net96),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__and2_1 _10831_ (.A(_03913_),
    .B(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__nor2_1 _10832_ (.A(_03913_),
    .B(_03915_),
    .Y(_03917_));
 sky130_fd_sc_hd__nor2_1 _10833_ (.A(_03916_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a22o_1 _10834_ (.A1(_00148_),
    .A2(net38),
    .B1(net36),
    .B2(_00157_),
    .X(_03919_));
 sky130_fd_sc_hd__xor2_1 _10835_ (.A(net90),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__xnor2_1 _10836_ (.A(_03918_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__o32a_1 _10837_ (.A1(net35),
    .A2(_00395_),
    .A3(_00397_),
    .B1(net33),
    .B2(net54),
    .X(_03922_));
 sky130_fd_sc_hd__xnor2_2 _10838_ (.A(net126),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__a22o_1 _10839_ (.A1(_06534_),
    .A2(net31),
    .B1(net29),
    .B2(_06538_),
    .X(_03924_));
 sky130_fd_sc_hd__xnor2_1 _10840_ (.A(net49),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _10841_ (.A(_03923_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__xor2_1 _10842_ (.A(_03923_),
    .B(_03925_),
    .X(_03927_));
 sky130_fd_sc_hd__o22a_1 _10843_ (.A1(net66),
    .A2(net27),
    .B1(net25),
    .B2(net64),
    .X(_03928_));
 sky130_fd_sc_hd__xnor2_1 _10844_ (.A(net88),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _10845_ (.A(_03927_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__xor2_1 _10846_ (.A(_03927_),
    .B(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__o22a_1 _10847_ (.A1(net84),
    .A2(net23),
    .B1(net15),
    .B2(net80),
    .X(_03932_));
 sky130_fd_sc_hd__xnor2_1 _10848_ (.A(net69),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__o22a_1 _10849_ (.A1(net76),
    .A2(net9),
    .B1(net4),
    .B2(net72),
    .X(_03934_));
 sky130_fd_sc_hd__xnor2_1 _10850_ (.A(net19),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__or2_1 _10851_ (.A(_03933_),
    .B(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__xor2_1 _10852_ (.A(_03933_),
    .B(_03935_),
    .X(_03937_));
 sky130_fd_sc_hd__nand2_1 _10853_ (.A(_03931_),
    .B(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__xnor2_1 _10854_ (.A(_03931_),
    .B(_03937_),
    .Y(_03939_));
 sky130_fd_sc_hd__or2_1 _10855_ (.A(_03921_),
    .B(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__nand2_1 _10856_ (.A(_03921_),
    .B(_03939_),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _10857_ (.A(_03940_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__a21oi_1 _10858_ (.A1(_03807_),
    .A2(_03809_),
    .B1(_03806_),
    .Y(_03943_));
 sky130_fd_sc_hd__nor2_1 _10859_ (.A(net120),
    .B(net19),
    .Y(_03944_));
 sky130_fd_sc_hd__xnor2_1 _10860_ (.A(_03943_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__o21ai_1 _10861_ (.A1(_03821_),
    .A2(_03823_),
    .B1(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__or3_1 _10862_ (.A(_03821_),
    .B(_03823_),
    .C(_03945_),
    .X(_03947_));
 sky130_fd_sc_hd__nand2_1 _10863_ (.A(_03946_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__xor2_1 _10864_ (.A(_03942_),
    .B(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_1 _10865_ (.A(_03911_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__or2_1 _10866_ (.A(_03911_),
    .B(_03949_),
    .X(_03951_));
 sky130_fd_sc_hd__and2_1 _10867_ (.A(_03950_),
    .B(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__o21a_1 _10868_ (.A1(_03783_),
    .A2(_03814_),
    .B1(_03830_),
    .X(_03953_));
 sky130_fd_sc_hd__a21o_1 _10869_ (.A1(_03816_),
    .A2(_03828_),
    .B1(_03827_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_1 _10870_ (.A(_03779_),
    .B(_03781_),
    .Y(_03955_));
 sky130_fd_sc_hd__o21a_1 _10871_ (.A1(_03793_),
    .A2(_03813_),
    .B1(_03811_),
    .X(_03956_));
 sky130_fd_sc_hd__a21oi_1 _10872_ (.A1(_03779_),
    .A2(_03781_),
    .B1(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__xnor2_2 _10873_ (.A(_03955_),
    .B(_03956_),
    .Y(_03958_));
 sky130_fd_sc_hd__xnor2_2 _10874_ (.A(_03954_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__a21boi_2 _10875_ (.A1(_03834_),
    .A2(_03838_),
    .B1_N(_03837_),
    .Y(_03960_));
 sky130_fd_sc_hd__xor2_2 _10876_ (.A(_03959_),
    .B(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__nand2b_1 _10877_ (.A_N(_03953_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__xnor2_2 _10878_ (.A(_03953_),
    .B(_03961_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _10879_ (.A(_03952_),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__xor2_2 _10880_ (.A(_03952_),
    .B(_03963_),
    .X(_03965_));
 sky130_fd_sc_hd__nand2_1 _10881_ (.A(_03898_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__xnor2_2 _10882_ (.A(_03898_),
    .B(_03965_),
    .Y(_03967_));
 sky130_fd_sc_hd__a21oi_1 _10883_ (.A1(_03844_),
    .A2(_03846_),
    .B1(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__a21o_1 _10884_ (.A1(_03844_),
    .A2(_03846_),
    .B1(_03967_),
    .X(_03969_));
 sky130_fd_sc_hd__and3_1 _10885_ (.A(_03844_),
    .B(_03846_),
    .C(_03967_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_2 _10886_ (.A(_03968_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__a21oi_1 _10887_ (.A1(_03731_),
    .A2(_03849_),
    .B1(_03850_),
    .Y(_03972_));
 sky130_fd_sc_hd__nor2_1 _10888_ (.A(_03733_),
    .B(_03851_),
    .Y(_03973_));
 sky130_fd_sc_hd__a21o_1 _10889_ (.A1(_03734_),
    .A2(_03973_),
    .B1(_03972_),
    .X(_03974_));
 sky130_fd_sc_hd__and2_1 _10890_ (.A(_03735_),
    .B(_03973_),
    .X(_03975_));
 sky130_fd_sc_hd__a21o_1 _10891_ (.A1(_03410_),
    .A2(_03975_),
    .B1(_03974_),
    .X(_03976_));
 sky130_fd_sc_hd__xor2_4 _10892_ (.A(_03971_),
    .B(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__o21ai_1 _10893_ (.A1(_03897_),
    .A2(_03977_),
    .B1(_02245_),
    .Y(_03978_));
 sky130_fd_sc_hd__a21oi_1 _10894_ (.A1(_03897_),
    .A2(_03977_),
    .B1(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21bo_1 _10895_ (.A1(net159),
    .A2(_01828_),
    .B1_N(_01831_),
    .X(_03980_));
 sky130_fd_sc_hd__or3b_1 _10896_ (.A(net157),
    .B(_01831_),
    .C_N(_01828_),
    .X(_03981_));
 sky130_fd_sc_hd__a21o_1 _10897_ (.A1(_06136_),
    .A2(_03863_),
    .B1(_06124_),
    .X(_03982_));
 sky130_fd_sc_hd__nand2_1 _10898_ (.A(net285),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__o21ai_1 _10899_ (.A1(net285),
    .A2(_06365_),
    .B1(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__o21ai_1 _10900_ (.A1(_06100_),
    .A2(_03984_),
    .B1(_02323_),
    .Y(_03985_));
 sky130_fd_sc_hd__a21o_1 _10901_ (.A1(_06100_),
    .A2(_03984_),
    .B1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__or2_1 _10902_ (.A(net219),
    .B(_02972_),
    .X(_03987_));
 sky130_fd_sc_hd__o211a_1 _10903_ (.A1(net217),
    .A2(_02970_),
    .B1(_03987_),
    .C1(_06318_),
    .X(_03988_));
 sky130_fd_sc_hd__a21oi_2 _10904_ (.A1(net220),
    .A2(_02831_),
    .B1(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_03990_));
 sky130_fd_sc_hd__or2_1 _10906_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_03991_));
 sky130_fd_sc_hd__a21bo_1 _10907_ (.A1(_03868_),
    .A2(_03869_),
    .B1_N(_03867_),
    .X(_03992_));
 sky130_fd_sc_hd__and3_1 _10908_ (.A(_03990_),
    .B(_03991_),
    .C(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__a21o_1 _10909_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03992_),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _10910_ (.A(net250),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__o22a_1 _10911_ (.A1(net250),
    .A2(_03989_),
    .B1(_03993_),
    .B2(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _10912_ (.A(\div_res[11] ),
    .B(_03877_),
    .X(_03997_));
 sky130_fd_sc_hd__a21oi_1 _10913_ (.A1(net165),
    .A2(_03997_),
    .B1(\div_res[12] ),
    .Y(_03998_));
 sky130_fd_sc_hd__a311o_1 _10914_ (.A1(\div_res[12] ),
    .A2(net165),
    .A3(_03997_),
    .B1(_03998_),
    .C1(net183),
    .X(_03999_));
 sky130_fd_sc_hd__or2_1 _10915_ (.A(\div_shifter[43] ),
    .B(_03882_),
    .X(_04000_));
 sky130_fd_sc_hd__a21oi_1 _10916_ (.A1(net228),
    .A2(_04000_),
    .B1(\div_shifter[44] ),
    .Y(_04001_));
 sky130_fd_sc_hd__a311o_1 _10917_ (.A1(\div_shifter[44] ),
    .A2(net228),
    .A3(_04000_),
    .B1(_04001_),
    .C1(net231),
    .X(_04002_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(net234),
    .A1(net185),
    .S(_06088_),
    .X(_04003_));
 sky130_fd_sc_hd__a21oi_1 _10919_ (.A1(net186),
    .A2(_04003_),
    .B1(_06094_),
    .Y(_04004_));
 sky130_fd_sc_hd__a21oi_1 _10920_ (.A1(_06081_),
    .A2(net242),
    .B1(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__and3_1 _10921_ (.A(_03999_),
    .B(_04002_),
    .C(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__o21ai_2 _10922_ (.A1(net220),
    .A2(_02821_),
    .B1(_02342_),
    .Y(_04007_));
 sky130_fd_sc_hd__o221a_1 _10923_ (.A1(_02320_),
    .A2(_03989_),
    .B1(_04007_),
    .B2(net168),
    .C1(_04006_),
    .X(_04008_));
 sky130_fd_sc_hd__o211ai_2 _10924_ (.A1(net196),
    .A2(_03996_),
    .B1(_04008_),
    .C1(_03986_),
    .Y(_04009_));
 sky130_fd_sc_hd__a311o_1 _10925_ (.A1(net233),
    .A2(_03980_),
    .A3(_03981_),
    .B1(_04009_),
    .C1(_03979_),
    .X(_04010_));
 sky130_fd_sc_hd__and3_2 _10926_ (.A(curr_PC[11]),
    .B(curr_PC[12]),
    .C(_03773_),
    .X(_04011_));
 sky130_fd_sc_hd__o21ai_1 _10927_ (.A1(curr_PC[12]),
    .A2(_03893_),
    .B1(net248),
    .Y(_04012_));
 sky130_fd_sc_hd__a2bb2o_4 _10928_ (.A1_N(_04011_),
    .A2_N(_04012_),
    .B1(net243),
    .B2(_04010_),
    .X(dest_val[12]));
 sky130_fd_sc_hd__a21o_1 _10929_ (.A1(_03896_),
    .A2(_03977_),
    .B1(net157),
    .X(_04013_));
 sky130_fd_sc_hd__o22a_1 _10930_ (.A1(net99),
    .A2(net22),
    .B1(net15),
    .B2(net84),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_1 _10931_ (.A(net69),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__a22o_1 _10932_ (.A1(_06522_),
    .A2(net38),
    .B1(net36),
    .B2(_00148_),
    .X(_04016_));
 sky130_fd_sc_hd__xor2_1 _10933_ (.A(net90),
    .B(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__nand2b_1 _10934_ (.A_N(_04015_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__xor2_1 _10935_ (.A(_04015_),
    .B(_04017_),
    .X(_04019_));
 sky130_fd_sc_hd__a22o_1 _10936_ (.A1(_00157_),
    .A2(net42),
    .B1(net40),
    .B2(net102),
    .X(_04020_));
 sky130_fd_sc_hd__xor2_1 _10937_ (.A(net94),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2b_1 _10938_ (.A_N(_04019_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__xnor2_1 _10939_ (.A(_04019_),
    .B(_04021_),
    .Y(_04023_));
 sky130_fd_sc_hd__o22a_1 _10940_ (.A1(net33),
    .A2(net16),
    .B1(net13),
    .B2(net35),
    .X(_04024_));
 sky130_fd_sc_hd__xnor2_2 _10941_ (.A(net126),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_2 _10942_ (.A(_00324_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__o22a_1 _10943_ (.A1(net74),
    .A2(net12),
    .B1(net6),
    .B2(_00346_),
    .X(_04027_));
 sky130_fd_sc_hd__xor2_2 _10944_ (.A(net122),
    .B(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__and2_1 _10945_ (.A(_04026_),
    .B(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__xor2_2 _10946_ (.A(_04026_),
    .B(_04028_),
    .X(_04030_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(_04023_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__or2_1 _10948_ (.A(_04023_),
    .B(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__o22a_1 _10949_ (.A1(net56),
    .A2(net46),
    .B1(net44),
    .B2(net63),
    .X(_04033_));
 sky130_fd_sc_hd__xnor2_1 _10950_ (.A(net96),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__o22a_1 _10951_ (.A1(net54),
    .A2(net27),
    .B1(net25),
    .B2(net66),
    .X(_04035_));
 sky130_fd_sc_hd__xnor2_1 _10952_ (.A(_00286_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__and2_1 _10953_ (.A(_04034_),
    .B(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_1 _10954_ (.A(_04034_),
    .B(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__nor2_1 _10955_ (.A(_04037_),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__a22o_1 _10956_ (.A1(_06500_),
    .A2(net31),
    .B1(net29),
    .B2(_06534_),
    .X(_04040_));
 sky130_fd_sc_hd__xnor2_1 _10957_ (.A(net49),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__xor2_1 _10958_ (.A(_04039_),
    .B(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__and3_1 _10959_ (.A(_04031_),
    .B(_04032_),
    .C(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__a21oi_1 _10960_ (.A1(_04031_),
    .A2(_04032_),
    .B1(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__o22a_1 _10961_ (.A1(net80),
    .A2(net9),
    .B1(net4),
    .B2(net76),
    .X(_04045_));
 sky130_fd_sc_hd__xnor2_1 _10962_ (.A(net20),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(_03906_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__and2_1 _10964_ (.A(_03906_),
    .B(_04046_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_1 _10965_ (.A(_04047_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nor2_1 _10966_ (.A(net72),
    .B(net19),
    .Y(_04050_));
 sky130_fd_sc_hd__xnor2_1 _10967_ (.A(_04049_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__or3_1 _10968_ (.A(_04043_),
    .B(_04044_),
    .C(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__o21ai_1 _10969_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04051_),
    .Y(_04053_));
 sky130_fd_sc_hd__a21o_1 _10970_ (.A1(_03918_),
    .A2(_03920_),
    .B1(_03916_),
    .X(_04054_));
 sky130_fd_sc_hd__a21oi_1 _10971_ (.A1(_03926_),
    .A2(_03930_),
    .B1(_03936_),
    .Y(_04055_));
 sky130_fd_sc_hd__and3_1 _10972_ (.A(_03926_),
    .B(_03930_),
    .C(_03936_),
    .X(_04056_));
 sky130_fd_sc_hd__or2_1 _10973_ (.A(_04055_),
    .B(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__and2b_1 _10974_ (.A_N(_04057_),
    .B(_04054_),
    .X(_04058_));
 sky130_fd_sc_hd__xnor2_1 _10975_ (.A(_04054_),
    .B(_04057_),
    .Y(_04059_));
 sky130_fd_sc_hd__and3_1 _10976_ (.A(_04052_),
    .B(_04053_),
    .C(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__a21oi_1 _10977_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04059_),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _10978_ (.A(_04060_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__o21ai_1 _10979_ (.A1(_03942_),
    .A2(_03948_),
    .B1(_03950_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21o_1 _10980_ (.A1(_03954_),
    .A2(_03958_),
    .B1(_03957_),
    .X(_04064_));
 sky130_fd_sc_hd__a21bo_1 _10981_ (.A1(_03900_),
    .A2(_03908_),
    .B1_N(_03910_),
    .X(_04065_));
 sky130_fd_sc_hd__nand2_1 _10982_ (.A(_03938_),
    .B(_03940_),
    .Y(_04066_));
 sky130_fd_sc_hd__o31a_1 _10983_ (.A1(net120),
    .A2(net19),
    .A3(_03943_),
    .B1(_03946_),
    .X(_04067_));
 sky130_fd_sc_hd__a21o_1 _10984_ (.A1(_03938_),
    .A2(_03940_),
    .B1(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__xor2_1 _10985_ (.A(_04066_),
    .B(_04067_),
    .X(_04069_));
 sky130_fd_sc_hd__nand2b_1 _10986_ (.A_N(_04069_),
    .B(_04065_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _10987_ (.A(_04065_),
    .B(_04069_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_04064_),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__xor2_1 _10989_ (.A(_04064_),
    .B(_04071_),
    .X(_04073_));
 sky130_fd_sc_hd__xor2_1 _10990_ (.A(_04063_),
    .B(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__nand2_1 _10991_ (.A(_04062_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__or2_1 _10992_ (.A(_04062_),
    .B(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_04075_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__o21a_1 _10994_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_03962_),
    .X(_04078_));
 sky130_fd_sc_hd__or2_1 _10995_ (.A(_04077_),
    .B(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__xnor2_1 _10996_ (.A(_04077_),
    .B(_04078_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21oi_2 _10997_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__and3_1 _10998_ (.A(_03964_),
    .B(_03966_),
    .C(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__or2_2 _10999_ (.A(_04081_),
    .B(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__a21oi_1 _11000_ (.A1(_03849_),
    .A2(_03969_),
    .B1(_03970_),
    .Y(_04084_));
 sky130_fd_sc_hd__nor2_1 _11001_ (.A(_03851_),
    .B(_03971_),
    .Y(_04085_));
 sky130_fd_sc_hd__a21o_1 _11002_ (.A1(_03852_),
    .A2(_04085_),
    .B1(_04084_),
    .X(_04086_));
 sky130_fd_sc_hd__and2_1 _11003_ (.A(_03853_),
    .B(_04085_),
    .X(_04087_));
 sky130_fd_sc_hd__inv_2 _11004_ (.A(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__a21oi_1 _11005_ (.A1(_03621_),
    .A2(_04087_),
    .B1(_04086_),
    .Y(_04089_));
 sky130_fd_sc_hd__o31a_2 _11006_ (.A1(_03091_),
    .A2(_03622_),
    .A3(_04088_),
    .B1(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__xnor2_4 _11007_ (.A(_04083_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21oi_1 _11008_ (.A1(_04013_),
    .A2(_04091_),
    .B1(net187),
    .Y(_04092_));
 sky130_fd_sc_hd__o21a_1 _11009_ (.A1(_04013_),
    .A2(_04091_),
    .B1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__o21ai_1 _11010_ (.A1(net157),
    .A2(_01832_),
    .B1(_01833_),
    .Y(_04094_));
 sky130_fd_sc_hd__or3_1 _11011_ (.A(net157),
    .B(_01832_),
    .C(_01833_),
    .X(_04095_));
 sky130_fd_sc_hd__a21o_1 _11012_ (.A1(_06100_),
    .A2(_03982_),
    .B1(_06088_),
    .X(_04096_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(_06367_),
    .A1(_04096_),
    .S(net285),
    .X(_04097_));
 sky130_fd_sc_hd__nand2_1 _11014_ (.A(_06059_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__o211a_1 _11015_ (.A1(_06059_),
    .A2(_04097_),
    .B1(_04098_),
    .C1(_02323_),
    .X(_04099_));
 sky130_fd_sc_hd__nand2_1 _11016_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .Y(_04100_));
 sky130_fd_sc_hd__or2_1 _11017_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .X(_04101_));
 sky130_fd_sc_hd__nand2_1 _11018_ (.A(_04100_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__a21o_1 _11019_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_03993_),
    .X(_04103_));
 sky130_fd_sc_hd__xnor2_1 _11020_ (.A(_04102_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(_03104_),
    .A1(_03106_),
    .S(net218),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(_02652_),
    .A1(_04105_),
    .S(_06318_),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(_04104_),
    .A1(_04106_),
    .S(net223),
    .X(_04107_));
 sky130_fd_sc_hd__or2_1 _11024_ (.A(\div_res[12] ),
    .B(_03997_),
    .X(_04108_));
 sky130_fd_sc_hd__a21oi_1 _11025_ (.A1(net165),
    .A2(_04108_),
    .B1(\div_res[13] ),
    .Y(_04109_));
 sky130_fd_sc_hd__a311o_1 _11026_ (.A1(\div_res[13] ),
    .A2(net165),
    .A3(_04108_),
    .B1(_04109_),
    .C1(net183),
    .X(_04110_));
 sky130_fd_sc_hd__or2_1 _11027_ (.A(\div_shifter[44] ),
    .B(_04000_),
    .X(_04111_));
 sky130_fd_sc_hd__a21oi_1 _11028_ (.A1(net228),
    .A2(_04111_),
    .B1(\div_shifter[45] ),
    .Y(_04112_));
 sky130_fd_sc_hd__a311o_1 _11029_ (.A1(\div_shifter[45] ),
    .A2(net228),
    .A3(_04111_),
    .B1(_04112_),
    .C1(net231),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(net234),
    .A1(net185),
    .S(_06037_),
    .X(_04114_));
 sky130_fd_sc_hd__a21oi_1 _11031_ (.A1(net186),
    .A2(_04114_),
    .B1(_06048_),
    .Y(_04115_));
 sky130_fd_sc_hd__a21oi_1 _11032_ (.A1(_06026_),
    .A2(net242),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand3_1 _11033_ (.A(_04110_),
    .B(_04113_),
    .C(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__o21a_1 _11034_ (.A1(net220),
    .A2(_02668_),
    .B1(_02342_),
    .X(_04118_));
 sky130_fd_sc_hd__a221o_1 _11035_ (.A1(_02319_),
    .A2(_04106_),
    .B1(_04118_),
    .B2(net170),
    .C1(_04117_),
    .X(_04119_));
 sky130_fd_sc_hd__a211o_1 _11036_ (.A1(net197),
    .A2(_04107_),
    .B1(_04119_),
    .C1(_04099_),
    .X(_04120_));
 sky130_fd_sc_hd__a311o_1 _11037_ (.A1(net233),
    .A2(_04094_),
    .A3(_04095_),
    .B1(_04120_),
    .C1(_04093_),
    .X(_04121_));
 sky130_fd_sc_hd__or2_1 _11038_ (.A(curr_PC[13]),
    .B(_04011_),
    .X(_04122_));
 sky130_fd_sc_hd__a21oi_1 _11039_ (.A1(curr_PC[13]),
    .A2(_04011_),
    .B1(net243),
    .Y(_04123_));
 sky130_fd_sc_hd__a22o_4 _11040_ (.A1(net244),
    .A2(_04121_),
    .B1(_04122_),
    .B2(_04123_),
    .X(dest_val[13]));
 sky130_fd_sc_hd__nand3_2 _11041_ (.A(_03895_),
    .B(_03977_),
    .C(_04091_),
    .Y(_04124_));
 sky130_fd_sc_hd__or2_1 _11042_ (.A(_03657_),
    .B(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__a21bo_1 _11043_ (.A1(_04063_),
    .A2(_04073_),
    .B1_N(_04072_),
    .X(_04126_));
 sky130_fd_sc_hd__a21o_1 _11044_ (.A1(_04039_),
    .A2(_04041_),
    .B1(_04037_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_1 _11045_ (.A(_04018_),
    .B(_04022_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21oi_2 _11046_ (.A1(net137),
    .A2(_04025_),
    .B1(_04029_),
    .Y(_04129_));
 sky130_fd_sc_hd__a21o_1 _11047_ (.A1(_04018_),
    .A2(_04022_),
    .B1(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__xor2_1 _11048_ (.A(_04128_),
    .B(_04129_),
    .X(_04131_));
 sky130_fd_sc_hd__nand2b_1 _11049_ (.A_N(_04131_),
    .B(_04127_),
    .Y(_04132_));
 sky130_fd_sc_hd__xnor2_1 _11050_ (.A(_04127_),
    .B(_04131_),
    .Y(_04133_));
 sky130_fd_sc_hd__o22a_1 _11051_ (.A1(net59),
    .A2(net46),
    .B1(net45),
    .B2(net57),
    .X(_04134_));
 sky130_fd_sc_hd__xnor2_1 _11052_ (.A(net96),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__o22a_1 _11053_ (.A1(net55),
    .A2(net25),
    .B1(net16),
    .B2(net27),
    .X(_04136_));
 sky130_fd_sc_hd__xnor2_1 _11054_ (.A(_00286_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_04135_),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__or2_1 _11056_ (.A(_04135_),
    .B(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__and2_1 _11057_ (.A(_04138_),
    .B(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__a22o_1 _11058_ (.A1(_06492_),
    .A2(net31),
    .B1(net29),
    .B2(_06500_),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_1 _11059_ (.A(net49),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__xor2_1 _11060_ (.A(_04140_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__a22o_1 _11061_ (.A1(_06515_),
    .A2(net38),
    .B1(net36),
    .B2(_06522_),
    .X(_04144_));
 sky130_fd_sc_hd__xor2_1 _11062_ (.A(net89),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__a22o_1 _11063_ (.A1(_00148_),
    .A2(net42),
    .B1(net41),
    .B2(_00157_),
    .X(_04146_));
 sky130_fd_sc_hd__xor2_1 _11064_ (.A(net92),
    .B(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__nand2_1 _11065_ (.A(_04145_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__or2_1 _11066_ (.A(_04145_),
    .B(_04147_),
    .X(_04149_));
 sky130_fd_sc_hd__and2_1 _11067_ (.A(_04148_),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__o22a_1 _11068_ (.A1(net33),
    .A2(net13),
    .B1(net12),
    .B2(net35),
    .X(_04151_));
 sky130_fd_sc_hd__xnor2_1 _11069_ (.A(net126),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__or2_1 _11070_ (.A(_00345_),
    .B(net6),
    .X(_04153_));
 sky130_fd_sc_hd__nor2_1 _11071_ (.A(_00344_),
    .B(net6),
    .Y(_04154_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(_04153_),
    .A1(_04154_),
    .S(net122),
    .X(_04155_));
 sky130_fd_sc_hd__nor2_1 _11073_ (.A(_04152_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__and2_1 _11074_ (.A(_04152_),
    .B(_04155_),
    .X(_04157_));
 sky130_fd_sc_hd__nor2_1 _11075_ (.A(_04156_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__and2b_1 _11076_ (.A_N(_04158_),
    .B(_04150_),
    .X(_04159_));
 sky130_fd_sc_hd__xnor2_1 _11077_ (.A(_04150_),
    .B(_04158_),
    .Y(_04160_));
 sky130_fd_sc_hd__xnor2_1 _11078_ (.A(_04143_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__o22a_1 _11079_ (.A1(net84),
    .A2(net10),
    .B1(net5),
    .B2(net80),
    .X(_04162_));
 sky130_fd_sc_hd__xnor2_1 _11080_ (.A(net19),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__o22a_1 _11081_ (.A1(net101),
    .A2(net22),
    .B1(net14),
    .B2(net99),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_1 _11082_ (.A(net69),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__nor2_1 _11083_ (.A(net76),
    .B(net20),
    .Y(_04166_));
 sky130_fd_sc_hd__xnor2_1 _11084_ (.A(_04165_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand2b_1 _11085_ (.A_N(_04163_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__xor2_1 _11086_ (.A(_04163_),
    .B(_04167_),
    .X(_04169_));
 sky130_fd_sc_hd__nor2_1 _11087_ (.A(_04161_),
    .B(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(_04161_),
    .B(_04169_),
    .Y(_04171_));
 sky130_fd_sc_hd__and2b_1 _11089_ (.A_N(_04170_),
    .B(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__xor2_1 _11090_ (.A(_04133_),
    .B(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__a21bo_1 _11091_ (.A1(_04053_),
    .A2(_04059_),
    .B1_N(_04052_),
    .X(_04174_));
 sky130_fd_sc_hd__or2_1 _11092_ (.A(_04055_),
    .B(_04058_),
    .X(_04175_));
 sky130_fd_sc_hd__a21o_1 _11093_ (.A1(_04023_),
    .A2(_04030_),
    .B1(_04043_),
    .X(_04176_));
 sky130_fd_sc_hd__a21o_1 _11094_ (.A1(_04049_),
    .A2(_04050_),
    .B1(_04047_),
    .X(_04177_));
 sky130_fd_sc_hd__nand2_1 _11095_ (.A(_04176_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__xor2_1 _11096_ (.A(_04176_),
    .B(_04177_),
    .X(_04179_));
 sky130_fd_sc_hd__xnor2_1 _11097_ (.A(_04175_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__and2_1 _11098_ (.A(_04068_),
    .B(_04070_),
    .X(_04181_));
 sky130_fd_sc_hd__xnor2_1 _11099_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2b_1 _11100_ (.A_N(_04182_),
    .B(_04174_),
    .Y(_04183_));
 sky130_fd_sc_hd__xnor2_2 _11101_ (.A(_04174_),
    .B(_04182_),
    .Y(_04184_));
 sky130_fd_sc_hd__nand2_1 _11102_ (.A(_04173_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__xnor2_1 _11103_ (.A(_04173_),
    .B(_04184_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2b_1 _11104_ (.A_N(_04186_),
    .B(_04126_),
    .Y(_04187_));
 sky130_fd_sc_hd__xor2_1 _11105_ (.A(_04126_),
    .B(_04186_),
    .X(_04188_));
 sky130_fd_sc_hd__a21oi_1 _11106_ (.A1(_04075_),
    .A2(_04079_),
    .B1(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__and3_1 _11107_ (.A(_04075_),
    .B(_04079_),
    .C(_04188_),
    .X(_04190_));
 sky130_fd_sc_hd__or2_2 _11108_ (.A(_04189_),
    .B(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__o21ba_1 _11109_ (.A1(_03968_),
    .A2(_04081_),
    .B1_N(_04082_),
    .X(_04192_));
 sky130_fd_sc_hd__nor2_1 _11110_ (.A(_03971_),
    .B(_04083_),
    .Y(_04193_));
 sky130_fd_sc_hd__a21oi_1 _11111_ (.A1(_03972_),
    .A2(_04193_),
    .B1(_04192_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _11112_ (.A(_03973_),
    .B(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__o21ai_4 _11113_ (.A1(_03739_),
    .A2(_04195_),
    .B1(_04194_),
    .Y(_04196_));
 sky130_fd_sc_hd__xnor2_4 _11114_ (.A(_04191_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__and3_1 _11115_ (.A(net165),
    .B(_04125_),
    .C(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__a21oi_1 _11116_ (.A1(net165),
    .A2(_04125_),
    .B1(_04197_),
    .Y(_04199_));
 sky130_fd_sc_hd__a22oi_2 _11117_ (.A1(net159),
    .A2(_01834_),
    .B1(_01836_),
    .B2(_01837_),
    .Y(_04200_));
 sky130_fd_sc_hd__a41o_1 _11118_ (.A1(net159),
    .A2(_01834_),
    .A3(_01836_),
    .A4(_01837_),
    .B1(_02330_),
    .X(_04201_));
 sky130_fd_sc_hd__a21o_1 _11119_ (.A1(_06059_),
    .A2(_04096_),
    .B1(_06037_),
    .X(_04202_));
 sky130_fd_sc_hd__nand2_1 _11120_ (.A(net284),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__o21ai_1 _11121_ (.A1(net284),
    .A2(_06369_),
    .B1(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ai_1 _11122_ (.A1(_05993_),
    .A2(_04204_),
    .B1(_02323_),
    .Y(_04205_));
 sky130_fd_sc_hd__a21o_1 _11123_ (.A1(_05993_),
    .A2(_04204_),
    .B1(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2_1 _11124_ (.A(net291),
    .B(curr_PC[14]),
    .Y(_04207_));
 sky130_fd_sc_hd__or2_1 _11125_ (.A(net291),
    .B(curr_PC[14]),
    .X(_04208_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21bo_1 _11127_ (.A1(_04101_),
    .A2(_04103_),
    .B1_N(_04100_),
    .X(_04210_));
 sky130_fd_sc_hd__xnor2_1 _11128_ (.A(_04209_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__nor2_1 _11129_ (.A(net223),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(_03239_),
    .A1(_03241_),
    .S(net217),
    .X(_04213_));
 sky130_fd_sc_hd__or2_1 _11131_ (.A(net220),
    .B(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__o21ai_2 _11132_ (.A1(_06318_),
    .A2(_02529_),
    .B1(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__a211o_1 _11133_ (.A1(net223),
    .A2(_04215_),
    .B1(_04212_),
    .C1(net196),
    .X(_04216_));
 sky130_fd_sc_hd__or2_1 _11134_ (.A(\div_res[13] ),
    .B(_04108_),
    .X(_04217_));
 sky130_fd_sc_hd__a21oi_1 _11135_ (.A1(net163),
    .A2(_04217_),
    .B1(\div_res[14] ),
    .Y(_04218_));
 sky130_fd_sc_hd__a31o_1 _11136_ (.A1(\div_res[14] ),
    .A2(net163),
    .A3(_04217_),
    .B1(net184),
    .X(_04219_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(net234),
    .A1(net185),
    .S(_05982_),
    .X(_04220_));
 sky130_fd_sc_hd__a2bb2o_1 _11138_ (.A1_N(net291),
    .A2_N(_05965_),
    .B1(net186),
    .B2(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__or2_1 _11139_ (.A(\div_shifter[45] ),
    .B(_04111_),
    .X(_04222_));
 sky130_fd_sc_hd__a21oi_1 _11140_ (.A1(net226),
    .A2(_04222_),
    .B1(\div_shifter[46] ),
    .Y(_04223_));
 sky130_fd_sc_hd__a31o_1 _11141_ (.A1(\div_shifter[46] ),
    .A2(net226),
    .A3(_04222_),
    .B1(net232),
    .X(_04224_));
 sky130_fd_sc_hd__o22a_1 _11142_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04223_),
    .B2(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__o21ai_2 _11143_ (.A1(net220),
    .A2(_02502_),
    .B1(_02342_),
    .Y(_04226_));
 sky130_fd_sc_hd__o211a_1 _11144_ (.A1(net168),
    .A2(_04226_),
    .B1(_04225_),
    .C1(_04221_),
    .X(_04227_));
 sky130_fd_sc_hd__o211a_1 _11145_ (.A1(_02320_),
    .A2(_04215_),
    .B1(_04216_),
    .C1(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__o211a_1 _11146_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04206_),
    .C1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__o31a_1 _11147_ (.A1(net187),
    .A2(_04198_),
    .A3(_04199_),
    .B1(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__o2bb2a_1 _11148_ (.A1_N(_05965_),
    .A2_N(net242),
    .B1(_06463_),
    .B2(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__and3_1 _11149_ (.A(curr_PC[13]),
    .B(curr_PC[14]),
    .C(_04011_),
    .X(_04232_));
 sky130_fd_sc_hd__a21oi_1 _11150_ (.A1(curr_PC[13]),
    .A2(_04011_),
    .B1(curr_PC[14]),
    .Y(_04233_));
 sky130_fd_sc_hd__or3_2 _11151_ (.A(net244),
    .B(_04232_),
    .C(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__o21ai_4 _11152_ (.A1(net248),
    .A2(_04231_),
    .B1(_04234_),
    .Y(dest_val[14]));
 sky130_fd_sc_hd__o21a_1 _11153_ (.A1(_04125_),
    .A2(_04197_),
    .B1(net165),
    .X(_04235_));
 sky130_fd_sc_hd__o22a_1 _11154_ (.A1(net99),
    .A2(net10),
    .B1(net5),
    .B2(net84),
    .X(_04236_));
 sky130_fd_sc_hd__xnor2_1 _11155_ (.A(net20),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__a22o_1 _11156_ (.A1(_06522_),
    .A2(net43),
    .B1(net41),
    .B2(_00148_),
    .X(_04238_));
 sky130_fd_sc_hd__xor2_1 _11157_ (.A(net93),
    .B(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__nand2b_1 _11158_ (.A_N(_04237_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2b_1 _11159_ (.A_N(_04239_),
    .B(_04237_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_1 _11160_ (.A(_04240_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__o22a_1 _11161_ (.A1(net51),
    .A2(net23),
    .B1(net15),
    .B2(net101),
    .X(_04243_));
 sky130_fd_sc_hd__xnor2_1 _11162_ (.A(net68),
    .B(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__or2_1 _11163_ (.A(_04242_),
    .B(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__nand2_1 _11164_ (.A(_04242_),
    .B(_04244_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _11165_ (.A(_04245_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__o22a_1 _11166_ (.A1(net25),
    .A2(net16),
    .B1(net13),
    .B2(net27),
    .X(_04248_));
 sky130_fd_sc_hd__xnor2_1 _11167_ (.A(net88),
    .B(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__and2_1 _11168_ (.A(net121),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nor2_1 _11169_ (.A(net122),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__nor2_1 _11170_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o22a_1 _11171_ (.A1(net33),
    .A2(net12),
    .B1(net6),
    .B2(net35),
    .X(_04253_));
 sky130_fd_sc_hd__xnor2_2 _11172_ (.A(net126),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__xor2_2 _11173_ (.A(_04252_),
    .B(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__a22o_1 _11174_ (.A1(_06538_),
    .A2(net38),
    .B1(net36),
    .B2(_06515_),
    .X(_04256_));
 sky130_fd_sc_hd__xor2_1 _11175_ (.A(net89),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__a22o_1 _11176_ (.A1(_06553_),
    .A2(net31),
    .B1(net29),
    .B2(_06492_),
    .X(_04258_));
 sky130_fd_sc_hd__xnor2_1 _11177_ (.A(net49),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__and2_1 _11178_ (.A(_04257_),
    .B(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__nor2_1 _11179_ (.A(_04257_),
    .B(_04259_),
    .Y(_04261_));
 sky130_fd_sc_hd__nor2_1 _11180_ (.A(_04260_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__o22a_1 _11181_ (.A1(net65),
    .A2(net46),
    .B1(net44),
    .B2(net59),
    .X(_04263_));
 sky130_fd_sc_hd__xnor2_2 _11182_ (.A(net95),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__xor2_2 _11183_ (.A(_04262_),
    .B(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__xnor2_2 _11184_ (.A(_04148_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__xnor2_2 _11185_ (.A(_04255_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__xnor2_1 _11186_ (.A(_04247_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21bo_1 _11187_ (.A1(_04140_),
    .A2(_04142_),
    .B1_N(_04138_),
    .X(_04269_));
 sky130_fd_sc_hd__nor2_1 _11188_ (.A(net80),
    .B(net19),
    .Y(_04270_));
 sky130_fd_sc_hd__xnor2_1 _11189_ (.A(_04269_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__or2_1 _11190_ (.A(_04156_),
    .B(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__nand2_1 _11191_ (.A(_04156_),
    .B(_04271_),
    .Y(_04273_));
 sky130_fd_sc_hd__and2_1 _11192_ (.A(_04272_),
    .B(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2b_1 _11193_ (.A_N(_04268_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_2 _11194_ (.A(_04268_),
    .B(_04274_),
    .Y(_04276_));
 sky130_fd_sc_hd__a21o_1 _11195_ (.A1(_04133_),
    .A2(_04171_),
    .B1(_04170_),
    .X(_04277_));
 sky130_fd_sc_hd__a21bo_1 _11196_ (.A1(_04175_),
    .A2(_04179_),
    .B1_N(_04178_),
    .X(_04278_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(_04130_),
    .B(_04132_),
    .Y(_04279_));
 sky130_fd_sc_hd__a21o_1 _11198_ (.A1(_04143_),
    .A2(_04160_),
    .B1(_04159_),
    .X(_04280_));
 sky130_fd_sc_hd__o31a_1 _11199_ (.A1(net76),
    .A2(net20),
    .A3(_04165_),
    .B1(_04168_),
    .X(_04281_));
 sky130_fd_sc_hd__inv_2 _11200_ (.A(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__and2_1 _11201_ (.A(_04280_),
    .B(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__xnor2_2 _11202_ (.A(_04280_),
    .B(_04282_),
    .Y(_04284_));
 sky130_fd_sc_hd__inv_2 _11203_ (.A(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__xnor2_2 _11204_ (.A(_04279_),
    .B(_04284_),
    .Y(_04286_));
 sky130_fd_sc_hd__xnor2_2 _11205_ (.A(_04278_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand2b_1 _11206_ (.A_N(_04287_),
    .B(_04277_),
    .Y(_04288_));
 sky130_fd_sc_hd__xnor2_2 _11207_ (.A(_04277_),
    .B(_04287_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(_04276_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_2 _11209_ (.A(_04276_),
    .B(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__o21ai_2 _11210_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04183_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand2b_1 _11211_ (.A_N(_04291_),
    .B(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__xor2_2 _11212_ (.A(_04291_),
    .B(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__a21oi_2 _11213_ (.A1(_04185_),
    .A2(_04187_),
    .B1(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand3_1 _11214_ (.A(_04185_),
    .B(_04187_),
    .C(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__nand2b_2 _11215_ (.A_N(_04295_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__o21ba_1 _11216_ (.A1(_04081_),
    .A2(_04189_),
    .B1_N(_04190_),
    .X(_04298_));
 sky130_fd_sc_hd__nor2_1 _11217_ (.A(_04083_),
    .B(_04191_),
    .Y(_04299_));
 sky130_fd_sc_hd__a21o_1 _11218_ (.A1(_04084_),
    .A2(_04299_),
    .B1(_04298_),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_1 _11219_ (.A(_04085_),
    .B(_04299_),
    .Y(_04301_));
 sky130_fd_sc_hd__o21ba_1 _11220_ (.A1(_03857_),
    .A2(_04301_),
    .B1_N(_04300_),
    .X(_04302_));
 sky130_fd_sc_hd__xor2_4 _11221_ (.A(_04297_),
    .B(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__a21oi_1 _11222_ (.A1(_04235_),
    .A2(_04303_),
    .B1(net187),
    .Y(_04304_));
 sky130_fd_sc_hd__o21a_1 _11223_ (.A1(_04235_),
    .A2(_04303_),
    .B1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__a21oi_1 _11224_ (.A1(net159),
    .A2(_01838_),
    .B1(_01840_),
    .Y(_04306_));
 sky130_fd_sc_hd__a311oi_4 _11225_ (.A1(net159),
    .A2(_01838_),
    .A3(_01840_),
    .B1(_02330_),
    .C1(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21o_1 _11226_ (.A1(_05993_),
    .A2(_04202_),
    .B1(_05982_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(_06371_),
    .A1(_04308_),
    .S(net284),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_05953_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__o211a_1 _11229_ (.A1(_05953_),
    .A2(_04309_),
    .B1(_04310_),
    .C1(_02323_),
    .X(_04311_));
 sky130_fd_sc_hd__and2_1 _11230_ (.A(net290),
    .B(curr_PC[15]),
    .X(_04312_));
 sky130_fd_sc_hd__or2_1 _11231_ (.A(net290),
    .B(curr_PC[15]),
    .X(_04313_));
 sky130_fd_sc_hd__and2b_1 _11232_ (.A_N(_04312_),
    .B(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__a21bo_1 _11233_ (.A1(_04208_),
    .A2(_04210_),
    .B1_N(_04207_),
    .X(_04315_));
 sky130_fd_sc_hd__xnor2_1 _11234_ (.A(_04314_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(_03374_),
    .A1(_03376_),
    .S(net217),
    .X(_04317_));
 sky130_fd_sc_hd__inv_2 _11236_ (.A(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(_02348_),
    .A1(_04318_),
    .S(_06318_),
    .X(_04319_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(_04316_),
    .A1(_04319_),
    .S(net224),
    .X(_04320_));
 sky130_fd_sc_hd__or2_1 _11239_ (.A(\div_res[14] ),
    .B(_04217_),
    .X(_04321_));
 sky130_fd_sc_hd__and3_1 _11240_ (.A(\div_res[15] ),
    .B(net163),
    .C(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__a21oi_1 _11241_ (.A1(net163),
    .A2(_04321_),
    .B1(\div_res[15] ),
    .Y(_04323_));
 sky130_fd_sc_hd__or3_1 _11242_ (.A(net184),
    .B(_04322_),
    .C(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__or3_1 _11243_ (.A(\div_shifter[46] ),
    .B(\div_shifter[45] ),
    .C(_04111_),
    .X(_04325_));
 sky130_fd_sc_hd__a21oi_1 _11244_ (.A1(net226),
    .A2(_04325_),
    .B1(\div_shifter[47] ),
    .Y(_04326_));
 sky130_fd_sc_hd__a311o_1 _11245_ (.A1(\div_shifter[47] ),
    .A2(net226),
    .A3(_04325_),
    .B1(_04326_),
    .C1(net231),
    .X(_04327_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(net234),
    .A1(net185),
    .S(_05941_),
    .X(_04328_));
 sky130_fd_sc_hd__a21oi_1 _11247_ (.A1(net186),
    .A2(_04328_),
    .B1(_05947_),
    .Y(_04329_));
 sky130_fd_sc_hd__a21oi_1 _11248_ (.A1(_05935_),
    .A2(net242),
    .B1(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__and3_1 _11249_ (.A(_04324_),
    .B(_04327_),
    .C(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__o21a_1 _11250_ (.A1(net220),
    .A2(_02312_),
    .B1(_02342_),
    .X(_04332_));
 sky130_fd_sc_hd__o2bb2a_1 _11251_ (.A1_N(net170),
    .A2_N(_04332_),
    .B1(_04319_),
    .B2(_02320_),
    .X(_04333_));
 sky130_fd_sc_hd__o211a_1 _11252_ (.A1(net196),
    .A2(_04320_),
    .B1(_04331_),
    .C1(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__or4b_2 _11253_ (.A(_04305_),
    .B(_04307_),
    .C(_04311_),
    .D_N(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__or2_1 _11254_ (.A(curr_PC[15]),
    .B(_04232_),
    .X(_04336_));
 sky130_fd_sc_hd__and2_1 _11255_ (.A(curr_PC[15]),
    .B(_04232_),
    .X(_04337_));
 sky130_fd_sc_hd__nor2_1 _11256_ (.A(net243),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a22o_4 _11257_ (.A1(net243),
    .A2(_04335_),
    .B1(_04336_),
    .B2(_04338_),
    .X(dest_val[15]));
 sky130_fd_sc_hd__or2_1 _11258_ (.A(_04197_),
    .B(_04303_),
    .X(_04339_));
 sky130_fd_sc_hd__or2_1 _11259_ (.A(_04125_),
    .B(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__a21oi_1 _11260_ (.A1(_04262_),
    .A2(_04264_),
    .B1(_04260_),
    .Y(_04341_));
 sky130_fd_sc_hd__o22a_1 _11261_ (.A1(net66),
    .A2(net46),
    .B1(net44),
    .B2(net65),
    .X(_04342_));
 sky130_fd_sc_hd__xnor2_1 _11262_ (.A(net95),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__a22oi_1 _11263_ (.A1(_06553_),
    .A2(net29),
    .B1(_00398_),
    .B2(net31),
    .Y(_04344_));
 sky130_fd_sc_hd__xnor2_1 _11264_ (.A(_00201_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_04343_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__or2_1 _11266_ (.A(_04343_),
    .B(_04345_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _11267_ (.A(_04346_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_1 _11268_ (.A(_04341_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__xnor2_1 _11269_ (.A(_04341_),
    .B(_04348_),
    .Y(_04351_));
 sky130_fd_sc_hd__o22a_1 _11270_ (.A1(net25),
    .A2(net13),
    .B1(net11),
    .B2(net27),
    .X(_04352_));
 sky130_fd_sc_hd__xnor2_1 _11271_ (.A(net88),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__o21ai_2 _11272_ (.A1(_00267_),
    .A2(net7),
    .B1(net125),
    .Y(_04354_));
 sky130_fd_sc_hd__o21ai_4 _11273_ (.A1(_00277_),
    .A2(net7),
    .B1(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__nor2_1 _11274_ (.A(_04353_),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__and2_1 _11275_ (.A(_04353_),
    .B(_04355_),
    .X(_04357_));
 sky130_fd_sc_hd__nor2_1 _11276_ (.A(_04356_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(_04351_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__and2_1 _11278_ (.A(_04351_),
    .B(_04358_),
    .X(_04360_));
 sky130_fd_sc_hd__or2_1 _11279_ (.A(_04359_),
    .B(_04360_),
    .X(_04362_));
 sky130_fd_sc_hd__o22a_1 _11280_ (.A1(net53),
    .A2(net22),
    .B1(net14),
    .B2(net51),
    .X(_04363_));
 sky130_fd_sc_hd__xnor2_1 _11281_ (.A(net68),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__inv_2 _11282_ (.A(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__a22o_1 _11283_ (.A1(_06534_),
    .A2(net38),
    .B1(net36),
    .B2(_06538_),
    .X(_04366_));
 sky130_fd_sc_hd__xor2_1 _11284_ (.A(net89),
    .B(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__xor2_1 _11285_ (.A(_04364_),
    .B(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__a22o_1 _11286_ (.A1(_06515_),
    .A2(net42),
    .B1(net40),
    .B2(_06522_),
    .X(_04369_));
 sky130_fd_sc_hd__xor2_1 _11287_ (.A(net92),
    .B(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__and2b_1 _11288_ (.A_N(_04368_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__and2b_1 _11289_ (.A_N(_04370_),
    .B(_04368_),
    .X(_04373_));
 sky130_fd_sc_hd__or2_1 _11290_ (.A(_04371_),
    .B(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__xnor2_2 _11291_ (.A(_04362_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__a21oi_2 _11292_ (.A1(_04252_),
    .A2(_04254_),
    .B1(_04250_),
    .Y(_04376_));
 sky130_fd_sc_hd__o22a_1 _11293_ (.A1(net101),
    .A2(net9),
    .B1(net4),
    .B2(net99),
    .X(_04377_));
 sky130_fd_sc_hd__xnor2_2 _11294_ (.A(net18),
    .B(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__xnor2_1 _11295_ (.A(_04376_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__or3_1 _11296_ (.A(net84),
    .B(net19),
    .C(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__o21ai_1 _11297_ (.A1(net84),
    .A2(net19),
    .B1(_04379_),
    .Y(_04381_));
 sky130_fd_sc_hd__and2_1 _11298_ (.A(_04380_),
    .B(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__and2b_1 _11299_ (.A_N(_04375_),
    .B(_04382_),
    .X(_04384_));
 sky130_fd_sc_hd__xnor2_2 _11300_ (.A(_04375_),
    .B(_04382_),
    .Y(_04385_));
 sky130_fd_sc_hd__o21ai_2 _11301_ (.A1(_04247_),
    .A2(_04267_),
    .B1(_04275_),
    .Y(_04386_));
 sky130_fd_sc_hd__a21bo_1 _11302_ (.A1(_04269_),
    .A2(_04270_),
    .B1_N(_04272_),
    .X(_04387_));
 sky130_fd_sc_hd__a32oi_2 _11303_ (.A1(_04145_),
    .A2(_04147_),
    .A3(_04265_),
    .B1(_04266_),
    .B2(_04255_),
    .Y(_04388_));
 sky130_fd_sc_hd__a21oi_1 _11304_ (.A1(_04240_),
    .A2(_04245_),
    .B1(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__and3_1 _11305_ (.A(_04240_),
    .B(_04245_),
    .C(_04388_),
    .X(_04390_));
 sky130_fd_sc_hd__nor2_1 _11306_ (.A(_04389_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__xnor2_2 _11307_ (.A(_04387_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__a21oi_2 _11308_ (.A1(_04279_),
    .A2(_04285_),
    .B1(_04283_),
    .Y(_04393_));
 sky130_fd_sc_hd__xnor2_2 _11309_ (.A(_04392_),
    .B(_04393_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2b_1 _11310_ (.A_N(_04395_),
    .B(_04386_),
    .Y(_04396_));
 sky130_fd_sc_hd__xnor2_2 _11311_ (.A(_04386_),
    .B(_04395_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _11312_ (.A(_04385_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__xnor2_2 _11313_ (.A(_04385_),
    .B(_04397_),
    .Y(_04399_));
 sky130_fd_sc_hd__a21boi_2 _11314_ (.A1(_04278_),
    .A2(_04286_),
    .B1_N(_04288_),
    .Y(_04400_));
 sky130_fd_sc_hd__or2_1 _11315_ (.A(_04399_),
    .B(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__xnor2_2 _11316_ (.A(_04399_),
    .B(_04400_),
    .Y(_04402_));
 sky130_fd_sc_hd__a21oi_2 _11317_ (.A1(_04290_),
    .A2(_04293_),
    .B1(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand3_2 _11318_ (.A(_04290_),
    .B(_04293_),
    .C(_04402_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2b_2 _11319_ (.A_N(_04403_),
    .B(_04404_),
    .Y(_04406_));
 sky130_fd_sc_hd__o21a_1 _11320_ (.A1(_04189_),
    .A2(_04295_),
    .B1(_04296_),
    .X(_04407_));
 sky130_fd_sc_hd__nor2_1 _11321_ (.A(_04191_),
    .B(_04297_),
    .Y(_04408_));
 sky130_fd_sc_hd__and2_1 _11322_ (.A(_04193_),
    .B(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__a221o_1 _11323_ (.A1(_04192_),
    .A2(_04408_),
    .B1(_04409_),
    .B2(_03974_),
    .C1(_04407_),
    .X(_04410_));
 sky130_fd_sc_hd__a31o_2 _11324_ (.A1(_03410_),
    .A2(_03975_),
    .A3(_04409_),
    .B1(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__xnor2_4 _11325_ (.A(_04406_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__a21oi_1 _11326_ (.A1(net165),
    .A2(_04340_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a31o_1 _11327_ (.A1(net165),
    .A2(_04340_),
    .A3(_04412_),
    .B1(net187),
    .X(_04414_));
 sky130_fd_sc_hd__a21oi_1 _11328_ (.A1(net159),
    .A2(_01841_),
    .B1(_01846_),
    .Y(_04415_));
 sky130_fd_sc_hd__a31o_1 _11329_ (.A1(net159),
    .A2(_01841_),
    .A3(_01846_),
    .B1(_02330_),
    .X(_04417_));
 sky130_fd_sc_hd__a21o_1 _11330_ (.A1(_05953_),
    .A2(_04308_),
    .B1(_05941_),
    .X(_04418_));
 sky130_fd_sc_hd__nand2_1 _11331_ (.A(net284),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__o21a_1 _11332_ (.A1(net284),
    .A2(_06373_),
    .B1(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__xnor2_1 _11333_ (.A(_05919_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__a21oi_1 _11334_ (.A1(_04313_),
    .A2(_04315_),
    .B1(_04312_),
    .Y(_04422_));
 sky130_fd_sc_hd__nor2_1 _11335_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04423_));
 sky130_fd_sc_hd__nand2_1 _11336_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2b_1 _11337_ (.A_N(_04423_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__xnor2_1 _11338_ (.A(_04422_),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(net250),
    .B(_04332_),
    .Y(_04428_));
 sky130_fd_sc_hd__a211o_1 _11340_ (.A1(net250),
    .A2(_04426_),
    .B1(_04428_),
    .C1(_06449_),
    .X(_04429_));
 sky130_fd_sc_hd__or2_1 _11341_ (.A(\div_shifter[47] ),
    .B(_04325_),
    .X(_04430_));
 sky130_fd_sc_hd__a21oi_1 _11342_ (.A1(net226),
    .A2(_04430_),
    .B1(\div_shifter[48] ),
    .Y(_04431_));
 sky130_fd_sc_hd__a311o_1 _11343_ (.A1(\div_shifter[48] ),
    .A2(net226),
    .A3(_04430_),
    .B1(_04431_),
    .C1(net231),
    .X(_04432_));
 sky130_fd_sc_hd__o21a_1 _11344_ (.A1(_05892_),
    .A2(net234),
    .B1(net186),
    .X(_04433_));
 sky130_fd_sc_hd__o2bb2a_1 _11345_ (.A1_N(_05892_),
    .A2_N(_02331_),
    .B1(net241),
    .B2(_05883_),
    .X(_04434_));
 sky130_fd_sc_hd__o211a_1 _11346_ (.A1(_05901_),
    .A2(_04433_),
    .B1(_04434_),
    .C1(_04432_),
    .X(_04435_));
 sky130_fd_sc_hd__or2_1 _11347_ (.A(\div_res[15] ),
    .B(_04321_),
    .X(_04436_));
 sky130_fd_sc_hd__a21oi_1 _11348_ (.A1(net163),
    .A2(_04436_),
    .B1(\div_res[16] ),
    .Y(_04437_));
 sky130_fd_sc_hd__a31o_1 _11349_ (.A1(\div_res[16] ),
    .A2(net164),
    .A3(_04436_),
    .B1(net183),
    .X(_04439_));
 sky130_fd_sc_hd__o2bb2a_1 _11350_ (.A1_N(_02319_),
    .A2_N(_04332_),
    .B1(_04437_),
    .B2(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__o211a_1 _11351_ (.A1(net168),
    .A2(_04319_),
    .B1(_04435_),
    .C1(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__o211a_1 _11352_ (.A1(net236),
    .A2(_04421_),
    .B1(_04429_),
    .C1(_04441_),
    .X(_04442_));
 sky130_fd_sc_hd__o221a_1 _11353_ (.A1(_04413_),
    .A2(_04414_),
    .B1(_04415_),
    .B2(_04417_),
    .C1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__nand2_1 _11354_ (.A(curr_PC[16]),
    .B(_04337_),
    .Y(_04444_));
 sky130_fd_sc_hd__o21a_1 _11355_ (.A1(curr_PC[16]),
    .A2(_04337_),
    .B1(net248),
    .X(_04445_));
 sky130_fd_sc_hd__a2bb2o_4 _11356_ (.A1_N(net248),
    .A2_N(_04443_),
    .B1(_04444_),
    .B2(_04445_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__o31a_1 _11357_ (.A1(_04125_),
    .A2(_04339_),
    .A3(_04412_),
    .B1(net166),
    .X(_04446_));
 sky130_fd_sc_hd__a22o_1 _11358_ (.A1(net29),
    .A2(_00398_),
    .B1(_00690_),
    .B2(net31),
    .X(_04447_));
 sky130_fd_sc_hd__xnor2_1 _11359_ (.A(net49),
    .B(_04447_),
    .Y(_04449_));
 sky130_fd_sc_hd__and2_1 _11360_ (.A(net124),
    .B(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__xnor2_1 _11361_ (.A(net124),
    .B(_04449_),
    .Y(_04451_));
 sky130_fd_sc_hd__o22a_1 _11362_ (.A1(net25),
    .A2(net11),
    .B1(_02070_),
    .B2(_00308_),
    .X(_04452_));
 sky130_fd_sc_hd__xnor2_1 _11363_ (.A(net88),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__and2b_1 _11364_ (.A_N(_04451_),
    .B(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__xor2_1 _11365_ (.A(_04451_),
    .B(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _11366_ (.A(_04356_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__xor2_1 _11367_ (.A(_04356_),
    .B(_04455_),
    .X(_04457_));
 sky130_fd_sc_hd__nand2b_1 _11368_ (.A_N(_04346_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__xnor2_1 _11369_ (.A(_04346_),
    .B(_04457_),
    .Y(_04460_));
 sky130_fd_sc_hd__a22o_1 _11370_ (.A1(_06538_),
    .A2(net42),
    .B1(net40),
    .B2(_06515_),
    .X(_04461_));
 sky130_fd_sc_hd__xor2_1 _11371_ (.A(net92),
    .B(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__o22a_1 _11372_ (.A1(net54),
    .A2(net46),
    .B1(net44),
    .B2(net66),
    .X(_04463_));
 sky130_fd_sc_hd__xnor2_1 _11373_ (.A(net95),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__and2_1 _11374_ (.A(_04462_),
    .B(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__nor2_1 _11375_ (.A(_04462_),
    .B(_04464_),
    .Y(_04466_));
 sky130_fd_sc_hd__nor2_1 _11376_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a22o_1 _11377_ (.A1(_06500_),
    .A2(net38),
    .B1(net36),
    .B2(_06534_),
    .X(_04468_));
 sky130_fd_sc_hd__xor2_2 _11378_ (.A(net89),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__xor2_1 _11379_ (.A(_04467_),
    .B(_04469_),
    .X(_04471_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(_04460_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__or2_1 _11381_ (.A(_04460_),
    .B(_04471_),
    .X(_04473_));
 sky130_fd_sc_hd__o22a_1 _11382_ (.A1(net51),
    .A2(net9),
    .B1(net4),
    .B2(net101),
    .X(_04474_));
 sky130_fd_sc_hd__xnor2_1 _11383_ (.A(net18),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__o22a_1 _11384_ (.A1(net61),
    .A2(net22),
    .B1(net14),
    .B2(net53),
    .X(_04476_));
 sky130_fd_sc_hd__xnor2_2 _11385_ (.A(net68),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_1 _11386_ (.A(net99),
    .B(net18),
    .Y(_04478_));
 sky130_fd_sc_hd__xnor2_1 _11387_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand2b_1 _11388_ (.A_N(_04475_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__xnor2_1 _11389_ (.A(_04475_),
    .B(_04479_),
    .Y(_04482_));
 sky130_fd_sc_hd__and3_1 _11390_ (.A(_04472_),
    .B(_04473_),
    .C(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__a21oi_1 _11391_ (.A1(_04472_),
    .A2(_04473_),
    .B1(_04482_),
    .Y(_04484_));
 sky130_fd_sc_hd__nor2_1 _11392_ (.A(_04483_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__o21ba_1 _11393_ (.A1(_04362_),
    .A2(_04374_),
    .B1_N(_04384_),
    .X(_04486_));
 sky130_fd_sc_hd__o21ai_2 _11394_ (.A1(_04376_),
    .A2(_04378_),
    .B1(_04380_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_1 _11395_ (.A1(_04365_),
    .A2(_04367_),
    .B1(_04371_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21ba_1 _11396_ (.A1(_04349_),
    .A2(_04359_),
    .B1_N(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__or3b_1 _11397_ (.A(_04349_),
    .B(_04359_),
    .C_N(_04488_),
    .X(_04490_));
 sky130_fd_sc_hd__and2b_1 _11398_ (.A_N(_04489_),
    .B(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__xnor2_1 _11399_ (.A(_04487_),
    .B(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21o_1 _11400_ (.A1(_04387_),
    .A2(_04391_),
    .B1(_04389_),
    .X(_04494_));
 sky130_fd_sc_hd__nand2b_1 _11401_ (.A_N(_04493_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__xnor2_2 _11402_ (.A(_04493_),
    .B(_04494_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand2b_1 _11403_ (.A_N(_04486_),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__xnor2_2 _11404_ (.A(_04486_),
    .B(_04496_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _11405_ (.A(_04485_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__xnor2_2 _11406_ (.A(_04485_),
    .B(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__o21ai_2 _11407_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04396_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand2b_1 _11408_ (.A_N(_04500_),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__xor2_2 _11409_ (.A(_04500_),
    .B(_04501_),
    .X(_04504_));
 sky130_fd_sc_hd__a21oi_2 _11410_ (.A1(_04398_),
    .A2(_04401_),
    .B1(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__nand3_2 _11411_ (.A(_04398_),
    .B(_04401_),
    .C(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2b_2 _11412_ (.A_N(_04505_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(_04297_),
    .B(_04406_),
    .Y(_04508_));
 sky130_fd_sc_hd__and2_1 _11414_ (.A(_04299_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__inv_2 _11415_ (.A(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__o21a_1 _11416_ (.A1(_04295_),
    .A2(_04403_),
    .B1(_04404_),
    .X(_04511_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(_04298_),
    .A2(_04508_),
    .B1(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__a21oi_1 _11418_ (.A1(_04086_),
    .A2(_04509_),
    .B1(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__o31ai_4 _11419_ (.A1(_03624_),
    .A2(_04088_),
    .A3(_04510_),
    .B1(_04513_),
    .Y(_04515_));
 sky130_fd_sc_hd__xnor2_4 _11420_ (.A(_04507_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__a21oi_1 _11421_ (.A1(_04446_),
    .A2(_04516_),
    .B1(net187),
    .Y(_04517_));
 sky130_fd_sc_hd__o21ai_1 _11422_ (.A1(_04446_),
    .A2(_04516_),
    .B1(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__o21a_1 _11423_ (.A1(net157),
    .A2(_01847_),
    .B1(_01850_),
    .X(_04519_));
 sky130_fd_sc_hd__o31ai_2 _11424_ (.A1(net157),
    .A2(_01847_),
    .A3(_01850_),
    .B1(net233),
    .Y(_04520_));
 sky130_fd_sc_hd__a21o_1 _11425_ (.A1(_05910_),
    .A2(_04418_),
    .B1(_05892_),
    .X(_04521_));
 sky130_fd_sc_hd__nand2_1 _11426_ (.A(net284),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21a_1 _11427_ (.A1(net284),
    .A2(_06375_),
    .B1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__xnor2_1 _11428_ (.A(_05857_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__o21a_1 _11429_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04424_),
    .X(_04525_));
 sky130_fd_sc_hd__nor2_1 _11430_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04526_));
 sky130_fd_sc_hd__nand2_1 _11431_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2b_1 _11432_ (.A_N(_04526_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__xnor2_1 _11433_ (.A(_04525_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(_04226_),
    .A1(_04529_),
    .S(net250),
    .X(_04530_));
 sky130_fd_sc_hd__a21o_1 _11435_ (.A1(_05838_),
    .A2(_02325_),
    .B1(_02321_),
    .X(_04531_));
 sky130_fd_sc_hd__o2bb2a_1 _11436_ (.A1_N(_05848_),
    .A2_N(_04531_),
    .B1(net185),
    .B2(_05838_),
    .X(_04532_));
 sky130_fd_sc_hd__o221a_1 _11437_ (.A1(net168),
    .A2(_04215_),
    .B1(_04226_),
    .B2(_02320_),
    .C1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__o21a_1 _11438_ (.A1(\div_shifter[48] ),
    .A2(_04430_),
    .B1(net226),
    .X(_04534_));
 sky130_fd_sc_hd__xnor2_1 _11439_ (.A(\div_shifter[49] ),
    .B(_04534_),
    .Y(_04536_));
 sky130_fd_sc_hd__o21a_1 _11440_ (.A1(\div_res[16] ),
    .A2(_04436_),
    .B1(net163),
    .X(_04537_));
 sky130_fd_sc_hd__xnor2_1 _11441_ (.A(\div_res[17] ),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__o22a_1 _11442_ (.A1(net231),
    .A2(_04536_),
    .B1(_04538_),
    .B2(net183),
    .X(_04539_));
 sky130_fd_sc_hd__o211a_1 _11443_ (.A1(net196),
    .A2(_04530_),
    .B1(_04533_),
    .C1(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__o221a_1 _11444_ (.A1(_04519_),
    .A2(_04520_),
    .B1(_04524_),
    .B2(net236),
    .C1(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__a21oi_1 _11445_ (.A1(_04518_),
    .A2(_04541_),
    .B1(_06463_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_1 _11446_ (.A(_05829_),
    .B(net241),
    .Y(_04543_));
 sky130_fd_sc_hd__a21oi_1 _11447_ (.A1(curr_PC[16]),
    .A2(_04337_),
    .B1(curr_PC[17]),
    .Y(_04544_));
 sky130_fd_sc_hd__and3_1 _11448_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04337_),
    .X(_04545_));
 sky130_fd_sc_hd__o21ai_2 _11449_ (.A1(_04544_),
    .A2(_04545_),
    .B1(net248),
    .Y(_04546_));
 sky130_fd_sc_hd__o31a_4 _11450_ (.A1(net248),
    .A2(_04542_),
    .A3(_04543_),
    .B1(_04546_),
    .X(dest_val[17]));
 sky130_fd_sc_hd__or2_1 _11451_ (.A(_04412_),
    .B(_04516_),
    .X(_04547_));
 sky130_fd_sc_hd__or4_2 _11452_ (.A(_03657_),
    .B(_04124_),
    .C(_04339_),
    .D(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_00307_),
    .B(net8),
    .Y(_04549_));
 sky130_fd_sc_hd__a22o_2 _11454_ (.A1(_00311_),
    .A2(net8),
    .B1(_04549_),
    .B2(net88),
    .X(_04550_));
 sky130_fd_sc_hd__o21a_1 _11455_ (.A1(net101),
    .A2(net18),
    .B1(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__nor3_1 _11456_ (.A(net101),
    .B(net18),
    .C(_04550_),
    .Y(_04552_));
 sky130_fd_sc_hd__nor2_1 _11457_ (.A(_04551_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__nor2_1 _11458_ (.A(_04450_),
    .B(_04454_),
    .Y(_04554_));
 sky130_fd_sc_hd__o21a_1 _11459_ (.A1(_04450_),
    .A2(_04454_),
    .B1(_04553_),
    .X(_04556_));
 sky130_fd_sc_hd__xnor2_2 _11460_ (.A(_04553_),
    .B(_04554_),
    .Y(_04557_));
 sky130_fd_sc_hd__a22o_1 _11461_ (.A1(_06492_),
    .A2(net38),
    .B1(net36),
    .B2(_06500_),
    .X(_04558_));
 sky130_fd_sc_hd__xor2_1 _11462_ (.A(net89),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__a22o_1 _11463_ (.A1(net29),
    .A2(_00690_),
    .B1(_01954_),
    .B2(net31),
    .X(_04560_));
 sky130_fd_sc_hd__xnor2_1 _11464_ (.A(_00202_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__and2_1 _11465_ (.A(_04559_),
    .B(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__nor2_1 _11466_ (.A(_04559_),
    .B(_04561_),
    .Y(_04563_));
 sky130_fd_sc_hd__nor2_1 _11467_ (.A(_04562_),
    .B(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__o22a_1 _11468_ (.A1(net54),
    .A2(net44),
    .B1(net16),
    .B2(net46),
    .X(_04565_));
 sky130_fd_sc_hd__xnor2_2 _11469_ (.A(net95),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__xor2_2 _11470_ (.A(_04564_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__nand2_1 _11471_ (.A(_04557_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__xnor2_2 _11472_ (.A(_04557_),
    .B(_04567_),
    .Y(_04569_));
 sky130_fd_sc_hd__o22a_1 _11473_ (.A1(net63),
    .A2(net22),
    .B1(net14),
    .B2(net61),
    .X(_04570_));
 sky130_fd_sc_hd__xnor2_2 _11474_ (.A(net68),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__o22a_1 _11475_ (.A1(net53),
    .A2(net9),
    .B1(net4),
    .B2(net51),
    .X(_04572_));
 sky130_fd_sc_hd__xnor2_1 _11476_ (.A(net18),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__a22o_1 _11477_ (.A1(_06534_),
    .A2(net42),
    .B1(net40),
    .B2(_06538_),
    .X(_04574_));
 sky130_fd_sc_hd__xor2_1 _11478_ (.A(net92),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__nand2b_1 _11479_ (.A_N(_04573_),
    .B(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__nand2b_1 _11480_ (.A_N(_04575_),
    .B(_04573_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _11481_ (.A(_04577_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__xnor2_2 _11482_ (.A(_04571_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__xor2_2 _11483_ (.A(_04569_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__a21o_1 _11484_ (.A1(_04460_),
    .A2(_04471_),
    .B1(_04483_),
    .X(_04582_));
 sky130_fd_sc_hd__o31ai_4 _11485_ (.A1(net99),
    .A2(net18),
    .A3(_04477_),
    .B1(_04480_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _11486_ (.A(_04456_),
    .B(_04458_),
    .Y(_04584_));
 sky130_fd_sc_hd__a21oi_2 _11487_ (.A1(_04467_),
    .A2(_04469_),
    .B1(_04465_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21o_1 _11488_ (.A1(_04456_),
    .A2(_04458_),
    .B1(_04585_),
    .X(_04586_));
 sky130_fd_sc_hd__xnor2_2 _11489_ (.A(_04584_),
    .B(_04585_),
    .Y(_04587_));
 sky130_fd_sc_hd__xnor2_2 _11490_ (.A(_04583_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__a21oi_2 _11491_ (.A1(_04487_),
    .A2(_04490_),
    .B1(_04489_),
    .Y(_04589_));
 sky130_fd_sc_hd__xnor2_2 _11492_ (.A(_04588_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2b_1 _11493_ (.A_N(_04590_),
    .B(_04582_),
    .Y(_04591_));
 sky130_fd_sc_hd__xnor2_2 _11494_ (.A(_04582_),
    .B(_04590_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2_1 _11495_ (.A(_04581_),
    .B(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__xnor2_2 _11496_ (.A(_04581_),
    .B(_04592_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _11497_ (.A(_04495_),
    .B(_04497_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2b_1 _11498_ (.A_N(_04594_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__xor2_2 _11499_ (.A(_04594_),
    .B(_04595_),
    .X(_04598_));
 sky130_fd_sc_hd__a21oi_2 _11500_ (.A1(_04499_),
    .A2(_04502_),
    .B1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand3_2 _11501_ (.A(_04499_),
    .B(_04502_),
    .C(_04598_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2b_4 _11502_ (.A_N(_04599_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__o21a_1 _11503_ (.A1(_04403_),
    .A2(_04505_),
    .B1(_04506_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_1 _11504_ (.A(_04406_),
    .B(_04507_),
    .Y(_04603_));
 sky130_fd_sc_hd__a21o_1 _11505_ (.A1(_04407_),
    .A2(_04603_),
    .B1(_04602_),
    .X(_04604_));
 sky130_fd_sc_hd__and2_1 _11506_ (.A(_04408_),
    .B(_04603_),
    .X(_04605_));
 sky130_fd_sc_hd__a21o_1 _11507_ (.A1(_04196_),
    .A2(_04605_),
    .B1(_04604_),
    .X(_04606_));
 sky130_fd_sc_hd__xnor2_4 _11508_ (.A(_04601_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__a21oi_1 _11509_ (.A1(net164),
    .A2(_04548_),
    .B1(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__a31o_1 _11510_ (.A1(net164),
    .A2(_04548_),
    .A3(_04607_),
    .B1(net187),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(net159),
    .B(_01851_),
    .Y(_04610_));
 sky130_fd_sc_hd__xnor2_2 _11512_ (.A(_01856_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__or2_1 _11513_ (.A(net284),
    .B(_06377_),
    .X(_04612_));
 sky130_fd_sc_hd__a21bo_1 _11514_ (.A1(_05848_),
    .A2(_04521_),
    .B1_N(_05838_),
    .X(_04613_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(net284),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__a21oi_1 _11516_ (.A1(_04612_),
    .A2(_04614_),
    .B1(_05802_),
    .Y(_04615_));
 sky130_fd_sc_hd__a31o_1 _11517_ (.A1(_05802_),
    .A2(_04612_),
    .A3(_04614_),
    .B1(net236),
    .X(_04616_));
 sky130_fd_sc_hd__nand2_1 _11518_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04617_));
 sky130_fd_sc_hd__or2_1 _11519_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .X(_04619_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_04617_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__o21ai_1 _11521_ (.A1(_04525_),
    .A2(_04526_),
    .B1(_04527_),
    .Y(_04621_));
 sky130_fd_sc_hd__xnor2_1 _11522_ (.A(_04620_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(_04118_),
    .A1(_04622_),
    .S(net250),
    .X(_04623_));
 sky130_fd_sc_hd__or3_1 _11524_ (.A(\div_shifter[49] ),
    .B(\div_shifter[48] ),
    .C(_04430_),
    .X(_04624_));
 sky130_fd_sc_hd__a21oi_1 _11525_ (.A1(net226),
    .A2(_04624_),
    .B1(\div_shifter[50] ),
    .Y(_04625_));
 sky130_fd_sc_hd__a31o_1 _11526_ (.A1(\div_shifter[50] ),
    .A2(net226),
    .A3(_04624_),
    .B1(net231),
    .X(_04626_));
 sky130_fd_sc_hd__nor2_1 _11527_ (.A(_04625_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__or3_1 _11528_ (.A(\div_res[17] ),
    .B(\div_res[16] ),
    .C(_04436_),
    .X(_04628_));
 sky130_fd_sc_hd__nand3_1 _11529_ (.A(\div_res[18] ),
    .B(net163),
    .C(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a21o_1 _11530_ (.A1(net163),
    .A2(_04628_),
    .B1(\div_res[18] ),
    .X(_04630_));
 sky130_fd_sc_hd__mux2_1 _11531_ (.A0(net234),
    .A1(net185),
    .S(_05775_),
    .X(_04631_));
 sky130_fd_sc_hd__a21oi_1 _11532_ (.A1(net186),
    .A2(_04631_),
    .B1(_05784_),
    .Y(_04632_));
 sky130_fd_sc_hd__a221o_1 _11533_ (.A1(net170),
    .A2(_04106_),
    .B1(_04118_),
    .B2(_02319_),
    .C1(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__a31o_1 _11534_ (.A1(_02334_),
    .A2(_04629_),
    .A3(_04630_),
    .B1(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__a211o_1 _11535_ (.A1(net197),
    .A2(_04623_),
    .B1(_04627_),
    .C1(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__o21ba_1 _11536_ (.A1(_04615_),
    .A2(_04616_),
    .B1_N(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__o221a_1 _11537_ (.A1(_04608_),
    .A2(_04609_),
    .B1(_04611_),
    .B2(_02330_),
    .C1(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a2bb2o_1 _11538_ (.A1_N(_06463_),
    .A2_N(_04637_),
    .B1(_05766_),
    .B2(net242),
    .X(_04638_));
 sky130_fd_sc_hd__and2_2 _11539_ (.A(curr_PC[18]),
    .B(_04545_),
    .X(_04639_));
 sky130_fd_sc_hd__o21ai_1 _11540_ (.A1(curr_PC[18]),
    .A2(_04545_),
    .B1(net249),
    .Y(_04640_));
 sky130_fd_sc_hd__a2bb2o_4 _11541_ (.A1_N(_04639_),
    .A2_N(_04640_),
    .B1(net244),
    .B2(_04638_),
    .X(dest_val[18]));
 sky130_fd_sc_hd__or2_1 _11542_ (.A(_04548_),
    .B(_04607_),
    .X(_04641_));
 sky130_fd_sc_hd__o21ai_2 _11543_ (.A1(_04588_),
    .A2(_04589_),
    .B1(_04591_),
    .Y(_04642_));
 sky130_fd_sc_hd__o22a_1 _11544_ (.A1(net57),
    .A2(net22),
    .B1(net14),
    .B2(net63),
    .X(_04643_));
 sky130_fd_sc_hd__xnor2_1 _11545_ (.A(net68),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__a22o_1 _11546_ (.A1(_06553_),
    .A2(net38),
    .B1(net36),
    .B2(_06492_),
    .X(_04645_));
 sky130_fd_sc_hd__xor2_1 _11547_ (.A(net89),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__nand2b_1 _11548_ (.A_N(_04644_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2b_1 _11549_ (.A_N(_04646_),
    .B(_04644_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _11550_ (.A(_04647_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__a22o_1 _11551_ (.A1(_06500_),
    .A2(net42),
    .B1(net40),
    .B2(_06534_),
    .X(_04651_));
 sky130_fd_sc_hd__xor2_2 _11552_ (.A(net92),
    .B(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__nand2b_1 _11553_ (.A_N(_04650_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__xnor2_2 _11554_ (.A(_04650_),
    .B(_04652_),
    .Y(_04654_));
 sky130_fd_sc_hd__o22a_1 _11555_ (.A1(net44),
    .A2(net16),
    .B1(net13),
    .B2(net46),
    .X(_04655_));
 sky130_fd_sc_hd__xor2_2 _11556_ (.A(net95),
    .B(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__xnor2_1 _11557_ (.A(net88),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__a22o_1 _11558_ (.A1(net29),
    .A2(_01954_),
    .B1(net8),
    .B2(_00290_),
    .X(_04658_));
 sky130_fd_sc_hd__xnor2_1 _11559_ (.A(_00201_),
    .B(_04658_),
    .Y(_04660_));
 sky130_fd_sc_hd__or2_1 _11560_ (.A(_04657_),
    .B(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(_04657_),
    .B(_04660_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(_04661_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__o22a_1 _11563_ (.A1(net61),
    .A2(net9),
    .B1(net4),
    .B2(net53),
    .X(_04664_));
 sky130_fd_sc_hd__xnor2_1 _11564_ (.A(net21),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand2_1 _11565_ (.A(_04550_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__or2_1 _11566_ (.A(_04550_),
    .B(_04665_),
    .X(_04667_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(_04666_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _11568_ (.A(_00157_),
    .B(_02081_),
    .Y(_04669_));
 sky130_fd_sc_hd__xor2_2 _11569_ (.A(_04668_),
    .B(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__xnor2_1 _11570_ (.A(_04663_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__xor2_1 _11571_ (.A(_04654_),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__o21ai_2 _11572_ (.A1(_04569_),
    .A2(_04580_),
    .B1(_04568_),
    .Y(_04674_));
 sky130_fd_sc_hd__o21ai_1 _11573_ (.A1(_04571_),
    .A2(_04579_),
    .B1(_04577_),
    .Y(_04675_));
 sky130_fd_sc_hd__a21oi_1 _11574_ (.A1(_04564_),
    .A2(_04566_),
    .B1(_04562_),
    .Y(_04676_));
 sky130_fd_sc_hd__o21bai_2 _11575_ (.A1(_04552_),
    .A2(_04556_),
    .B1_N(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__or3b_1 _11576_ (.A(_04552_),
    .B(_04556_),
    .C_N(_04676_),
    .X(_04678_));
 sky130_fd_sc_hd__nand2_1 _11577_ (.A(_04677_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2b_1 _11578_ (.A_N(_04679_),
    .B(_04675_),
    .Y(_04680_));
 sky130_fd_sc_hd__xor2_1 _11579_ (.A(_04675_),
    .B(_04679_),
    .X(_04682_));
 sky130_fd_sc_hd__a21boi_1 _11580_ (.A1(_04583_),
    .A2(_04587_),
    .B1_N(_04586_),
    .Y(_04683_));
 sky130_fd_sc_hd__or2_1 _11581_ (.A(_04682_),
    .B(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__xnor2_1 _11582_ (.A(_04682_),
    .B(_04683_),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2b_1 _11583_ (.A_N(_04685_),
    .B(_04674_),
    .Y(_04686_));
 sky130_fd_sc_hd__xnor2_1 _11584_ (.A(_04674_),
    .B(_04685_),
    .Y(_04687_));
 sky130_fd_sc_hd__nand2_1 _11585_ (.A(_04673_),
    .B(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__or2_1 _11586_ (.A(_04673_),
    .B(_04687_),
    .X(_04689_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(_04688_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2b_1 _11588_ (.A_N(_04690_),
    .B(_04642_),
    .Y(_04691_));
 sky130_fd_sc_hd__xor2_2 _11589_ (.A(_04642_),
    .B(_04690_),
    .X(_04693_));
 sky130_fd_sc_hd__a21o_2 _11590_ (.A1(_04593_),
    .A2(_04596_),
    .B1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__inv_2 _11591_ (.A(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand3_2 _11592_ (.A(_04593_),
    .B(_04596_),
    .C(_04693_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_4 _11593_ (.A(_04694_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__o21a_1 _11594_ (.A1(_04505_),
    .A2(_04599_),
    .B1(_04600_),
    .X(_04698_));
 sky130_fd_sc_hd__nor2_1 _11595_ (.A(_04507_),
    .B(_04601_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_1 _11596_ (.A1(_04511_),
    .A2(_04699_),
    .B1(_04698_),
    .Y(_04700_));
 sky130_fd_sc_hd__and2_1 _11597_ (.A(_04508_),
    .B(_04699_),
    .X(_04701_));
 sky130_fd_sc_hd__inv_2 _11598_ (.A(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2_1 _11599_ (.A(_04300_),
    .B(_04701_),
    .Y(_04704_));
 sky130_fd_sc_hd__o311a_2 _11600_ (.A1(_03857_),
    .A2(_04301_),
    .A3(_04702_),
    .B1(_04704_),
    .C1(_04700_),
    .X(_04705_));
 sky130_fd_sc_hd__xor2_4 _11601_ (.A(_04697_),
    .B(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__a21oi_1 _11602_ (.A1(net164),
    .A2(_04641_),
    .B1(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__a31o_1 _11603_ (.A1(net164),
    .A2(_04641_),
    .A3(_04706_),
    .B1(net187),
    .X(_04708_));
 sky130_fd_sc_hd__or3_1 _11604_ (.A(net157),
    .B(_01857_),
    .C(_01860_),
    .X(_04709_));
 sky130_fd_sc_hd__o21ai_1 _11605_ (.A1(net157),
    .A2(_01857_),
    .B1(_01860_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_2 _11606_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__or2_1 _11607_ (.A(net284),
    .B(_06379_),
    .X(_04712_));
 sky130_fd_sc_hd__a21oi_1 _11608_ (.A1(_05793_),
    .A2(_04613_),
    .B1(_05775_),
    .Y(_04713_));
 sky130_fd_sc_hd__or2_1 _11609_ (.A(instruction[7]),
    .B(_04713_),
    .X(_04715_));
 sky130_fd_sc_hd__a21oi_1 _11610_ (.A1(_04712_),
    .A2(_04715_),
    .B1(_05728_),
    .Y(_04716_));
 sky130_fd_sc_hd__and3_1 _11611_ (.A(_05728_),
    .B(_04712_),
    .C(_04715_),
    .X(_04717_));
 sky130_fd_sc_hd__or3_1 _11612_ (.A(net236),
    .B(_04716_),
    .C(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04719_));
 sky130_fd_sc_hd__or2_1 _11614_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .X(_04720_));
 sky130_fd_sc_hd__nand2_1 _11615_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21bo_1 _11616_ (.A1(_04619_),
    .A2(_04621_),
    .B1_N(_04617_),
    .X(_04722_));
 sky130_fd_sc_hd__xnor2_1 _11617_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nor2_1 _11618_ (.A(net223),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__a211o_1 _11619_ (.A1(net224),
    .A2(_04007_),
    .B1(_04724_),
    .C1(_06449_),
    .X(_04726_));
 sky130_fd_sc_hd__or2_1 _11620_ (.A(\div_res[18] ),
    .B(_04628_),
    .X(_04727_));
 sky130_fd_sc_hd__a21oi_1 _11621_ (.A1(net163),
    .A2(_04727_),
    .B1(\div_res[19] ),
    .Y(_04728_));
 sky130_fd_sc_hd__a311o_1 _11622_ (.A1(\div_res[19] ),
    .A2(net163),
    .A3(_04727_),
    .B1(_04728_),
    .C1(net183),
    .X(_04729_));
 sky130_fd_sc_hd__or2_1 _11623_ (.A(\div_shifter[50] ),
    .B(_04624_),
    .X(_04730_));
 sky130_fd_sc_hd__a21oi_1 _11624_ (.A1(net226),
    .A2(_04730_),
    .B1(\div_shifter[51] ),
    .Y(_04731_));
 sky130_fd_sc_hd__a31o_1 _11625_ (.A1(\div_shifter[51] ),
    .A2(net226),
    .A3(_04730_),
    .B1(net231),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(net234),
    .A1(net185),
    .S(_05709_),
    .X(_04733_));
 sky130_fd_sc_hd__a21o_1 _11627_ (.A1(net186),
    .A2(_04733_),
    .B1(_05719_),
    .X(_04734_));
 sky130_fd_sc_hd__o221a_1 _11628_ (.A1(net168),
    .A2(_03989_),
    .B1(_04007_),
    .B2(_02320_),
    .C1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__o21a_1 _11629_ (.A1(_04731_),
    .A2(_04732_),
    .B1(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__and4_1 _11630_ (.A(_04718_),
    .B(_04726_),
    .C(_04729_),
    .D(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__o221a_1 _11631_ (.A1(_04707_),
    .A2(_04708_),
    .B1(_04711_),
    .B2(_02330_),
    .C1(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__o22a_1 _11632_ (.A1(_05700_),
    .A2(net241),
    .B1(_06463_),
    .B2(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__a21oi_1 _11633_ (.A1(curr_PC[19]),
    .A2(_04639_),
    .B1(net244),
    .Y(_04741_));
 sky130_fd_sc_hd__o21ai_2 _11634_ (.A1(curr_PC[19]),
    .A2(_04639_),
    .B1(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21ai_4 _11635_ (.A1(net248),
    .A2(_04740_),
    .B1(_04742_),
    .Y(dest_val[19]));
 sky130_fd_sc_hd__o31a_1 _11636_ (.A1(_04548_),
    .A2(_04607_),
    .A3(_04706_),
    .B1(net166),
    .X(_04743_));
 sky130_fd_sc_hd__o22a_1 _11637_ (.A1(net44),
    .A2(net13),
    .B1(net11),
    .B2(net46),
    .X(_04744_));
 sky130_fd_sc_hd__xnor2_1 _11638_ (.A(net95),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__a21oi_1 _11639_ (.A1(net29),
    .A2(net8),
    .B1(_00201_),
    .Y(_04747_));
 sky130_fd_sc_hd__a31o_1 _11640_ (.A1(_00201_),
    .A2(_00288_),
    .A3(net8),
    .B1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__and2b_1 _11641_ (.A_N(_04745_),
    .B(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__and2b_1 _11642_ (.A_N(_04748_),
    .B(_04745_),
    .X(_04750_));
 sky130_fd_sc_hd__nor2_1 _11643_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__o22a_1 _11644_ (.A1(net63),
    .A2(net9),
    .B1(net4),
    .B2(net61),
    .X(_04752_));
 sky130_fd_sc_hd__nand2_1 _11645_ (.A(net53),
    .B(net21),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_1 _11646_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__or2_1 _11647_ (.A(_04751_),
    .B(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__nand2_1 _11648_ (.A(_04751_),
    .B(_04754_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(_04755_),
    .B(_04756_),
    .Y(_04758_));
 sky130_fd_sc_hd__o22a_1 _11650_ (.A1(net59),
    .A2(net22),
    .B1(net14),
    .B2(net57),
    .X(_04759_));
 sky130_fd_sc_hd__xnor2_1 _11651_ (.A(net68),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__o22a_1 _11652_ (.A1(net54),
    .A2(_00252_),
    .B1(net16),
    .B2(_00248_),
    .X(_04761_));
 sky130_fd_sc_hd__xnor2_1 _11653_ (.A(net89),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__and2b_1 _11654_ (.A_N(_04760_),
    .B(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__xor2_1 _11655_ (.A(_04760_),
    .B(_04762_),
    .X(_04764_));
 sky130_fd_sc_hd__a22o_1 _11656_ (.A1(_06492_),
    .A2(net42),
    .B1(net40),
    .B2(_06500_),
    .X(_04765_));
 sky130_fd_sc_hd__xor2_1 _11657_ (.A(net92),
    .B(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__and2b_1 _11658_ (.A_N(_04764_),
    .B(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__and2b_1 _11659_ (.A_N(_04766_),
    .B(_04764_),
    .X(_04769_));
 sky130_fd_sc_hd__or2_1 _11660_ (.A(_04767_),
    .B(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__xor2_1 _11661_ (.A(_04758_),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__a32oi_2 _11662_ (.A1(_04661_),
    .A2(_04662_),
    .A3(_04671_),
    .B1(_04672_),
    .B2(_04654_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_04647_),
    .B(_04653_),
    .Y(_04773_));
 sky130_fd_sc_hd__o21ai_1 _11664_ (.A1(net88),
    .A2(_04656_),
    .B1(_04661_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21a_1 _11665_ (.A1(_04668_),
    .A2(_04669_),
    .B1(_04666_),
    .X(_04775_));
 sky130_fd_sc_hd__inv_2 _11666_ (.A(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand2_1 _11667_ (.A(_04774_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__xor2_1 _11668_ (.A(_04774_),
    .B(_04775_),
    .X(_04778_));
 sky130_fd_sc_hd__nand2b_1 _11669_ (.A_N(_04778_),
    .B(_04773_),
    .Y(_04780_));
 sky130_fd_sc_hd__xor2_1 _11670_ (.A(_04773_),
    .B(_04778_),
    .X(_04781_));
 sky130_fd_sc_hd__a21oi_1 _11671_ (.A1(_04677_),
    .A2(_04680_),
    .B1(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__and3_1 _11672_ (.A(_04677_),
    .B(_04680_),
    .C(_04781_),
    .X(_04783_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(_04782_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__and2b_1 _11674_ (.A_N(_04772_),
    .B(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__xnor2_1 _11675_ (.A(_04772_),
    .B(_04784_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_1 _11676_ (.A(_04771_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__xnor2_1 _11677_ (.A(_04771_),
    .B(_04786_),
    .Y(_04788_));
 sky130_fd_sc_hd__a21o_1 _11678_ (.A1(_04684_),
    .A2(_04686_),
    .B1(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__nand3_1 _11679_ (.A(_04684_),
    .B(_04686_),
    .C(_04788_),
    .Y(_04791_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(_04789_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__a21oi_1 _11681_ (.A1(_04688_),
    .A2(_04691_),
    .B1(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21o_1 _11682_ (.A1(_04688_),
    .A2(_04691_),
    .B1(_04792_),
    .X(_04794_));
 sky130_fd_sc_hd__and3_1 _11683_ (.A(_04688_),
    .B(_04691_),
    .C(_04792_),
    .X(_04795_));
 sky130_fd_sc_hd__or2_2 _11684_ (.A(_04793_),
    .B(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__o21a_1 _11685_ (.A1(_04599_),
    .A2(_04695_),
    .B1(_04696_),
    .X(_04797_));
 sky130_fd_sc_hd__nor2_2 _11686_ (.A(_04601_),
    .B(_04697_),
    .Y(_04798_));
 sky130_fd_sc_hd__a21o_1 _11687_ (.A1(_04602_),
    .A2(_04798_),
    .B1(_04797_),
    .X(_04799_));
 sky130_fd_sc_hd__a31oi_4 _11688_ (.A1(_04411_),
    .A2(_04603_),
    .A3(_04798_),
    .B1(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__xor2_2 _11689_ (.A(_04796_),
    .B(_04800_),
    .X(_04802_));
 sky130_fd_sc_hd__nor2_1 _11690_ (.A(_04743_),
    .B(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21o_1 _11691_ (.A1(_04743_),
    .A2(_04802_),
    .B1(net187),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_2 _11692_ (.A(net159),
    .B(_01861_),
    .Y(_04805_));
 sky130_fd_sc_hd__xnor2_4 _11693_ (.A(_01866_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__o21bai_1 _11694_ (.A1(_05728_),
    .A2(_04713_),
    .B1_N(_05709_),
    .Y(_04807_));
 sky130_fd_sc_hd__mux2_1 _11695_ (.A0(_06381_),
    .A1(_04807_),
    .S(net284),
    .X(_04808_));
 sky130_fd_sc_hd__o21ai_1 _11696_ (.A1(_05582_),
    .A2(_04808_),
    .B1(_02323_),
    .Y(_04809_));
 sky130_fd_sc_hd__a21o_1 _11697_ (.A1(_05582_),
    .A2(_04808_),
    .B1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__nand2_1 _11698_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04811_));
 sky130_fd_sc_hd__or2_1 _11699_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _11700_ (.A(_04811_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__a21bo_1 _11701_ (.A1(_04720_),
    .A2(_04722_),
    .B1_N(_04719_),
    .X(_04815_));
 sky130_fd_sc_hd__xnor2_1 _11702_ (.A(_04814_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nor2_1 _11703_ (.A(net223),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__a211o_1 _11704_ (.A1(net224),
    .A2(_03887_),
    .B1(_04817_),
    .C1(_06449_),
    .X(_04818_));
 sky130_fd_sc_hd__or2_1 _11705_ (.A(\div_res[19] ),
    .B(_04727_),
    .X(_04819_));
 sky130_fd_sc_hd__a21oi_1 _11706_ (.A1(net163),
    .A2(_04819_),
    .B1(\div_res[20] ),
    .Y(_04820_));
 sky130_fd_sc_hd__a311o_1 _11707_ (.A1(\div_res[20] ),
    .A2(net163),
    .A3(_04819_),
    .B1(_04820_),
    .C1(net184),
    .X(_04821_));
 sky130_fd_sc_hd__or2_1 _11708_ (.A(\div_shifter[51] ),
    .B(_04730_),
    .X(_04822_));
 sky130_fd_sc_hd__a21oi_1 _11709_ (.A1(net226),
    .A2(_04822_),
    .B1(\div_shifter[52] ),
    .Y(_04824_));
 sky130_fd_sc_hd__a31o_1 _11710_ (.A1(\div_shifter[52] ),
    .A2(net226),
    .A3(_04822_),
    .B1(net231),
    .X(_04825_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(net234),
    .A1(net185),
    .S(_05561_),
    .X(_04826_));
 sky130_fd_sc_hd__a21o_1 _11712_ (.A1(net186),
    .A2(_04826_),
    .B1(_05572_),
    .X(_04827_));
 sky130_fd_sc_hd__o221a_1 _11713_ (.A1(net168),
    .A2(_03875_),
    .B1(_03887_),
    .B2(_02320_),
    .C1(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__o21a_1 _11714_ (.A1(_04824_),
    .A2(_04825_),
    .B1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__and4_1 _11715_ (.A(_04810_),
    .B(_04818_),
    .C(_04821_),
    .D(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__o221a_1 _11716_ (.A1(_04803_),
    .A2(_04804_),
    .B1(_04806_),
    .B2(_02330_),
    .C1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__o22a_1 _11717_ (.A1(_05550_),
    .A2(net241),
    .B1(_06463_),
    .B2(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__and3_1 _11718_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04639_),
    .X(_04833_));
 sky130_fd_sc_hd__a21oi_1 _11719_ (.A1(curr_PC[19]),
    .A2(_04639_),
    .B1(curr_PC[20]),
    .Y(_04835_));
 sky130_fd_sc_hd__or3_2 _11720_ (.A(net244),
    .B(_04833_),
    .C(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__o21ai_4 _11721_ (.A1(net248),
    .A2(_04832_),
    .B1(_04836_),
    .Y(dest_val[20]));
 sky130_fd_sc_hd__o41a_1 _11722_ (.A1(_04548_),
    .A2(_04607_),
    .A3(_04706_),
    .A4(_04802_),
    .B1(net166),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _11723_ (.A(_04782_),
    .B(_04785_),
    .X(_04838_));
 sky130_fd_sc_hd__o22a_1 _11724_ (.A1(net65),
    .A2(net22),
    .B1(net14),
    .B2(net59),
    .X(_04839_));
 sky130_fd_sc_hd__xnor2_1 _11725_ (.A(net68),
    .B(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__o22a_1 _11726_ (.A1(net57),
    .A2(net9),
    .B1(net4),
    .B2(net63),
    .X(_04841_));
 sky130_fd_sc_hd__xnor2_1 _11727_ (.A(net18),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(_06553_),
    .A2(net42),
    .B1(net40),
    .B2(_06492_),
    .X(_04843_));
 sky130_fd_sc_hd__xor2_1 _11729_ (.A(net92),
    .B(_04843_),
    .X(_04845_));
 sky130_fd_sc_hd__nand2b_1 _11730_ (.A_N(_04842_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2b_1 _11731_ (.A_N(_04845_),
    .B(_04842_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _11732_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__xor2_1 _11733_ (.A(_04840_),
    .B(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__and3_1 _11734_ (.A(_00148_),
    .B(_02081_),
    .C(_04752_),
    .X(_04850_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_04849_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__or2_1 _11736_ (.A(_04849_),
    .B(_04850_),
    .X(_04852_));
 sky130_fd_sc_hd__nand2_1 _11737_ (.A(_04851_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__o22a_1 _11738_ (.A1(_00252_),
    .A2(net16),
    .B1(_00689_),
    .B2(_00248_),
    .X(_04854_));
 sky130_fd_sc_hd__xnor2_1 _11739_ (.A(net89),
    .B(_04854_),
    .Y(_04856_));
 sky130_fd_sc_hd__xnor2_1 _11740_ (.A(_00202_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__o22a_1 _11741_ (.A1(net44),
    .A2(net11),
    .B1(_02070_),
    .B2(net46),
    .X(_04858_));
 sky130_fd_sc_hd__xnor2_1 _11742_ (.A(net95),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__and2b_1 _11743_ (.A_N(_04857_),
    .B(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__and2b_1 _11744_ (.A_N(_04859_),
    .B(_04857_),
    .X(_04861_));
 sky130_fd_sc_hd__or2_1 _11745_ (.A(_04860_),
    .B(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__xor2_1 _11746_ (.A(_04853_),
    .B(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__o21a_1 _11747_ (.A1(_04758_),
    .A2(_04770_),
    .B1(_04755_),
    .X(_04864_));
 sky130_fd_sc_hd__nor2_1 _11748_ (.A(_04763_),
    .B(_04767_),
    .Y(_04865_));
 sky130_fd_sc_hd__nand2_1 _11749_ (.A(_06522_),
    .B(_02081_),
    .Y(_04867_));
 sky130_fd_sc_hd__nor2_1 _11750_ (.A(_04865_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__xnor2_1 _11751_ (.A(_04865_),
    .B(_04867_),
    .Y(_04869_));
 sky130_fd_sc_hd__nor2_1 _11752_ (.A(_04749_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__and2_1 _11753_ (.A(_04749_),
    .B(_04869_),
    .X(_04871_));
 sky130_fd_sc_hd__or2_1 _11754_ (.A(_04870_),
    .B(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__a21oi_1 _11755_ (.A1(_04777_),
    .A2(_04780_),
    .B1(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__and3_1 _11756_ (.A(_04777_),
    .B(_04780_),
    .C(_04872_),
    .X(_04874_));
 sky130_fd_sc_hd__nor2_1 _11757_ (.A(_04873_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__xnor2_1 _11758_ (.A(_04864_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__nand2_1 _11759_ (.A(_04863_),
    .B(_04876_),
    .Y(_04878_));
 sky130_fd_sc_hd__xor2_1 _11760_ (.A(_04863_),
    .B(_04876_),
    .X(_04879_));
 sky130_fd_sc_hd__nand2_1 _11761_ (.A(_04838_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__xnor2_1 _11762_ (.A(_04838_),
    .B(_04879_),
    .Y(_04881_));
 sky130_fd_sc_hd__a21o_1 _11763_ (.A1(_04787_),
    .A2(_04789_),
    .B1(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__and3_1 _11764_ (.A(_04787_),
    .B(_04789_),
    .C(_04881_),
    .X(_04883_));
 sky130_fd_sc_hd__inv_2 _11765_ (.A(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_2 _11766_ (.A(_04882_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nor2_1 _11767_ (.A(_04697_),
    .B(_04796_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_1 _11768_ (.A(_04699_),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__nand2b_1 _11769_ (.A_N(_04887_),
    .B(_04512_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21oi_2 _11770_ (.A1(_04694_),
    .A2(_04794_),
    .B1(_04795_),
    .Y(_04890_));
 sky130_fd_sc_hd__a21oi_1 _11771_ (.A1(_04698_),
    .A2(_04886_),
    .B1(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o311a_2 _11772_ (.A1(_04090_),
    .A2(_04510_),
    .A3(_04887_),
    .B1(_04889_),
    .C1(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__xor2_2 _11773_ (.A(_04885_),
    .B(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__nor2_1 _11774_ (.A(_04837_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a21o_1 _11775_ (.A1(_04837_),
    .A2(_04893_),
    .B1(net187),
    .X(_04895_));
 sky130_fd_sc_hd__or2_1 _11776_ (.A(net157),
    .B(_01867_),
    .X(_04896_));
 sky130_fd_sc_hd__nor2_1 _11777_ (.A(_01870_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__a21o_1 _11778_ (.A1(_01870_),
    .A2(_04896_),
    .B1(_02330_),
    .X(_04898_));
 sky130_fd_sc_hd__o21a_1 _11779_ (.A1(_05582_),
    .A2(_06381_),
    .B1(_06383_),
    .X(_04900_));
 sky130_fd_sc_hd__a21o_1 _11780_ (.A1(_05582_),
    .A2(_04807_),
    .B1(_05561_),
    .X(_04901_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(_04900_),
    .A1(_04901_),
    .S(net284),
    .X(_04902_));
 sky130_fd_sc_hd__xnor2_1 _11782_ (.A(_05652_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _11783_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04904_));
 sky130_fd_sc_hd__or2_1 _11784_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .X(_04905_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_04904_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21bo_1 _11786_ (.A1(_04813_),
    .A2(_04815_),
    .B1_N(_04811_),
    .X(_04907_));
 sky130_fd_sc_hd__xnor2_1 _11787_ (.A(_04906_),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(net223),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a211o_1 _11789_ (.A1(net224),
    .A2(_03769_),
    .B1(_04909_),
    .C1(net196),
    .X(_04911_));
 sky130_fd_sc_hd__or2_1 _11790_ (.A(\div_shifter[52] ),
    .B(_04822_),
    .X(_04912_));
 sky130_fd_sc_hd__a21oi_1 _11791_ (.A1(net226),
    .A2(_04912_),
    .B1(\div_shifter[53] ),
    .Y(_04913_));
 sky130_fd_sc_hd__a31o_1 _11792_ (.A1(\div_shifter[53] ),
    .A2(net227),
    .A3(_04912_),
    .B1(net231),
    .X(_04914_));
 sky130_fd_sc_hd__or2_1 _11793_ (.A(_04913_),
    .B(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__or2_1 _11794_ (.A(\div_res[20] ),
    .B(_04819_),
    .X(_04916_));
 sky130_fd_sc_hd__a21oi_1 _11795_ (.A1(net163),
    .A2(_04916_),
    .B1(\div_res[21] ),
    .Y(_04917_));
 sky130_fd_sc_hd__a31o_1 _11796_ (.A1(\div_res[21] ),
    .A2(net163),
    .A3(_04916_),
    .B1(net184),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(net234),
    .A1(net185),
    .S(_05633_),
    .X(_04919_));
 sky130_fd_sc_hd__a21o_1 _11798_ (.A1(net186),
    .A2(_04919_),
    .B1(_05642_),
    .X(_04920_));
 sky130_fd_sc_hd__o221a_1 _11799_ (.A1(net168),
    .A2(_03756_),
    .B1(_03769_),
    .B2(_02320_),
    .C1(_04920_),
    .X(_04922_));
 sky130_fd_sc_hd__o211a_1 _11800_ (.A1(_04917_),
    .A2(_04918_),
    .B1(_04922_),
    .C1(_04915_),
    .X(_04923_));
 sky130_fd_sc_hd__o211a_1 _11801_ (.A1(net236),
    .A2(_04903_),
    .B1(_04911_),
    .C1(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__o221a_1 _11802_ (.A1(_04894_),
    .A2(_04895_),
    .B1(_04897_),
    .B2(_04898_),
    .C1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o22a_1 _11803_ (.A1(_05614_),
    .A2(net241),
    .B1(_06463_),
    .B2(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__nor2_1 _11804_ (.A(curr_PC[21]),
    .B(_04833_),
    .Y(_04927_));
 sky130_fd_sc_hd__and2_1 _11805_ (.A(curr_PC[21]),
    .B(_04833_),
    .X(_04928_));
 sky130_fd_sc_hd__or3_2 _11806_ (.A(net246),
    .B(_04927_),
    .C(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__o21ai_4 _11807_ (.A1(net249),
    .A2(_04926_),
    .B1(_04929_),
    .Y(dest_val[21]));
 sky130_fd_sc_hd__nor4_1 _11808_ (.A(_04547_),
    .B(_04607_),
    .C(_04802_),
    .D(_04893_),
    .Y(_04930_));
 sky130_fd_sc_hd__nor4_1 _11809_ (.A(_03657_),
    .B(_04124_),
    .C(_04339_),
    .D(_04706_),
    .Y(_04932_));
 sky130_fd_sc_hd__a21o_1 _11810_ (.A1(_04930_),
    .A2(_04932_),
    .B1(net158),
    .X(_04933_));
 sky130_fd_sc_hd__o21bai_1 _11811_ (.A1(_04864_),
    .A2(_04874_),
    .B1_N(_04873_),
    .Y(_04934_));
 sky130_fd_sc_hd__o22a_1 _11812_ (.A1(net66),
    .A2(net22),
    .B1(net14),
    .B2(net65),
    .X(_04935_));
 sky130_fd_sc_hd__xnor2_1 _11813_ (.A(_00668_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__a22oi_1 _11814_ (.A1(_06553_),
    .A2(net40),
    .B1(_00398_),
    .B2(net42),
    .Y(_04937_));
 sky130_fd_sc_hd__xnor2_1 _11815_ (.A(net92),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _11816_ (.A(_04936_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__or2_1 _11817_ (.A(_04936_),
    .B(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__nand2_1 _11818_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21a_1 _11819_ (.A1(_04840_),
    .A2(_04848_),
    .B1(_04846_),
    .X(_04943_));
 sky130_fd_sc_hd__xnor2_1 _11820_ (.A(_04941_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a22o_1 _11821_ (.A1(net37),
    .A2(_00690_),
    .B1(_01954_),
    .B2(net38),
    .X(_04945_));
 sky130_fd_sc_hd__xor2_1 _11822_ (.A(net89),
    .B(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__or2_1 _11823_ (.A(_00207_),
    .B(net6),
    .X(_04947_));
 sky130_fd_sc_hd__a22o_1 _11824_ (.A1(_00213_),
    .A2(net8),
    .B1(_04947_),
    .B2(net95),
    .X(_04948_));
 sky130_fd_sc_hd__or2_1 _11825_ (.A(_04946_),
    .B(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__nand2_1 _11826_ (.A(_04946_),
    .B(_04948_),
    .Y(_04950_));
 sky130_fd_sc_hd__and2_1 _11827_ (.A(_04949_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__or2_1 _11828_ (.A(_04944_),
    .B(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__nand2_1 _11829_ (.A(_04944_),
    .B(_04951_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _11830_ (.A(_04952_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__o21ai_1 _11831_ (.A1(_04853_),
    .A2(_04862_),
    .B1(_04851_),
    .Y(_04956_));
 sky130_fd_sc_hd__a21oi_1 _11832_ (.A1(_00202_),
    .A2(_04856_),
    .B1(_04860_),
    .Y(_04957_));
 sky130_fd_sc_hd__o22a_1 _11833_ (.A1(net59),
    .A2(net9),
    .B1(net4),
    .B2(net57),
    .X(_04958_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(net17),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nor2_1 _11835_ (.A(_04957_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__xnor2_1 _11836_ (.A(_04957_),
    .B(_04959_),
    .Y(_04961_));
 sky130_fd_sc_hd__nor2_1 _11837_ (.A(net63),
    .B(net18),
    .Y(_04962_));
 sky130_fd_sc_hd__and2b_1 _11838_ (.A_N(_04961_),
    .B(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__xnor2_1 _11839_ (.A(_04961_),
    .B(_04962_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21a_1 _11840_ (.A1(_04868_),
    .A2(_04870_),
    .B1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__nor3_1 _11841_ (.A(_04868_),
    .B(_04870_),
    .C(_04965_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor2_1 _11842_ (.A(_04966_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__xnor2_1 _11843_ (.A(_04956_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__or2_1 _11844_ (.A(_04955_),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_04955_),
    .B(_04969_),
    .Y(_04971_));
 sky130_fd_sc_hd__and2_1 _11846_ (.A(_04970_),
    .B(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(_04934_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__xnor2_1 _11848_ (.A(_04934_),
    .B(_04972_),
    .Y(_04974_));
 sky130_fd_sc_hd__a21o_1 _11849_ (.A1(_04878_),
    .A2(_04880_),
    .B1(_04974_),
    .X(_04976_));
 sky130_fd_sc_hd__and3_1 _11850_ (.A(_04878_),
    .B(_04880_),
    .C(_04974_),
    .X(_04977_));
 sky130_fd_sc_hd__inv_2 _11851_ (.A(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand2_2 _11852_ (.A(_04976_),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__a21oi_2 _11853_ (.A1(_04794_),
    .A2(_04882_),
    .B1(_04883_),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_2 _11854_ (.A(_04796_),
    .B(_04885_),
    .Y(_04981_));
 sky130_fd_sc_hd__a21o_1 _11855_ (.A1(_04797_),
    .A2(_04981_),
    .B1(_04980_),
    .X(_04982_));
 sky130_fd_sc_hd__nand2_1 _11856_ (.A(_04798_),
    .B(_04981_),
    .Y(_04983_));
 sky130_fd_sc_hd__inv_2 _11857_ (.A(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__a31o_1 _11858_ (.A1(_04604_),
    .A2(_04798_),
    .A3(_04981_),
    .B1(_04982_),
    .X(_04985_));
 sky130_fd_sc_hd__a31oi_4 _11859_ (.A1(_04196_),
    .A2(_04605_),
    .A3(_04984_),
    .B1(_04985_),
    .Y(_04987_));
 sky130_fd_sc_hd__xnor2_2 _11860_ (.A(_04979_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__and2_1 _11861_ (.A(_04933_),
    .B(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(_04933_),
    .B(_04988_),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _11863_ (.A(net159),
    .B(_01871_),
    .Y(_04991_));
 sky130_fd_sc_hd__xnor2_2 _11864_ (.A(_01877_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__a21o_1 _11865_ (.A1(_05652_),
    .A2(_04901_),
    .B1(_05633_),
    .X(_04993_));
 sky130_fd_sc_hd__o21a_1 _11866_ (.A1(_05652_),
    .A2(_04900_),
    .B1(_06382_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(_04993_),
    .A1(_04994_),
    .S(instruction[7]),
    .X(_04995_));
 sky130_fd_sc_hd__o21ai_1 _11868_ (.A1(_05518_),
    .A2(_04995_),
    .B1(_02323_),
    .Y(_04996_));
 sky130_fd_sc_hd__a21o_1 _11869_ (.A1(_05518_),
    .A2(_04995_),
    .B1(_04996_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _11870_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_04999_));
 sky130_fd_sc_hd__or2_1 _11871_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .X(_05000_));
 sky130_fd_sc_hd__nand2_1 _11872_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21bo_1 _11873_ (.A1(_04905_),
    .A2(_04907_),
    .B1_N(_04904_),
    .X(_05002_));
 sky130_fd_sc_hd__xnor2_1 _11874_ (.A(_05001_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(net223),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__a211o_1 _11876_ (.A1(net223),
    .A2(_03652_),
    .B1(_05004_),
    .C1(_06449_),
    .X(_05005_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(\div_shifter[53] ),
    .B(_04912_),
    .X(_05006_));
 sky130_fd_sc_hd__a21oi_1 _11878_ (.A1(net226),
    .A2(_05006_),
    .B1(\div_shifter[54] ),
    .Y(_05007_));
 sky130_fd_sc_hd__a31o_1 _11879_ (.A1(\div_shifter[54] ),
    .A2(net226),
    .A3(_05006_),
    .B1(net231),
    .X(_05009_));
 sky130_fd_sc_hd__or2_1 _11880_ (.A(\div_res[21] ),
    .B(_04916_),
    .X(_05010_));
 sky130_fd_sc_hd__a21oi_1 _11881_ (.A1(net163),
    .A2(_05010_),
    .B1(\div_res[22] ),
    .Y(_05011_));
 sky130_fd_sc_hd__a31o_1 _11882_ (.A1(\div_res[22] ),
    .A2(net163),
    .A3(_05010_),
    .B1(net184),
    .X(_05012_));
 sky130_fd_sc_hd__mux2_1 _11883_ (.A0(_02325_),
    .A1(_02331_),
    .S(_05496_),
    .X(_05013_));
 sky130_fd_sc_hd__o22a_1 _11884_ (.A1(reg1_val[22]),
    .A2(_05485_),
    .B1(_02321_),
    .B2(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__a221o_1 _11885_ (.A1(net170),
    .A2(_03640_),
    .B1(_03653_),
    .B2(_02319_),
    .C1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__o21ba_1 _11886_ (.A1(_05011_),
    .A2(_05012_),
    .B1_N(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__o211a_1 _11887_ (.A1(_05007_),
    .A2(_05009_),
    .B1(_05016_),
    .C1(_05005_),
    .X(_05017_));
 sky130_fd_sc_hd__o211a_1 _11888_ (.A1(_02330_),
    .A2(_04992_),
    .B1(_04998_),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__o31a_1 _11889_ (.A1(net187),
    .A2(_04989_),
    .A3(_04990_),
    .B1(_05018_),
    .X(_05020_));
 sky130_fd_sc_hd__o22a_1 _11890_ (.A1(_05474_),
    .A2(net241),
    .B1(_06463_),
    .B2(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__nor2_1 _11891_ (.A(curr_PC[22]),
    .B(_04928_),
    .Y(_05022_));
 sky130_fd_sc_hd__and3_1 _11892_ (.A(curr_PC[21]),
    .B(curr_PC[22]),
    .C(_04833_),
    .X(_05023_));
 sky130_fd_sc_hd__or3_2 _11893_ (.A(net246),
    .B(_05022_),
    .C(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o21ai_4 _11894_ (.A1(net249),
    .A2(_05021_),
    .B1(_05024_),
    .Y(dest_val[22]));
 sky130_fd_sc_hd__a31o_1 _11895_ (.A1(_04930_),
    .A2(_04932_),
    .A3(_04988_),
    .B1(net158),
    .X(_05025_));
 sky130_fd_sc_hd__a21o_1 _11896_ (.A1(_04956_),
    .A2(_04968_),
    .B1(_04966_),
    .X(_05026_));
 sky130_fd_sc_hd__a22o_1 _11897_ (.A1(net40),
    .A2(_00398_),
    .B1(_00690_),
    .B2(net42),
    .X(_05027_));
 sky130_fd_sc_hd__xor2_1 _11898_ (.A(net92),
    .B(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__and2b_1 _11899_ (.A_N(net95),
    .B(_05028_),
    .X(_05030_));
 sky130_fd_sc_hd__xor2_1 _11900_ (.A(net95),
    .B(_05028_),
    .X(_05031_));
 sky130_fd_sc_hd__o22a_1 _11901_ (.A1(_00252_),
    .A2(net11),
    .B1(net6),
    .B2(_00248_),
    .X(_05032_));
 sky130_fd_sc_hd__xnor2_1 _11902_ (.A(net89),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__and2b_1 _11903_ (.A_N(_05031_),
    .B(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__and2b_1 _11904_ (.A_N(_05033_),
    .B(_05031_),
    .X(_05035_));
 sky130_fd_sc_hd__or2_1 _11905_ (.A(_05034_),
    .B(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__nand2b_1 _11906_ (.A_N(_05036_),
    .B(_04949_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2b_1 _11907_ (.A_N(_04949_),
    .B(_05036_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _11908_ (.A(_05037_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__or2_1 _11909_ (.A(_04939_),
    .B(_05039_),
    .X(_05041_));
 sky130_fd_sc_hd__nand2_1 _11910_ (.A(_04939_),
    .B(_05039_),
    .Y(_05042_));
 sky130_fd_sc_hd__and2_1 _11911_ (.A(_05041_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__o21a_1 _11912_ (.A1(_04941_),
    .A2(_04943_),
    .B1(_04952_),
    .X(_05044_));
 sky130_fd_sc_hd__o22a_1 _11913_ (.A1(net65),
    .A2(net9),
    .B1(net4),
    .B2(net59),
    .X(_05045_));
 sky130_fd_sc_hd__xnor2_1 _11914_ (.A(net18),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__o22a_1 _11915_ (.A1(net54),
    .A2(net22),
    .B1(net14),
    .B2(net66),
    .X(_05047_));
 sky130_fd_sc_hd__xnor2_1 _11916_ (.A(net68),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__and3b_1 _11917_ (.A_N(_05048_),
    .B(_06538_),
    .C(_02081_),
    .X(_05049_));
 sky130_fd_sc_hd__o21a_1 _11918_ (.A1(net57),
    .A2(net18),
    .B1(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__nor2_1 _11919_ (.A(_05049_),
    .B(_05050_),
    .Y(_05052_));
 sky130_fd_sc_hd__and2b_1 _11920_ (.A_N(_05046_),
    .B(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__xnor2_1 _11921_ (.A(_05046_),
    .B(_05052_),
    .Y(_05054_));
 sky130_fd_sc_hd__o21ai_1 _11922_ (.A1(_04960_),
    .A2(_04963_),
    .B1(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__or3_1 _11923_ (.A(_04960_),
    .B(_04963_),
    .C(_05054_),
    .X(_05056_));
 sky130_fd_sc_hd__and2_1 _11924_ (.A(_05055_),
    .B(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__nand2b_1 _11925_ (.A_N(_05044_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__xnor2_1 _11926_ (.A(_05044_),
    .B(_05057_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11927_ (.A(_05043_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__xor2_1 _11928_ (.A(_05043_),
    .B(_05059_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_1 _11929_ (.A(_05026_),
    .B(_05061_),
    .Y(_05063_));
 sky130_fd_sc_hd__or2_1 _11930_ (.A(_05026_),
    .B(_05061_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _11931_ (.A(_05063_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__a21o_1 _11932_ (.A1(_04970_),
    .A2(_04973_),
    .B1(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__and3_1 _11933_ (.A(_04970_),
    .B(_04973_),
    .C(_05065_),
    .X(_05067_));
 sky130_fd_sc_hd__inv_2 _11934_ (.A(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__nand2_2 _11935_ (.A(_05066_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__a21oi_1 _11936_ (.A1(_04882_),
    .A2(_04976_),
    .B1(_04977_),
    .Y(_05070_));
 sky130_fd_sc_hd__nor2_1 _11937_ (.A(_04885_),
    .B(_04979_),
    .Y(_05071_));
 sky130_fd_sc_hd__a21o_1 _11938_ (.A1(_04890_),
    .A2(_05071_),
    .B1(_05070_),
    .X(_05072_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(_04886_),
    .B(_05071_),
    .Y(_05074_));
 sky130_fd_sc_hd__o21ba_1 _11940_ (.A1(_04705_),
    .A2(_05074_),
    .B1_N(_05072_),
    .X(_05075_));
 sky130_fd_sc_hd__xnor2_2 _11941_ (.A(_05069_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a21oi_1 _11942_ (.A1(_05025_),
    .A2(_05076_),
    .B1(_02246_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21a_1 _11943_ (.A1(_05025_),
    .A2(_05076_),
    .B1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a31o_1 _11944_ (.A1(_01867_),
    .A2(_01870_),
    .A3(_01877_),
    .B1(net157),
    .X(_05079_));
 sky130_fd_sc_hd__xor2_1 _11945_ (.A(_01879_),
    .B(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__nor2_2 _11946_ (.A(_02330_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__or2_1 _11947_ (.A(_05518_),
    .B(_04994_),
    .X(_05082_));
 sky130_fd_sc_hd__a21oi_1 _11948_ (.A1(reg1_val[22]),
    .A2(_05474_),
    .B1(net285),
    .Y(_05083_));
 sky130_fd_sc_hd__a21o_1 _11949_ (.A1(_05518_),
    .A2(_04993_),
    .B1(_05496_),
    .X(_05085_));
 sky130_fd_sc_hd__a22o_1 _11950_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_05085_),
    .B2(net286),
    .X(_05086_));
 sky130_fd_sc_hd__nand2_1 _11951_ (.A(_05442_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__o211a_1 _11952_ (.A1(_05442_),
    .A2(_05086_),
    .B1(_05087_),
    .C1(_02323_),
    .X(_05088_));
 sky130_fd_sc_hd__and2_1 _11953_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05089_));
 sky130_fd_sc_hd__or2_1 _11954_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05090_));
 sky130_fd_sc_hd__nand2b_1 _11955_ (.A_N(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21bo_1 _11956_ (.A1(_05000_),
    .A2(_05002_),
    .B1_N(_04999_),
    .X(_05092_));
 sky130_fd_sc_hd__xnor2_1 _11957_ (.A(_05091_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__nor2_1 _11958_ (.A(net223),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__a211o_1 _11959_ (.A1(net223),
    .A2(_03523_),
    .B1(_05094_),
    .C1(_06449_),
    .X(_05096_));
 sky130_fd_sc_hd__or2_1 _11960_ (.A(\div_res[22] ),
    .B(_05010_),
    .X(_05097_));
 sky130_fd_sc_hd__a21oi_1 _11961_ (.A1(net164),
    .A2(_05097_),
    .B1(\div_res[23] ),
    .Y(_05098_));
 sky130_fd_sc_hd__a311o_1 _11962_ (.A1(\div_res[23] ),
    .A2(net164),
    .A3(_05097_),
    .B1(_05098_),
    .C1(net184),
    .X(_05099_));
 sky130_fd_sc_hd__or2_1 _11963_ (.A(\div_shifter[54] ),
    .B(_05006_),
    .X(_05100_));
 sky130_fd_sc_hd__a21oi_1 _11964_ (.A1(net227),
    .A2(_05100_),
    .B1(\div_shifter[55] ),
    .Y(_05101_));
 sky130_fd_sc_hd__a31o_1 _11965_ (.A1(\div_shifter[55] ),
    .A2(net227),
    .A3(_05100_),
    .B1(net231),
    .X(_05102_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_05420_),
    .B(_02331_),
    .Y(_05103_));
 sky130_fd_sc_hd__o211a_1 _11967_ (.A1(_05420_),
    .A2(net235),
    .B1(_05103_),
    .C1(_02322_),
    .X(_05104_));
 sky130_fd_sc_hd__o22a_1 _11968_ (.A1(_05410_),
    .A2(net241),
    .B1(_05104_),
    .B2(_05431_),
    .X(_05105_));
 sky130_fd_sc_hd__o221a_1 _11969_ (.A1(net168),
    .A2(_03512_),
    .B1(_03523_),
    .B2(_02320_),
    .C1(_05105_),
    .X(_05107_));
 sky130_fd_sc_hd__o21a_1 _11970_ (.A1(_05101_),
    .A2(_05102_),
    .B1(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__and3_1 _11971_ (.A(_05096_),
    .B(_05099_),
    .C(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__or4b_2 _11972_ (.A(_05078_),
    .B(_05081_),
    .C(_05088_),
    .D_N(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__or2_1 _11973_ (.A(curr_PC[23]),
    .B(_05023_),
    .X(_05111_));
 sky130_fd_sc_hd__and2_1 _11974_ (.A(curr_PC[23]),
    .B(_05023_),
    .X(_05112_));
 sky130_fd_sc_hd__nor2_1 _11975_ (.A(net247),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__a22o_4 _11976_ (.A1(net247),
    .A2(_05110_),
    .B1(_05111_),
    .B2(_05113_),
    .X(dest_val[23]));
 sky130_fd_sc_hd__o31a_1 _11977_ (.A1(net95),
    .A2(_00244_),
    .A3(net6),
    .B1(net89),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_1 _11978_ (.A(net89),
    .B(net6),
    .Y(_05115_));
 sky130_fd_sc_hd__a21o_1 _11979_ (.A1(_00245_),
    .A2(_05115_),
    .B1(_05114_),
    .X(_05117_));
 sky130_fd_sc_hd__nor2_1 _11980_ (.A(net59),
    .B(net17),
    .Y(_05118_));
 sky130_fd_sc_hd__xnor2_1 _11981_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__o21ai_1 _11982_ (.A1(_05030_),
    .A2(_05034_),
    .B1(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__or3_1 _11983_ (.A(_05030_),
    .B(_05034_),
    .C(_05119_),
    .X(_05121_));
 sky130_fd_sc_hd__and2_1 _11984_ (.A(_05120_),
    .B(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__o22a_1 _11985_ (.A1(net16),
    .A2(net22),
    .B1(net14),
    .B2(net54),
    .X(_05123_));
 sky130_fd_sc_hd__xnor2_1 _11986_ (.A(net69),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__o22a_1 _11987_ (.A1(net67),
    .A2(net9),
    .B1(net4),
    .B2(net65),
    .X(_05125_));
 sky130_fd_sc_hd__xnor2_1 _11988_ (.A(net18),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__a22o_1 _11989_ (.A1(net40),
    .A2(_00690_),
    .B1(_01954_),
    .B2(net42),
    .X(_05128_));
 sky130_fd_sc_hd__xnor2_1 _11990_ (.A(net92),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(_05126_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__and2_1 _11992_ (.A(_05126_),
    .B(_05129_),
    .X(_05131_));
 sky130_fd_sc_hd__or2_1 _11993_ (.A(_05130_),
    .B(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(_05124_),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__and2_1 _11995_ (.A(_05124_),
    .B(_05132_),
    .X(_05134_));
 sky130_fd_sc_hd__nor2_1 _11996_ (.A(_05133_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_1 _11997_ (.A1(_05049_),
    .A2(_05053_),
    .B1(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__or3_1 _11998_ (.A(_05049_),
    .B(_05053_),
    .C(_05135_),
    .X(_05137_));
 sky130_fd_sc_hd__nand2_1 _11999_ (.A(_05136_),
    .B(_05137_),
    .Y(_05139_));
 sky130_fd_sc_hd__a21o_1 _12000_ (.A1(_05037_),
    .A2(_05041_),
    .B1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nand3_1 _12001_ (.A(_05037_),
    .B(_05041_),
    .C(_05139_),
    .Y(_05141_));
 sky130_fd_sc_hd__and2_1 _12002_ (.A(_05140_),
    .B(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__nand2_1 _12003_ (.A(_05122_),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__or2_1 _12004_ (.A(_05122_),
    .B(_05142_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(_05143_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__a21o_1 _12006_ (.A1(_05055_),
    .A2(_05058_),
    .B1(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__nand3_1 _12007_ (.A(_05055_),
    .B(_05058_),
    .C(_05145_),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__a21oi_1 _12009_ (.A1(_05060_),
    .A2(_05063_),
    .B1(_05148_),
    .Y(_05150_));
 sky130_fd_sc_hd__inv_2 _12010_ (.A(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__and3_1 _12011_ (.A(_05060_),
    .B(_05063_),
    .C(_05148_),
    .X(_05152_));
 sky130_fd_sc_hd__or2_2 _12012_ (.A(_05150_),
    .B(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__a21o_1 _12013_ (.A1(_04976_),
    .A2(_05066_),
    .B1(_05067_),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_1 _12014_ (.A(_04979_),
    .B(_05069_),
    .Y(_05155_));
 sky130_fd_sc_hd__a21bo_1 _12015_ (.A1(_04980_),
    .A2(_05155_),
    .B1_N(_05154_),
    .X(_05156_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(_04981_),
    .B(_05155_),
    .Y(_05157_));
 sky130_fd_sc_hd__o21bai_2 _12017_ (.A1(_04800_),
    .A2(_05157_),
    .B1_N(_05156_),
    .Y(_05158_));
 sky130_fd_sc_hd__xnor2_2 _12018_ (.A(_05153_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__inv_2 _12019_ (.A(_05159_),
    .Y(_05161_));
 sky130_fd_sc_hd__and4_2 _12020_ (.A(_04930_),
    .B(_04932_),
    .C(_04988_),
    .D(_05076_),
    .X(_05162_));
 sky130_fd_sc_hd__nor2_1 _12021_ (.A(net158),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__o31a_1 _12022_ (.A1(net158),
    .A2(_05161_),
    .A3(_05162_),
    .B1(_02245_),
    .X(_05164_));
 sky130_fd_sc_hd__o21a_1 _12023_ (.A1(_05159_),
    .A2(_05163_),
    .B1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__a21oi_1 _12024_ (.A1(_05442_),
    .A2(_05085_),
    .B1(_05420_),
    .Y(_05166_));
 sky130_fd_sc_hd__mux2_1 _12025_ (.A0(_06388_),
    .A1(_05166_),
    .S(net285),
    .X(_05167_));
 sky130_fd_sc_hd__a21oi_1 _12026_ (.A1(_05225_),
    .A2(_05167_),
    .B1(_02324_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21a_1 _12027_ (.A1(_05225_),
    .A2(_05167_),
    .B1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__a21o_1 _12028_ (.A1(net161),
    .A2(_01880_),
    .B1(_01887_),
    .X(_05170_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(net233),
    .B(_05170_),
    .Y(_05172_));
 sky130_fd_sc_hd__a31oi_4 _12030_ (.A1(net161),
    .A2(_01880_),
    .A3(_01887_),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21oi_1 _12031_ (.A1(_05090_),
    .A2(_05092_),
    .B1(_05089_),
    .Y(_05174_));
 sky130_fd_sc_hd__nor2_1 _12032_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05176_));
 sky130_fd_sc_hd__and2b_1 _12034_ (.A_N(_05175_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__xnor2_1 _12035_ (.A(_05174_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(_03372_),
    .A1(_05178_),
    .S(net251),
    .X(_05179_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(\div_res[23] ),
    .B(_05097_),
    .X(_05180_));
 sky130_fd_sc_hd__a21oi_1 _12038_ (.A1(net164),
    .A2(_05180_),
    .B1(\div_res[24] ),
    .Y(_05181_));
 sky130_fd_sc_hd__a311o_1 _12039_ (.A1(\div_res[24] ),
    .A2(net164),
    .A3(_05180_),
    .B1(_05181_),
    .C1(net184),
    .X(_05183_));
 sky130_fd_sc_hd__or2_1 _12040_ (.A(\div_shifter[55] ),
    .B(_05100_),
    .X(_05184_));
 sky130_fd_sc_hd__a21oi_1 _12041_ (.A1(net227),
    .A2(_05184_),
    .B1(\div_shifter[56] ),
    .Y(_05185_));
 sky130_fd_sc_hd__a31o_1 _12042_ (.A1(\div_shifter[56] ),
    .A2(net227),
    .A3(_05184_),
    .B1(net231),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_1 _12043_ (.A0(_02331_),
    .A1(_02325_),
    .S(_05203_),
    .X(_05187_));
 sky130_fd_sc_hd__o21a_1 _12044_ (.A1(_02321_),
    .A2(_05187_),
    .B1(_05214_),
    .X(_05188_));
 sky130_fd_sc_hd__a221o_1 _12045_ (.A1(_05193_),
    .A2(net242),
    .B1(_02319_),
    .B2(_03372_),
    .C1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__a21oi_1 _12046_ (.A1(net170),
    .A2(_03378_),
    .B1(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__o211ai_1 _12047_ (.A1(_05185_),
    .A2(_05186_),
    .B1(_05190_),
    .C1(_05183_),
    .Y(_05191_));
 sky130_fd_sc_hd__a211o_1 _12048_ (.A1(net197),
    .A2(_05179_),
    .B1(_05191_),
    .C1(_05173_),
    .X(_05192_));
 sky130_fd_sc_hd__o31a_1 _12049_ (.A1(_05165_),
    .A2(_05169_),
    .A3(_05192_),
    .B1(net247),
    .X(_05194_));
 sky130_fd_sc_hd__or2_1 _12050_ (.A(curr_PC[24]),
    .B(_05112_),
    .X(_05195_));
 sky130_fd_sc_hd__and3_1 _12051_ (.A(curr_PC[23]),
    .B(curr_PC[24]),
    .C(_05023_),
    .X(_05196_));
 sky130_fd_sc_hd__inv_2 _12052_ (.A(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a31o_4 _12053_ (.A1(net248),
    .A2(_05195_),
    .A3(_05197_),
    .B1(_05194_),
    .X(dest_val[24]));
 sky130_fd_sc_hd__o22a_1 _12054_ (.A1(net54),
    .A2(net9),
    .B1(net4),
    .B2(net67),
    .X(_05198_));
 sky130_fd_sc_hd__xnor2_1 _12055_ (.A(net17),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2b_1 _12056_ (.A_N(_05199_),
    .B(_05117_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2b_1 _12057_ (.A_N(_05117_),
    .B(_05199_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _12058_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__nor2_1 _12059_ (.A(net65),
    .B(net17),
    .Y(_05204_));
 sky130_fd_sc_hd__xnor2_1 _12060_ (.A(_05202_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__o31ai_2 _12061_ (.A1(net59),
    .A2(net17),
    .A3(_05117_),
    .B1(_05120_),
    .Y(_05206_));
 sky130_fd_sc_hd__o22a_1 _12062_ (.A1(net16),
    .A2(net14),
    .B1(_00689_),
    .B2(net22),
    .X(_05207_));
 sky130_fd_sc_hd__xnor2_1 _12063_ (.A(net68),
    .B(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(net89),
    .B(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__nand2_1 _12065_ (.A(net89),
    .B(_05208_),
    .Y(_05210_));
 sky130_fd_sc_hd__and2_1 _12066_ (.A(_05209_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__a22o_1 _12067_ (.A1(net40),
    .A2(_01954_),
    .B1(net8),
    .B2(net42),
    .X(_05212_));
 sky130_fd_sc_hd__xor2_1 _12068_ (.A(net92),
    .B(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__nand2_1 _12069_ (.A(_05211_),
    .B(_05213_),
    .Y(_05215_));
 sky130_fd_sc_hd__or2_1 _12070_ (.A(_05211_),
    .B(_05213_),
    .X(_05216_));
 sky130_fd_sc_hd__and2_1 _12071_ (.A(_05215_),
    .B(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__o21a_1 _12072_ (.A1(_05130_),
    .A2(_05133_),
    .B1(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__nor3_1 _12073_ (.A(_05130_),
    .B(_05133_),
    .C(_05217_),
    .Y(_05219_));
 sky130_fd_sc_hd__nor2_1 _12074_ (.A(_05218_),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__xor2_1 _12075_ (.A(_05206_),
    .B(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_05205_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(_05205_),
    .B(_05221_),
    .X(_05223_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_05222_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21o_1 _12079_ (.A1(_05136_),
    .A2(_05140_),
    .B1(_05224_),
    .X(_05226_));
 sky130_fd_sc_hd__nand3_1 _12080_ (.A(_05136_),
    .B(_05140_),
    .C(_05224_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__a21oi_2 _12082_ (.A1(_05143_),
    .A2(_05146_),
    .B1(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand3_1 _12083_ (.A(_05143_),
    .B(_05146_),
    .C(_05228_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand2b_2 _12084_ (.A_N(_05229_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nor2_1 _12085_ (.A(_05069_),
    .B(_05153_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_05071_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__nor2_1 _12087_ (.A(_04887_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__nor2_1 _12088_ (.A(_04891_),
    .B(_05233_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21oi_1 _12089_ (.A1(_05066_),
    .A2(_05151_),
    .B1(_05152_),
    .Y(_05237_));
 sky130_fd_sc_hd__a21o_1 _12090_ (.A1(_05070_),
    .A2(_05232_),
    .B1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a211o_1 _12091_ (.A1(_04515_),
    .A2(_05234_),
    .B1(_05235_),
    .C1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__xnor2_2 _12092_ (.A(_05231_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__a21oi_1 _12093_ (.A1(_05161_),
    .A2(_05162_),
    .B1(net158),
    .Y(_05241_));
 sky130_fd_sc_hd__nor2_1 _12094_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__a21o_1 _12095_ (.A1(_05240_),
    .A2(_05241_),
    .B1(_02246_),
    .X(_05243_));
 sky130_fd_sc_hd__o21a_1 _12096_ (.A1(_05225_),
    .A2(_05166_),
    .B1(_05203_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(_06406_),
    .A1(_05244_),
    .S(net286),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_1 _12098_ (.A(_05149_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21o_1 _12099_ (.A1(_05149_),
    .A2(_05245_),
    .B1(net236),
    .X(_05248_));
 sky130_fd_sc_hd__a21oi_1 _12100_ (.A1(net162),
    .A2(_01888_),
    .B1(_01802_),
    .Y(_05249_));
 sky130_fd_sc_hd__a31o_1 _12101_ (.A1(net162),
    .A2(_01802_),
    .A3(_01888_),
    .B1(_02330_),
    .X(_05250_));
 sky130_fd_sc_hd__o21a_1 _12102_ (.A1(_05174_),
    .A2(_05175_),
    .B1(_05176_),
    .X(_05251_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05253_));
 sky130_fd_sc_hd__and2b_1 _12105_ (.A_N(_05252_),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__xnor2_1 _12106_ (.A(_05251_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__o21a_1 _12107_ (.A1(net250),
    .A2(_03237_),
    .B1(net197),
    .X(_05256_));
 sky130_fd_sc_hd__o21ai_1 _12108_ (.A1(net224),
    .A2(_05255_),
    .B1(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__or2_1 _12109_ (.A(\div_shifter[56] ),
    .B(_05184_),
    .X(_05259_));
 sky130_fd_sc_hd__a21oi_1 _12110_ (.A1(net227),
    .A2(_05259_),
    .B1(\div_shifter[57] ),
    .Y(_05260_));
 sky130_fd_sc_hd__a311o_1 _12111_ (.A1(\div_shifter[57] ),
    .A2(net227),
    .A3(_05259_),
    .B1(_05260_),
    .C1(net231),
    .X(_05261_));
 sky130_fd_sc_hd__or2_1 _12112_ (.A(\div_res[24] ),
    .B(_05180_),
    .X(_05262_));
 sky130_fd_sc_hd__a21oi_1 _12113_ (.A1(net164),
    .A2(_05262_),
    .B1(\div_res[25] ),
    .Y(_05263_));
 sky130_fd_sc_hd__a311o_1 _12114_ (.A1(\div_res[25] ),
    .A2(net164),
    .A3(_05262_),
    .B1(_05263_),
    .C1(net184),
    .X(_05264_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(net235),
    .A1(_02332_),
    .S(_05127_),
    .X(_05265_));
 sky130_fd_sc_hd__a21o_1 _12116_ (.A1(_02322_),
    .A2(_05265_),
    .B1(_05138_),
    .X(_05266_));
 sky130_fd_sc_hd__o21ai_1 _12117_ (.A1(_05116_),
    .A2(_06461_),
    .B1(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__a221o_1 _12118_ (.A1(_02319_),
    .A2(_03237_),
    .B1(_03243_),
    .B2(net170),
    .C1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__and3b_1 _12119_ (.A_N(_05268_),
    .B(_05264_),
    .C(_05261_),
    .X(_05270_));
 sky130_fd_sc_hd__o211a_1 _12120_ (.A1(_05249_),
    .A2(_05250_),
    .B1(_05257_),
    .C1(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__o221a_1 _12121_ (.A1(_05242_),
    .A2(_05243_),
    .B1(_05246_),
    .B2(_05248_),
    .C1(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__nor2_1 _12122_ (.A(curr_PC[25]),
    .B(_05196_),
    .Y(_05273_));
 sky130_fd_sc_hd__and2_1 _12123_ (.A(curr_PC[25]),
    .B(_05196_),
    .X(_05274_));
 sky130_fd_sc_hd__or3_1 _12124_ (.A(net245),
    .B(_05273_),
    .C(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__o21ai_4 _12125_ (.A1(net249),
    .A2(_05272_),
    .B1(_05275_),
    .Y(dest_val[25]));
 sky130_fd_sc_hd__nor2_1 _12126_ (.A(_05159_),
    .B(_05240_),
    .Y(_05276_));
 sky130_fd_sc_hd__a21o_1 _12127_ (.A1(_05162_),
    .A2(_05276_),
    .B1(net158),
    .X(_05277_));
 sky130_fd_sc_hd__a21o_1 _12128_ (.A1(_05206_),
    .A2(_05220_),
    .B1(_05218_),
    .X(_05278_));
 sky130_fd_sc_hd__a21bo_1 _12129_ (.A1(_05201_),
    .A2(_05204_),
    .B1_N(_05200_),
    .X(_05280_));
 sky130_fd_sc_hd__o22a_1 _12130_ (.A1(net14),
    .A2(_00689_),
    .B1(net12),
    .B2(net22),
    .X(_05281_));
 sky130_fd_sc_hd__xnor2_1 _12131_ (.A(net69),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(_00233_),
    .B(net8),
    .Y(_05283_));
 sky130_fd_sc_hd__a22o_1 _12133_ (.A1(_00235_),
    .A2(net8),
    .B1(_05283_),
    .B2(net93),
    .X(_05284_));
 sky130_fd_sc_hd__and2b_1 _12134_ (.A_N(_05284_),
    .B(_05282_),
    .X(_05285_));
 sky130_fd_sc_hd__and2b_1 _12135_ (.A_N(_05282_),
    .B(_05284_),
    .X(_05286_));
 sky130_fd_sc_hd__nor2_1 _12136_ (.A(_05285_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__a21oi_1 _12137_ (.A1(_05209_),
    .A2(_05215_),
    .B1(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__and3_1 _12138_ (.A(_05209_),
    .B(_05215_),
    .C(_05287_),
    .X(_05289_));
 sky130_fd_sc_hd__nor2_1 _12139_ (.A(_05288_),
    .B(_05289_),
    .Y(_05291_));
 sky130_fd_sc_hd__and2_1 _12140_ (.A(_05280_),
    .B(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__xnor2_1 _12141_ (.A(_05280_),
    .B(_05291_),
    .Y(_05293_));
 sky130_fd_sc_hd__a22o_1 _12142_ (.A1(_00398_),
    .A2(_01970_),
    .B1(_02085_),
    .B2(_06553_),
    .X(_05294_));
 sky130_fd_sc_hd__nor2_1 _12143_ (.A(_06492_),
    .B(net17),
    .Y(_05295_));
 sky130_fd_sc_hd__xnor2_1 _12144_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__nor2_1 _12145_ (.A(_05293_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__and2_1 _12146_ (.A(_05293_),
    .B(_05296_),
    .X(_05298_));
 sky130_fd_sc_hd__or2_1 _12147_ (.A(_05297_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__and2b_1 _12148_ (.A_N(_05299_),
    .B(_05278_),
    .X(_05300_));
 sky130_fd_sc_hd__xor2_1 _12149_ (.A(_05278_),
    .B(_05299_),
    .X(_05302_));
 sky130_fd_sc_hd__a21oi_2 _12150_ (.A1(_05222_),
    .A2(_05226_),
    .B1(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__and3_1 _12151_ (.A(_05222_),
    .B(_05226_),
    .C(_05302_),
    .X(_05304_));
 sky130_fd_sc_hd__nor2_2 _12152_ (.A(_05303_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21ai_1 _12153_ (.A1(_05150_),
    .A2(_05229_),
    .B1(_05230_),
    .Y(_05306_));
 sky130_fd_sc_hd__or2_1 _12154_ (.A(_05153_),
    .B(_05231_),
    .X(_05307_));
 sky130_fd_sc_hd__o21a_1 _12155_ (.A1(_05154_),
    .A2(_05307_),
    .B1(_05306_),
    .X(_05308_));
 sky130_fd_sc_hd__o41a_1 _12156_ (.A1(_04979_),
    .A2(_04987_),
    .A3(_05069_),
    .A4(_05307_),
    .B1(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__xor2_2 _12157_ (.A(_05305_),
    .B(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__nor2_1 _12158_ (.A(_05277_),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__a21o_1 _12159_ (.A1(_05277_),
    .A2(_05310_),
    .B1(_02246_),
    .X(_05313_));
 sky130_fd_sc_hd__o21ba_1 _12160_ (.A1(_05149_),
    .A2(_05244_),
    .B1_N(_05127_),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(_06407_),
    .A1(_05314_),
    .S(net286),
    .X(_05315_));
 sky130_fd_sc_hd__nor2_1 _12162_ (.A(_05355_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__a211o_1 _12163_ (.A1(_05355_),
    .A2(_05315_),
    .B1(_05316_),
    .C1(net236),
    .X(_05317_));
 sky130_fd_sc_hd__o21a_1 _12164_ (.A1(net156),
    .A2(_01889_),
    .B1(_01894_),
    .X(_05318_));
 sky130_fd_sc_hd__o31ai_2 _12165_ (.A1(net156),
    .A2(_01889_),
    .A3(_01894_),
    .B1(net233),
    .Y(_05319_));
 sky130_fd_sc_hd__o21a_1 _12166_ (.A1(_05251_),
    .A2(_05252_),
    .B1(_05253_),
    .X(_05320_));
 sky130_fd_sc_hd__nor2_1 _12167_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2_1 _12168_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2b_1 _12169_ (.A_N(_05321_),
    .B(_05322_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_1 _12170_ (.A(_05320_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nor2_1 _12171_ (.A(net250),
    .B(_03102_),
    .Y(_05326_));
 sky130_fd_sc_hd__a211o_1 _12172_ (.A1(net250),
    .A2(_05325_),
    .B1(_05326_),
    .C1(_06449_),
    .X(_05327_));
 sky130_fd_sc_hd__or2_1 _12173_ (.A(\div_shifter[57] ),
    .B(_05259_),
    .X(_05328_));
 sky130_fd_sc_hd__a21oi_1 _12174_ (.A1(net227),
    .A2(_05328_),
    .B1(\div_shifter[58] ),
    .Y(_05329_));
 sky130_fd_sc_hd__a311o_1 _12175_ (.A1(\div_shifter[58] ),
    .A2(net227),
    .A3(_05328_),
    .B1(_05329_),
    .C1(net231),
    .X(_05330_));
 sky130_fd_sc_hd__or2_1 _12176_ (.A(\div_res[25] ),
    .B(_05262_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _12177_ (.A1(net166),
    .A2(_05331_),
    .B1(\div_res[26] ),
    .Y(_05332_));
 sky130_fd_sc_hd__a311o_1 _12178_ (.A1(\div_res[26] ),
    .A2(net164),
    .A3(_05331_),
    .B1(_05332_),
    .C1(net184),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(net235),
    .A1(_02332_),
    .S(_05323_),
    .X(_05335_));
 sky130_fd_sc_hd__a21o_1 _12180_ (.A1(_02322_),
    .A2(_05335_),
    .B1(_05344_),
    .X(_05336_));
 sky130_fd_sc_hd__o21ai_1 _12181_ (.A1(_05312_),
    .A2(net241),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__a221o_1 _12182_ (.A1(_02319_),
    .A2(_03102_),
    .B1(_03108_),
    .B2(net170),
    .C1(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__and4b_1 _12183_ (.A_N(_05338_),
    .B(_05333_),
    .C(_05330_),
    .D(_05327_),
    .X(_05339_));
 sky130_fd_sc_hd__o211a_1 _12184_ (.A1(_05318_),
    .A2(_05319_),
    .B1(_05339_),
    .C1(_05317_),
    .X(_05340_));
 sky130_fd_sc_hd__o21ai_1 _12185_ (.A1(_05311_),
    .A2(_05313_),
    .B1(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__and3_1 _12186_ (.A(curr_PC[25]),
    .B(curr_PC[26]),
    .C(_05196_),
    .X(_05342_));
 sky130_fd_sc_hd__o21ai_1 _12187_ (.A1(curr_PC[26]),
    .A2(_05274_),
    .B1(net249),
    .Y(_05343_));
 sky130_fd_sc_hd__a2bb2o_4 _12188_ (.A1_N(_05342_),
    .A2_N(_05343_),
    .B1(net247),
    .B2(_05341_),
    .X(dest_val[26]));
 sky130_fd_sc_hd__xor2_1 _12189_ (.A(curr_PC[27]),
    .B(_05342_),
    .X(_05345_));
 sky130_fd_sc_hd__o22a_1 _12190_ (.A1(_00689_),
    .A2(net9),
    .B1(net4),
    .B2(_00399_),
    .X(_05346_));
 sky130_fd_sc_hd__xnor2_1 _12191_ (.A(net17),
    .B(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__or2_1 _12192_ (.A(net93),
    .B(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(net93),
    .B(_05347_),
    .Y(_05349_));
 sky130_fd_sc_hd__and2_1 _12194_ (.A(_05348_),
    .B(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__o22a_1 _12195_ (.A1(net14),
    .A2(net12),
    .B1(net6),
    .B2(net22),
    .X(_05351_));
 sky130_fd_sc_hd__xnor2_1 _12196_ (.A(net68),
    .B(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__inv_2 _12197_ (.A(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_05350_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__or2_1 _12199_ (.A(_05350_),
    .B(_05353_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _12200_ (.A(_05354_),
    .B(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__o21a_1 _12201_ (.A1(net66),
    .A2(_05294_),
    .B1(net54),
    .X(_05358_));
 sky130_fd_sc_hd__or4_1 _12202_ (.A(net66),
    .B(net54),
    .C(net17),
    .D(_05294_),
    .X(_05359_));
 sky130_fd_sc_hd__or3b_1 _12203_ (.A(net17),
    .B(_05358_),
    .C_N(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__xor2_1 _12204_ (.A(_05285_),
    .B(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__and3_1 _12205_ (.A(_05354_),
    .B(_05356_),
    .C(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__xnor2_1 _12206_ (.A(_05357_),
    .B(_05361_),
    .Y(_05363_));
 sky130_fd_sc_hd__o21a_1 _12207_ (.A1(_05288_),
    .A2(_05292_),
    .B1(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__nor3_1 _12208_ (.A(_05288_),
    .B(_05292_),
    .C(_05363_),
    .Y(_05365_));
 sky130_fd_sc_hd__nor2_1 _12209_ (.A(_05364_),
    .B(_05365_),
    .Y(_05367_));
 sky130_fd_sc_hd__o21ai_2 _12210_ (.A1(_05297_),
    .A2(_05300_),
    .B1(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__inv_2 _12211_ (.A(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__or3_1 _12212_ (.A(_05297_),
    .B(_05300_),
    .C(_05367_),
    .X(_05370_));
 sky130_fd_sc_hd__and2_1 _12213_ (.A(_05368_),
    .B(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__and2b_1 _12214_ (.A_N(_05231_),
    .B(_05305_),
    .X(_05372_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05232_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__o21ba_1 _12216_ (.A1(_05229_),
    .A2(_05303_),
    .B1_N(_05304_),
    .X(_05374_));
 sky130_fd_sc_hd__inv_2 _12217_ (.A(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__a21oi_1 _12218_ (.A1(_05237_),
    .A2(_05372_),
    .B1(_05374_),
    .Y(_05376_));
 sky130_fd_sc_hd__o21ai_2 _12219_ (.A1(_05075_),
    .A2(_05373_),
    .B1(_05376_),
    .Y(_05378_));
 sky130_fd_sc_hd__xnor2_2 _12220_ (.A(_05371_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__a31o_1 _12221_ (.A1(_05162_),
    .A2(_05276_),
    .A3(_05310_),
    .B1(net158),
    .X(_05380_));
 sky130_fd_sc_hd__a21oi_1 _12222_ (.A1(_05379_),
    .A2(_05380_),
    .B1(_02246_),
    .Y(_05381_));
 sky130_fd_sc_hd__o21a_1 _12223_ (.A1(_05379_),
    .A2(_05380_),
    .B1(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__o211a_1 _12224_ (.A1(_05355_),
    .A2(_05314_),
    .B1(net286),
    .C1(_05334_),
    .X(_05383_));
 sky130_fd_sc_hd__a21o_1 _12225_ (.A1(net294),
    .A2(_06408_),
    .B1(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__a21oi_1 _12226_ (.A1(_05073_),
    .A2(_05384_),
    .B1(net236),
    .Y(_05385_));
 sky130_fd_sc_hd__o21a_1 _12227_ (.A1(_05073_),
    .A2(_05384_),
    .B1(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__a21bo_1 _12228_ (.A1(net161),
    .A2(_01895_),
    .B1_N(_01896_),
    .X(_05387_));
 sky130_fd_sc_hd__or3b_1 _12229_ (.A(net158),
    .B(_01896_),
    .C_N(_01895_),
    .X(_05389_));
 sky130_fd_sc_hd__o21a_1 _12230_ (.A1(_05320_),
    .A2(_05321_),
    .B1(_05322_),
    .X(_05390_));
 sky130_fd_sc_hd__nor2_1 _12231_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _12232_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05392_));
 sky130_fd_sc_hd__and2b_1 _12233_ (.A_N(_05391_),
    .B(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12234_ (.A(_05390_),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(_02968_),
    .A1(_05394_),
    .S(net251),
    .X(_05395_));
 sky130_fd_sc_hd__or2_1 _12236_ (.A(\div_res[26] ),
    .B(_05331_),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _12237_ (.A1(net166),
    .A2(_05396_),
    .B1(\div_res[27] ),
    .X(_05397_));
 sky130_fd_sc_hd__nand3_1 _12238_ (.A(\div_res[27] ),
    .B(net166),
    .C(_05396_),
    .Y(_05398_));
 sky130_fd_sc_hd__or2_1 _12239_ (.A(\div_shifter[58] ),
    .B(_05328_),
    .X(_05400_));
 sky130_fd_sc_hd__a21oi_1 _12240_ (.A1(net229),
    .A2(_05400_),
    .B1(\div_shifter[59] ),
    .Y(_05401_));
 sky130_fd_sc_hd__a31o_1 _12241_ (.A1(\div_shifter[59] ),
    .A2(net229),
    .A3(_05400_),
    .B1(net232),
    .X(_05402_));
 sky130_fd_sc_hd__nor2_1 _12242_ (.A(_05401_),
    .B(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a21oi_1 _12243_ (.A1(_05062_),
    .A2(_02325_),
    .B1(_02321_),
    .Y(_05404_));
 sky130_fd_sc_hd__o221a_1 _12244_ (.A1(_05040_),
    .A2(net241),
    .B1(_02332_),
    .B2(_05062_),
    .C1(net247),
    .X(_05405_));
 sky130_fd_sc_hd__o21ai_1 _12245_ (.A1(_05051_),
    .A2(_05404_),
    .B1(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__a221o_1 _12246_ (.A1(_02319_),
    .A2(_02968_),
    .B1(_02974_),
    .B2(net170),
    .C1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__a31o_1 _12247_ (.A1(_02334_),
    .A2(_05397_),
    .A3(_05398_),
    .B1(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__a211o_1 _12248_ (.A1(_06448_),
    .A2(_05395_),
    .B1(_05403_),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a31o_1 _12249_ (.A1(net233),
    .A2(_05387_),
    .A3(_05389_),
    .B1(_05409_),
    .X(_05411_));
 sky130_fd_sc_hd__o32a_4 _12250_ (.A1(_05382_),
    .A2(_05386_),
    .A3(_05411_),
    .B1(_05345_),
    .B2(net247),
    .X(dest_val[27]));
 sky130_fd_sc_hd__o31a_1 _12251_ (.A1(net17),
    .A2(_05285_),
    .A3(_05358_),
    .B1(_05359_),
    .X(_05412_));
 sky130_fd_sc_hd__o22a_1 _12252_ (.A1(net12),
    .A2(net9),
    .B1(net4),
    .B2(_00689_),
    .X(_05413_));
 sky130_fd_sc_hd__xnor2_1 _12253_ (.A(net17),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__a21oi_1 _12254_ (.A1(_05348_),
    .A2(_05354_),
    .B1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__and3_1 _12255_ (.A(_05348_),
    .B(_05354_),
    .C(_05414_),
    .X(_05416_));
 sky130_fd_sc_hd__nor2_1 _12256_ (.A(_05415_),
    .B(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__nor2_1 _12257_ (.A(net16),
    .B(net17),
    .Y(_05418_));
 sky130_fd_sc_hd__xnor2_1 _12258_ (.A(_05417_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__o21a_1 _12259_ (.A1(net14),
    .A2(net6),
    .B1(_00668_),
    .X(_05421_));
 sky130_fd_sc_hd__a31o_1 _12260_ (.A1(net69),
    .A2(_00676_),
    .A3(net8),
    .B1(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__nor2_1 _12261_ (.A(_05419_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__and2_1 _12262_ (.A(_05419_),
    .B(_05422_),
    .X(_05424_));
 sky130_fd_sc_hd__nor3_1 _12263_ (.A(_05412_),
    .B(_05423_),
    .C(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__o21a_1 _12264_ (.A1(_05423_),
    .A2(_05424_),
    .B1(_05412_),
    .X(_05426_));
 sky130_fd_sc_hd__nor2_1 _12265_ (.A(_05425_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__o21ai_2 _12266_ (.A1(_05362_),
    .A2(_05364_),
    .B1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nor3_1 _12267_ (.A(_05362_),
    .B(_05364_),
    .C(_05427_),
    .Y(_05429_));
 sky130_fd_sc_hd__inv_2 _12268_ (.A(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_05428_),
    .B(_05430_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_1 _12270_ (.A(_05305_),
    .B(_05371_),
    .Y(_05433_));
 sky130_fd_sc_hd__or3_1 _12271_ (.A(_05157_),
    .B(_05307_),
    .C(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__o21ai_1 _12272_ (.A1(_05303_),
    .A2(_05369_),
    .B1(_05370_),
    .Y(_05435_));
 sky130_fd_sc_hd__nand2b_1 _12273_ (.A_N(_05307_),
    .B(_05156_),
    .Y(_05436_));
 sky130_fd_sc_hd__a21o_1 _12274_ (.A1(_05306_),
    .A2(_05436_),
    .B1(_05433_),
    .X(_05437_));
 sky130_fd_sc_hd__o211a_1 _12275_ (.A1(_04800_),
    .A2(_05434_),
    .B1(_05435_),
    .C1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__xnor2_2 _12276_ (.A(_05432_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__inv_2 _12277_ (.A(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__or4bb_1 _12278_ (.A(_05159_),
    .B(_05240_),
    .C_N(_05310_),
    .D_N(_05379_),
    .X(_05441_));
 sky130_fd_sc_hd__and4_1 _12279_ (.A(_05162_),
    .B(_05276_),
    .C(_05310_),
    .D(_05379_),
    .X(_05443_));
 sky130_fd_sc_hd__or3_1 _12280_ (.A(net158),
    .B(_05439_),
    .C(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__o21ai_1 _12281_ (.A1(net158),
    .A2(_05443_),
    .B1(_05439_),
    .Y(_05445_));
 sky130_fd_sc_hd__a21o_1 _12282_ (.A1(_05062_),
    .A2(_05334_),
    .B1(_05051_),
    .X(_05446_));
 sky130_fd_sc_hd__o31ai_1 _12283_ (.A1(_05073_),
    .A2(_05355_),
    .A3(_05314_),
    .B1(_05446_),
    .Y(_05447_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(_06409_),
    .A1(_05447_),
    .S(net286),
    .X(_05448_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(_04931_),
    .B(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__o211a_1 _12286_ (.A1(_04931_),
    .A2(_05448_),
    .B1(_05449_),
    .C1(_02323_),
    .X(_05450_));
 sky130_fd_sc_hd__o21ai_1 _12287_ (.A1(net158),
    .A2(_01897_),
    .B1(_01904_),
    .Y(_05451_));
 sky130_fd_sc_hd__o311a_1 _12288_ (.A1(net156),
    .A2(_01897_),
    .A3(_01904_),
    .B1(_02329_),
    .C1(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__o21ai_2 _12289_ (.A1(_05390_),
    .A2(_05391_),
    .B1(_05392_),
    .Y(_05454_));
 sky130_fd_sc_hd__xor2_1 _12290_ (.A(reg1_val[28]),
    .B(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__or2_1 _12291_ (.A(net251),
    .B(_02832_),
    .X(_05456_));
 sky130_fd_sc_hd__o211a_1 _12292_ (.A1(net224),
    .A2(_05455_),
    .B1(_05456_),
    .C1(_06448_),
    .X(_05457_));
 sky130_fd_sc_hd__or2_1 _12293_ (.A(\div_res[27] ),
    .B(_05396_),
    .X(_05458_));
 sky130_fd_sc_hd__a21oi_1 _12294_ (.A1(net166),
    .A2(_05458_),
    .B1(\div_res[28] ),
    .Y(_05459_));
 sky130_fd_sc_hd__a31o_1 _12295_ (.A1(\div_res[28] ),
    .A2(net166),
    .A3(_05458_),
    .B1(net183),
    .X(_05460_));
 sky130_fd_sc_hd__or2_1 _12296_ (.A(\div_shifter[59] ),
    .B(_05400_),
    .X(_05461_));
 sky130_fd_sc_hd__a21oi_1 _12297_ (.A1(net229),
    .A2(_05461_),
    .B1(\div_shifter[60] ),
    .Y(_05462_));
 sky130_fd_sc_hd__a31o_1 _12298_ (.A1(\div_shifter[60] ),
    .A2(net229),
    .A3(_05461_),
    .B1(net232),
    .X(_05463_));
 sky130_fd_sc_hd__o21ai_1 _12299_ (.A1(_04910_),
    .A2(net235),
    .B1(_02322_),
    .Y(_05465_));
 sky130_fd_sc_hd__a221o_1 _12300_ (.A1(_04910_),
    .A2(_02331_),
    .B1(_05465_),
    .B2(_04921_),
    .C1(net242),
    .X(_05466_));
 sky130_fd_sc_hd__a221o_1 _12301_ (.A1(net170),
    .A2(_02822_),
    .B1(_02832_),
    .B2(_02319_),
    .C1(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__o21ba_1 _12302_ (.A1(_05462_),
    .A2(_05463_),
    .B1_N(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__o21ai_1 _12303_ (.A1(_05459_),
    .A2(_05460_),
    .B1(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__or4_1 _12304_ (.A(_05450_),
    .B(_05452_),
    .C(_05457_),
    .D(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__a31o_1 _12305_ (.A1(_02245_),
    .A2(_05444_),
    .A3(_05445_),
    .B1(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__o211a_4 _12306_ (.A1(_04899_),
    .A2(_06461_),
    .B1(_05471_),
    .C1(net247),
    .X(dest_val[28]));
 sky130_fd_sc_hd__o22a_1 _12307_ (.A1(net9),
    .A2(net6),
    .B1(net4),
    .B2(net12),
    .X(_05472_));
 sky130_fd_sc_hd__xnor2_1 _12308_ (.A(net17),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(_00689_),
    .B(net17),
    .Y(_05475_));
 sky130_fd_sc_hd__xnor2_1 _12310_ (.A(net68),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nor2_1 _12311_ (.A(_05473_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__and2_1 _12312_ (.A(_05473_),
    .B(_05476_),
    .X(_05478_));
 sky130_fd_sc_hd__nor2_1 _12313_ (.A(_05477_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _12314_ (.A(_05422_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__or2_1 _12315_ (.A(_05422_),
    .B(_05479_),
    .X(_05481_));
 sky130_fd_sc_hd__nand2_1 _12316_ (.A(_05480_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__a31o_1 _12317_ (.A1(_00398_),
    .A2(_02081_),
    .A3(_05417_),
    .B1(_05415_),
    .X(_05483_));
 sky130_fd_sc_hd__nand2b_1 _12318_ (.A_N(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__xnor2_1 _12319_ (.A(_05482_),
    .B(_05483_),
    .Y(_05486_));
 sky130_fd_sc_hd__nor3_1 _12320_ (.A(_05423_),
    .B(_05425_),
    .C(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__o21ai_2 _12321_ (.A1(_05423_),
    .A2(_05425_),
    .B1(_05486_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2b_1 _12322_ (.A_N(_05487_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__or3b_1 _12323_ (.A(_05369_),
    .B(_05432_),
    .C_N(_05370_),
    .X(_05490_));
 sky130_fd_sc_hd__or4_1 _12324_ (.A(_05231_),
    .B(_05303_),
    .C(_05304_),
    .D(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__nand2b_1 _12325_ (.A_N(_05491_),
    .B(_05238_),
    .Y(_05492_));
 sky130_fd_sc_hd__a21o_1 _12326_ (.A1(_05368_),
    .A2(_05428_),
    .B1(_05429_),
    .X(_05493_));
 sky130_fd_sc_hd__o211a_1 _12327_ (.A1(_05375_),
    .A2(_05490_),
    .B1(_05492_),
    .C1(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__o31a_1 _12328_ (.A1(_04892_),
    .A2(_05233_),
    .A3(_05491_),
    .B1(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__xnor2_1 _12329_ (.A(_05489_),
    .B(_05495_),
    .Y(_05497_));
 sky130_fd_sc_hd__nor3b_1 _12330_ (.A(_05440_),
    .B(_05441_),
    .C_N(_05162_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_1 _12331_ (.A1(net158),
    .A2(_05498_),
    .B1(_05497_),
    .Y(_05499_));
 sky130_fd_sc_hd__o31a_1 _12332_ (.A1(_06465_),
    .A2(_05497_),
    .A3(_05498_),
    .B1(_02245_),
    .X(_05500_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(_05499_),
    .B(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__a21o_1 _12334_ (.A1(_04921_),
    .A2(_05447_),
    .B1(_04910_),
    .X(_05502_));
 sky130_fd_sc_hd__nand2_1 _12335_ (.A(net295),
    .B(_06410_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21a_1 _12336_ (.A1(net295),
    .A2(_05502_),
    .B1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__o21ai_1 _12337_ (.A1(_04844_),
    .A2(_05504_),
    .B1(_02323_),
    .Y(_05505_));
 sky130_fd_sc_hd__a21oi_1 _12338_ (.A1(_04844_),
    .A2(_05504_),
    .B1(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__a21oi_1 _12339_ (.A1(net162),
    .A2(_01905_),
    .B1(_01801_),
    .Y(_05508_));
 sky130_fd_sc_hd__a311oi_2 _12340_ (.A1(net161),
    .A2(_01801_),
    .A3(_01905_),
    .B1(_02330_),
    .C1(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__and3_1 _12341_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05454_),
    .X(_05510_));
 sky130_fd_sc_hd__a21oi_1 _12342_ (.A1(reg1_val[28]),
    .A2(_05454_),
    .B1(reg1_val[29]),
    .Y(_05511_));
 sky130_fd_sc_hd__o21a_1 _12343_ (.A1(_05510_),
    .A2(_05511_),
    .B1(net251),
    .X(_05512_));
 sky130_fd_sc_hd__a211o_1 _12344_ (.A1(net224),
    .A2(_02653_),
    .B1(_05512_),
    .C1(net196),
    .X(_05513_));
 sky130_fd_sc_hd__or2_1 _12345_ (.A(\div_res[28] ),
    .B(_05458_),
    .X(_05514_));
 sky130_fd_sc_hd__a21o_1 _12346_ (.A1(net166),
    .A2(_05514_),
    .B1(\div_res[29] ),
    .X(_05515_));
 sky130_fd_sc_hd__nand3_1 _12347_ (.A(\div_res[29] ),
    .B(net166),
    .C(_05514_),
    .Y(_05516_));
 sky130_fd_sc_hd__or2_1 _12348_ (.A(\div_shifter[60] ),
    .B(_05461_),
    .X(_05517_));
 sky130_fd_sc_hd__and2_1 _12349_ (.A(net229),
    .B(_05517_),
    .X(_05519_));
 sky130_fd_sc_hd__o21ai_1 _12350_ (.A1(\div_shifter[61] ),
    .A2(_05519_),
    .B1(_02336_),
    .Y(_05520_));
 sky130_fd_sc_hd__a21oi_1 _12351_ (.A1(\div_shifter[61] ),
    .A2(_05519_),
    .B1(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_1 _12352_ (.A1(_04823_),
    .A2(net235),
    .B1(net186),
    .Y(_05522_));
 sky130_fd_sc_hd__a221o_1 _12353_ (.A1(_04823_),
    .A2(_02331_),
    .B1(_05522_),
    .B2(_04834_),
    .C1(_06460_),
    .X(_05523_));
 sky130_fd_sc_hd__a221o_1 _12354_ (.A1(_02319_),
    .A2(_02654_),
    .B1(_02669_),
    .B2(net170),
    .C1(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a311o_1 _12355_ (.A1(_02334_),
    .A2(_05515_),
    .A3(_05516_),
    .B1(_05521_),
    .C1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__or4b_1 _12356_ (.A(_05506_),
    .B(_05509_),
    .C(_05525_),
    .D_N(_05513_),
    .X(_05526_));
 sky130_fd_sc_hd__o221a_4 _12357_ (.A1(_04812_),
    .A2(net241),
    .B1(_05501_),
    .B2(_05526_),
    .C1(net247),
    .X(dest_val[29]));
 sky130_fd_sc_hd__a21o_1 _12358_ (.A1(net68),
    .A2(_05475_),
    .B1(_05477_),
    .X(_05527_));
 sky130_fd_sc_hd__o21ai_1 _12359_ (.A1(_01968_),
    .A2(net6),
    .B1(net17),
    .Y(_05529_));
 sky130_fd_sc_hd__or2_1 _12360_ (.A(net6),
    .B(_02083_),
    .X(_05530_));
 sky130_fd_sc_hd__o21ai_1 _12361_ (.A1(_01954_),
    .A2(_05530_),
    .B1(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__a31o_1 _12362_ (.A1(_01954_),
    .A2(_02081_),
    .A3(_05530_),
    .B1(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__nand2_1 _12363_ (.A(_05527_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__or2_1 _12364_ (.A(_05527_),
    .B(_05532_),
    .X(_05534_));
 sky130_fd_sc_hd__nand2_1 _12365_ (.A(_05533_),
    .B(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(_05480_),
    .B(_05484_),
    .C(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__a21oi_1 _12367_ (.A1(_05480_),
    .A2(_05484_),
    .B1(_05535_),
    .Y(_05537_));
 sky130_fd_sc_hd__or2_1 _12368_ (.A(_05536_),
    .B(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__or2_1 _12369_ (.A(_05432_),
    .B(_05489_),
    .X(_05540_));
 sky130_fd_sc_hd__o221a_1 _12370_ (.A1(_05428_),
    .A2(_05487_),
    .B1(_05540_),
    .B2(_05435_),
    .C1(_05488_),
    .X(_05541_));
 sky130_fd_sc_hd__o31a_1 _12371_ (.A1(_05309_),
    .A2(_05433_),
    .A3(_05540_),
    .B1(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__xor2_1 _12372_ (.A(_05538_),
    .B(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__inv_2 _12373_ (.A(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__and4bb_1 _12374_ (.A_N(_05440_),
    .B_N(_05441_),
    .C(_05497_),
    .D(_05162_),
    .X(_05545_));
 sky130_fd_sc_hd__o21ai_1 _12375_ (.A1(net158),
    .A2(_05545_),
    .B1(_05544_),
    .Y(_05546_));
 sky130_fd_sc_hd__o31a_1 _12376_ (.A1(net158),
    .A2(_05544_),
    .A3(_05545_),
    .B1(_02245_),
    .X(_05547_));
 sky130_fd_sc_hd__a21oi_1 _12377_ (.A1(_04834_),
    .A2(_05502_),
    .B1(_04823_),
    .Y(_05548_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(_06411_),
    .A1(_05548_),
    .S(net286),
    .X(_05549_));
 sky130_fd_sc_hd__or2_1 _12379_ (.A(_05008_),
    .B(_05549_),
    .X(_05551_));
 sky130_fd_sc_hd__a21oi_1 _12380_ (.A1(_05008_),
    .A2(_05549_),
    .B1(net236),
    .Y(_05552_));
 sky130_fd_sc_hd__or2_1 _12381_ (.A(_05008_),
    .B(_05548_),
    .X(_05553_));
 sky130_fd_sc_hd__o21a_1 _12382_ (.A1(_01801_),
    .A2(_01905_),
    .B1(net161),
    .X(_05554_));
 sky130_fd_sc_hd__nand2_1 _12383_ (.A(_02018_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21a_1 _12384_ (.A1(_02018_),
    .A2(_05554_),
    .B1(net233),
    .X(_05556_));
 sky130_fd_sc_hd__xnor2_1 _12385_ (.A(reg1_val[30]),
    .B(_05510_),
    .Y(_05557_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(_02530_),
    .A1(_05557_),
    .S(net251),
    .X(_05558_));
 sky130_fd_sc_hd__or2_1 _12387_ (.A(\div_res[29] ),
    .B(_05514_),
    .X(_05559_));
 sky130_fd_sc_hd__a21oi_1 _12388_ (.A1(net166),
    .A2(_05559_),
    .B1(\div_res[30] ),
    .Y(_05560_));
 sky130_fd_sc_hd__a31o_1 _12389_ (.A1(\div_res[30] ),
    .A2(net166),
    .A3(_05559_),
    .B1(net184),
    .X(_05562_));
 sky130_fd_sc_hd__or2_1 _12390_ (.A(_05560_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__or2_1 _12391_ (.A(\div_shifter[61] ),
    .B(_05517_),
    .X(_05564_));
 sky130_fd_sc_hd__a21oi_1 _12392_ (.A1(net229),
    .A2(_05564_),
    .B1(\div_shifter[62] ),
    .Y(_05565_));
 sky130_fd_sc_hd__a31o_1 _12393_ (.A1(\div_shifter[62] ),
    .A2(net229),
    .A3(_05564_),
    .B1(net232),
    .X(_05566_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(net235),
    .A1(net185),
    .S(_04986_),
    .X(_05567_));
 sky130_fd_sc_hd__a21oi_1 _12395_ (.A1(net186),
    .A2(_05567_),
    .B1(_04997_),
    .Y(_05568_));
 sky130_fd_sc_hd__nor2_1 _12396_ (.A(_06460_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__o221a_2 _12397_ (.A1(net168),
    .A2(_02504_),
    .B1(_02530_),
    .B2(_02320_),
    .C1(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__o211a_1 _12398_ (.A1(_05565_),
    .A2(_05566_),
    .B1(_05570_),
    .C1(_05563_),
    .X(_05571_));
 sky130_fd_sc_hd__o21ai_1 _12399_ (.A1(net196),
    .A2(_05558_),
    .B1(_05571_),
    .Y(_05573_));
 sky130_fd_sc_hd__a21o_1 _12400_ (.A1(_05555_),
    .A2(_05556_),
    .B1(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__a221o_1 _12401_ (.A1(_05546_),
    .A2(_05547_),
    .B1(_05551_),
    .B2(_05552_),
    .C1(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__o211a_4 _12402_ (.A1(_04975_),
    .A2(net241),
    .B1(_05575_),
    .C1(net245),
    .X(dest_val[30]));
 sky130_fd_sc_hd__a21o_1 _12403_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_06465_),
    .X(_05576_));
 sky130_fd_sc_hd__nor2_1 _12404_ (.A(_02069_),
    .B(net17),
    .Y(_05577_));
 sky130_fd_sc_hd__or2_1 _12405_ (.A(_05489_),
    .B(_05538_),
    .X(_05578_));
 sky130_fd_sc_hd__nor2_1 _12406_ (.A(_05490_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__o22ai_1 _12407_ (.A1(_05488_),
    .A2(_05536_),
    .B1(_05578_),
    .B2(_05493_),
    .Y(_05580_));
 sky130_fd_sc_hd__a211oi_1 _12408_ (.A1(_05378_),
    .A2(_05579_),
    .B1(_05580_),
    .C1(_05537_),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_1 _12409_ (.A(_05577_),
    .B(_05581_),
    .Y(_05583_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(_05533_),
    .A1(_05527_),
    .S(_05531_),
    .X(_05584_));
 sky130_fd_sc_hd__nand2_1 _12411_ (.A(_05583_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__or2_1 _12412_ (.A(_05583_),
    .B(_05584_),
    .X(_05586_));
 sky130_fd_sc_hd__a221oi_1 _12413_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05585_),
    .B2(_05586_),
    .C1(_06465_),
    .Y(_05587_));
 sky130_fd_sc_hd__a311o_2 _12414_ (.A1(_05576_),
    .A2(_05585_),
    .A3(_05586_),
    .B1(_05587_),
    .C1(_02246_),
    .X(_05588_));
 sky130_fd_sc_hd__nor2_1 _12415_ (.A(net294),
    .B(_04986_),
    .Y(_05589_));
 sky130_fd_sc_hd__a22o_1 _12416_ (.A1(net295),
    .A2(_06412_),
    .B1(_05553_),
    .B2(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__nor2_1 _12417_ (.A(_05279_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__a211o_1 _12418_ (.A1(_05279_),
    .A2(_05590_),
    .B1(_05591_),
    .C1(net236),
    .X(_05592_));
 sky130_fd_sc_hd__a21oi_1 _12419_ (.A1(net161),
    .A2(_02019_),
    .B1(_02134_),
    .Y(_05594_));
 sky130_fd_sc_hd__and3_1 _12420_ (.A(net161),
    .B(_02019_),
    .C(_02134_),
    .X(_05595_));
 sky130_fd_sc_hd__nand3_1 _12421_ (.A(reg1_val[30]),
    .B(net251),
    .C(_05510_),
    .Y(_05596_));
 sky130_fd_sc_hd__a21oi_1 _12422_ (.A1(_02349_),
    .A2(_05596_),
    .B1(net196),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_1 _12423_ (.A1(_02349_),
    .A2(_05596_),
    .B1(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__o21a_1 _12424_ (.A1(\div_res[30] ),
    .A2(_05559_),
    .B1(net166),
    .X(_05599_));
 sky130_fd_sc_hd__xnor2_1 _12425_ (.A(\div_res[31] ),
    .B(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21a_1 _12426_ (.A1(\div_shifter[62] ),
    .A2(_05564_),
    .B1(net229),
    .X(_05601_));
 sky130_fd_sc_hd__o21ai_1 _12427_ (.A1(\div_shifter[63] ),
    .A2(_05601_),
    .B1(_02336_),
    .Y(_05602_));
 sky130_fd_sc_hd__a21o_1 _12428_ (.A1(\div_shifter[63] ),
    .A2(_05601_),
    .B1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__o21ai_1 _12429_ (.A1(reg1_val[31]),
    .A2(_05258_),
    .B1(_02321_),
    .Y(_05605_));
 sky130_fd_sc_hd__o311a_1 _12430_ (.A1(_04427_),
    .A2(_05247_),
    .A3(_02332_),
    .B1(_05605_),
    .C1(net241),
    .X(_05606_));
 sky130_fd_sc_hd__o221a_1 _12431_ (.A1(_05279_),
    .A2(net235),
    .B1(_02349_),
    .B2(_02320_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__o211a_1 _12432_ (.A1(net168),
    .A2(_02314_),
    .B1(_05603_),
    .C1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__o211a_1 _12433_ (.A1(net183),
    .A2(_05600_),
    .B1(_05608_),
    .C1(_05598_),
    .X(_05609_));
 sky130_fd_sc_hd__o31a_1 _12434_ (.A1(_02330_),
    .A2(_05594_),
    .A3(_05595_),
    .B1(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__o21ai_1 _12435_ (.A1(_05258_),
    .A2(net241),
    .B1(net245),
    .Y(_05611_));
 sky130_fd_sc_hd__a31oi_4 _12436_ (.A1(_05588_),
    .A2(_05592_),
    .A3(_05610_),
    .B1(_05611_),
    .Y(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(net293),
    .A1(curr_PC[0]),
    .S(net244),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _12438_ (.A(_04703_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__or2_1 _12439_ (.A(_04703_),
    .B(_05612_),
    .X(_05615_));
 sky130_fd_sc_hd__and2_4 _12440_ (.A(_05613_),
    .B(_05615_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(net289),
    .A1(curr_PC[1]),
    .S(net244),
    .X(_05616_));
 sky130_fd_sc_hd__nand2_1 _12442_ (.A(_05865_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__or2_1 _12443_ (.A(_05865_),
    .B(_05616_),
    .X(_05618_));
 sky130_fd_sc_hd__nand2_1 _12444_ (.A(_05617_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _12445_ (.A(_05613_),
    .B(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _12446_ (.A(_05613_),
    .B(_05619_),
    .Y(_05621_));
 sky130_fd_sc_hd__and2_4 _12447_ (.A(_05620_),
    .B(_05621_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12448_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net244),
    .X(_05622_));
 sky130_fd_sc_hd__nand2_1 _12449_ (.A(_05811_),
    .B(_05622_),
    .Y(_05624_));
 sky130_fd_sc_hd__or2_1 _12450_ (.A(_05811_),
    .B(_05622_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a21o_1 _12452_ (.A1(_05617_),
    .A2(_05620_),
    .B1(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__nand3_1 _12453_ (.A(_05617_),
    .B(_05620_),
    .C(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__and2_4 _12454_ (.A(_05627_),
    .B(_05628_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net245),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _12456_ (.A(_05738_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__or2_1 _12457_ (.A(_05738_),
    .B(_05629_),
    .X(_05631_));
 sky130_fd_sc_hd__nand2_1 _12458_ (.A(_05630_),
    .B(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__a21o_1 _12459_ (.A1(_05624_),
    .A2(_05627_),
    .B1(_05632_),
    .X(_05634_));
 sky130_fd_sc_hd__nand3_1 _12460_ (.A(_05624_),
    .B(_05627_),
    .C(_05632_),
    .Y(_05635_));
 sky130_fd_sc_hd__and2_4 _12461_ (.A(_05634_),
    .B(_05635_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net245),
    .X(_05636_));
 sky130_fd_sc_hd__nand2_1 _12463_ (.A(_05681_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(_05681_),
    .B(_05636_),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a21o_1 _12466_ (.A1(_05630_),
    .A2(_05634_),
    .B1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__nand3_1 _12467_ (.A(_05630_),
    .B(_05634_),
    .C(_05639_),
    .Y(_05641_));
 sky130_fd_sc_hd__and2_4 _12468_ (.A(_05640_),
    .B(_05641_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net245),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _12470_ (.A(_05528_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__or2_1 _12471_ (.A(_05528_),
    .B(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _12472_ (.A(_05644_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__a21o_1 _12473_ (.A1(_05637_),
    .A2(_05640_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand3_1 _12474_ (.A(_05637_),
    .B(_05640_),
    .C(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__and2_4 _12475_ (.A(_05647_),
    .B(_05648_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net245),
    .X(_05649_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_05593_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__or2_1 _12478_ (.A(_05593_),
    .B(_05649_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2_1 _12479_ (.A(_05650_),
    .B(_05651_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21o_1 _12480_ (.A1(_05644_),
    .A2(_05647_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__nand3_1 _12481_ (.A(_05644_),
    .B(_05647_),
    .C(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_4 _12482_ (.A(_05654_),
    .B(_05655_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(reg1_val[7]),
    .A1(curr_PC[7]),
    .S(net244),
    .X(_05656_));
 sky130_fd_sc_hd__nand2_1 _12484_ (.A(_05453_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__or2_1 _12485_ (.A(_05453_),
    .B(_05656_),
    .X(_05658_));
 sky130_fd_sc_hd__nand2_1 _12486_ (.A(_05657_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a21o_1 _12487_ (.A1(_05650_),
    .A2(_05654_),
    .B1(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__nand3_1 _12488_ (.A(_05650_),
    .B(_05654_),
    .C(_05659_),
    .Y(_05661_));
 sky130_fd_sc_hd__and2_4 _12489_ (.A(_05660_),
    .B(_05661_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net243),
    .X(_05663_));
 sky130_fd_sc_hd__nand2_1 _12491_ (.A(_05388_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__or2_1 _12492_ (.A(_05388_),
    .B(_05663_),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _12493_ (.A(_05664_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__a21o_1 _12494_ (.A1(_05657_),
    .A2(_05660_),
    .B1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__nand3_1 _12495_ (.A(_05657_),
    .B(_05660_),
    .C(_05666_),
    .Y(_05668_));
 sky130_fd_sc_hd__and2_4 _12496_ (.A(_05667_),
    .B(_05668_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_2 _12497_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net244),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_1 _12498_ (.A(_05160_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__or2_1 _12499_ (.A(_05160_),
    .B(_05669_),
    .X(_05672_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_05670_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21o_1 _12501_ (.A1(_05664_),
    .A2(_05667_),
    .B1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__nand3_1 _12502_ (.A(_05664_),
    .B(_05667_),
    .C(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__and2_4 _12503_ (.A(_05674_),
    .B(_05675_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net245),
    .X(_05676_));
 sky130_fd_sc_hd__nand2_1 _12505_ (.A(_05095_),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__or2_1 _12506_ (.A(_05095_),
    .B(_05676_),
    .X(_05678_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_05677_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__a21o_1 _12508_ (.A1(_05670_),
    .A2(_05674_),
    .B1(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__nand3_1 _12509_ (.A(_05670_),
    .B(_05674_),
    .C(_05679_),
    .Y(_05682_));
 sky130_fd_sc_hd__and2_4 _12510_ (.A(_05680_),
    .B(_05682_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_2 _12511_ (.A0(reg1_val[11]),
    .A1(curr_PC[11]),
    .S(net244),
    .X(_05683_));
 sky130_fd_sc_hd__nand2_1 _12512_ (.A(_05290_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__or2_1 _12513_ (.A(_05290_),
    .B(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _12514_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__a21o_1 _12515_ (.A1(_05677_),
    .A2(_05680_),
    .B1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__nand3_1 _12516_ (.A(_05677_),
    .B(_05680_),
    .C(_05686_),
    .Y(_05688_));
 sky130_fd_sc_hd__and2_4 _12517_ (.A(_05687_),
    .B(_05688_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net244),
    .X(_05689_));
 sky130_fd_sc_hd__nand2_1 _12519_ (.A(_05019_),
    .B(_05689_),
    .Y(_05691_));
 sky130_fd_sc_hd__or2_1 _12520_ (.A(_05019_),
    .B(_05689_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _12521_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _12522_ (.A1(_05684_),
    .A2(_05687_),
    .B1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__nand3_1 _12523_ (.A(_05684_),
    .B(_05687_),
    .C(_05693_),
    .Y(_05695_));
 sky130_fd_sc_hd__and2_4 _12524_ (.A(_05694_),
    .B(_05695_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(reg1_val[13]),
    .A1(curr_PC[13]),
    .S(net244),
    .X(_05696_));
 sky130_fd_sc_hd__nand2_1 _12526_ (.A(_04866_),
    .B(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(_04866_),
    .B(_05696_),
    .X(_05698_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_05697_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__a21o_1 _12529_ (.A1(_05691_),
    .A2(_05694_),
    .B1(_05699_),
    .X(_05701_));
 sky130_fd_sc_hd__nand3_1 _12530_ (.A(_05691_),
    .B(_05694_),
    .C(_05699_),
    .Y(_05702_));
 sky130_fd_sc_hd__and2_4 _12531_ (.A(_05701_),
    .B(_05702_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(net291),
    .A1(curr_PC[14]),
    .S(net246),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _12533_ (.A(_04779_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__or2_1 _12534_ (.A(_04779_),
    .B(_05703_),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _12535_ (.A(_05704_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__a21o_1 _12536_ (.A1(_05697_),
    .A2(_05701_),
    .B1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__nand3_1 _12537_ (.A(_05697_),
    .B(_05701_),
    .C(_05706_),
    .Y(_05708_));
 sky130_fd_sc_hd__and2_4 _12538_ (.A(_05707_),
    .B(_05708_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(net290),
    .A1(curr_PC[15]),
    .S(net246),
    .X(_05710_));
 sky130_fd_sc_hd__nand2_1 _12540_ (.A(_04942_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _12541_ (.A(_04942_),
    .B(_05710_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _12542_ (.A(_05711_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21o_1 _12543_ (.A1(_05704_),
    .A2(_05707_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nand3_1 _12544_ (.A(_05704_),
    .B(_05707_),
    .C(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__and2_4 _12545_ (.A(_05714_),
    .B(_05715_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_2 _12546_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net246),
    .X(_05716_));
 sky130_fd_sc_hd__xnor2_1 _12547_ (.A(net264),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__a21o_1 _12548_ (.A1(_05711_),
    .A2(_05714_),
    .B1(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nand3_1 _12549_ (.A(_05711_),
    .B(_05714_),
    .C(_05717_),
    .Y(_05720_));
 sky130_fd_sc_hd__and2_4 _12550_ (.A(_05718_),
    .B(_05720_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12551_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net246),
    .X(_05721_));
 sky130_fd_sc_hd__xnor2_4 _12552_ (.A(net264),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a21bo_1 _12553_ (.A1(net264),
    .A2(_05716_),
    .B1_N(_05718_),
    .X(_05723_));
 sky130_fd_sc_hd__xnor2_4 _12554_ (.A(_05722_),
    .B(_05723_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net246),
    .X(_05724_));
 sky130_fd_sc_hd__nand2_1 _12556_ (.A(net264),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(net264),
    .B(_05724_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_05725_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__or2_1 _12559_ (.A(_05718_),
    .B(_05722_),
    .X(_05729_));
 sky130_fd_sc_hd__o21ai_1 _12560_ (.A1(_05716_),
    .A2(_05721_),
    .B1(net264),
    .Y(_05730_));
 sky130_fd_sc_hd__a21o_1 _12561_ (.A1(_05729_),
    .A2(_05730_),
    .B1(_05727_),
    .X(_05731_));
 sky130_fd_sc_hd__nand3_1 _12562_ (.A(_05727_),
    .B(_05729_),
    .C(_05730_),
    .Y(_05732_));
 sky130_fd_sc_hd__and2_4 _12563_ (.A(_05731_),
    .B(_05732_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net246),
    .X(_05733_));
 sky130_fd_sc_hd__nand2_1 _12565_ (.A(net264),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__or2_1 _12566_ (.A(net264),
    .B(_05733_),
    .X(_05735_));
 sky130_fd_sc_hd__nand2_2 _12567_ (.A(_05734_),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2_2 _12568_ (.A(_05725_),
    .B(_05731_),
    .Y(_05737_));
 sky130_fd_sc_hd__xnor2_4 _12569_ (.A(_05736_),
    .B(_05737_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net246),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_1 _12571_ (.A(net265),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__or2_1 _12572_ (.A(net265),
    .B(_05739_),
    .X(_05741_));
 sky130_fd_sc_hd__nand2_2 _12573_ (.A(_05740_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__or3_1 _12574_ (.A(_05727_),
    .B(_05729_),
    .C(_05736_),
    .X(_05743_));
 sky130_fd_sc_hd__and3_1 _12575_ (.A(_05725_),
    .B(_05730_),
    .C(_05734_),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_2 _12576_ (.A(_05743_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__inv_2 _12577_ (.A(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__xnor2_4 _12578_ (.A(_05742_),
    .B(_05745_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_2 _12579_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net246),
    .X(_05748_));
 sky130_fd_sc_hd__xnor2_4 _12580_ (.A(net264),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_2 _12581_ (.A1(_05742_),
    .A2(_05746_),
    .B1(_05740_),
    .Y(_05750_));
 sky130_fd_sc_hd__xnor2_4 _12582_ (.A(_05749_),
    .B(_05750_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net246),
    .X(_05751_));
 sky130_fd_sc_hd__and2_1 _12584_ (.A(net265),
    .B(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__or2_1 _12585_ (.A(net264),
    .B(_05751_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2b_2 _12586_ (.A_N(_05752_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__o21ai_2 _12587_ (.A1(_05739_),
    .A2(_05748_),
    .B1(net264),
    .Y(_05755_));
 sky130_fd_sc_hd__nor2_1 _12588_ (.A(_05742_),
    .B(_05749_),
    .Y(_05756_));
 sky130_fd_sc_hd__inv_2 _12589_ (.A(_05756_),
    .Y(_05758_));
 sky130_fd_sc_hd__o21ai_4 _12590_ (.A1(_05746_),
    .A2(_05758_),
    .B1(_05755_),
    .Y(_05759_));
 sky130_fd_sc_hd__xnor2_4 _12591_ (.A(_05754_),
    .B(_05759_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_2 _12592_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net246),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_4 _12593_ (.A(net264),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__a21o_1 _12594_ (.A1(_05753_),
    .A2(_05759_),
    .B1(_05752_),
    .X(_05762_));
 sky130_fd_sc_hd__xnor2_4 _12595_ (.A(_05761_),
    .B(_05762_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_2 _12596_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net246),
    .X(_05763_));
 sky130_fd_sc_hd__xnor2_4 _12597_ (.A(net265),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__or4_1 _12598_ (.A(_05743_),
    .B(_05754_),
    .C(_05758_),
    .D(_05761_),
    .X(_05765_));
 sky130_fd_sc_hd__o21ai_1 _12599_ (.A1(_05751_),
    .A2(_05760_),
    .B1(net265),
    .Y(_05767_));
 sky130_fd_sc_hd__and4_2 _12600_ (.A(_05744_),
    .B(_05755_),
    .C(_05765_),
    .D(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__xor2_4 _12601_ (.A(_05764_),
    .B(_05768_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net246),
    .X(_05769_));
 sky130_fd_sc_hd__and2_1 _12603_ (.A(net265),
    .B(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__nor2_1 _12604_ (.A(net264),
    .B(_05769_),
    .Y(_05771_));
 sky130_fd_sc_hd__nor2_2 _12605_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__o2bb2a_2 _12606_ (.A1_N(net264),
    .A2_N(_05763_),
    .B1(_05764_),
    .B2(_05768_),
    .X(_05773_));
 sky130_fd_sc_hd__xnor2_4 _12607_ (.A(_05772_),
    .B(_05773_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net246),
    .X(_05774_));
 sky130_fd_sc_hd__and2_1 _12609_ (.A(net264),
    .B(_05774_),
    .X(_05776_));
 sky130_fd_sc_hd__nor2_1 _12610_ (.A(net264),
    .B(_05774_),
    .Y(_05777_));
 sky130_fd_sc_hd__nor2_2 _12611_ (.A(_05776_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__o21ba_2 _12612_ (.A1(_05771_),
    .A2(_05773_),
    .B1_N(_05770_),
    .X(_05779_));
 sky130_fd_sc_hd__xnor2_4 _12613_ (.A(_05778_),
    .B(_05779_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_2 _12614_ (.A1(_05777_),
    .A2(_05779_),
    .B1_N(_05776_),
    .X(_05780_));
 sky130_fd_sc_hd__mux2_2 _12615_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net246),
    .X(_05781_));
 sky130_fd_sc_hd__xor2_2 _12616_ (.A(net265),
    .B(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__xnor2_4 _12617_ (.A(_05780_),
    .B(_05782_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__nand2_2 _12618_ (.A(net292),
    .B(_04703_),
    .Y(_05783_));
 sky130_fd_sc_hd__or2_1 _12619_ (.A(net292),
    .B(_04703_),
    .X(_05785_));
 sky130_fd_sc_hd__and2_4 _12620_ (.A(_05783_),
    .B(_05785_),
    .X(loadstore_address[0]));
 sky130_fd_sc_hd__or2_1 _12621_ (.A(net289),
    .B(_05865_),
    .X(_05786_));
 sky130_fd_sc_hd__nand2_1 _12622_ (.A(reg1_val[1]),
    .B(_05865_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_2 _12623_ (.A(_05786_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__xor2_4 _12624_ (.A(_05783_),
    .B(_05788_),
    .X(loadstore_address[1]));
 sky130_fd_sc_hd__o21a_2 _12625_ (.A1(_05783_),
    .A2(_05788_),
    .B1(_05787_),
    .X(_05789_));
 sky130_fd_sc_hd__nor2_1 _12626_ (.A(reg1_val[2]),
    .B(_05811_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(reg1_val[2]),
    .B(_05811_),
    .Y(_05791_));
 sky130_fd_sc_hd__and2b_1 _12628_ (.A_N(_05790_),
    .B(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__xnor2_4 _12629_ (.A(_05789_),
    .B(_05792_),
    .Y(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12630_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_05791_),
    .X(_05794_));
 sky130_fd_sc_hd__nor2_1 _12631_ (.A(reg1_val[3]),
    .B(_05738_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_1 _12632_ (.A(reg1_val[3]),
    .B(_05738_),
    .Y(_05796_));
 sky130_fd_sc_hd__and2b_2 _12633_ (.A_N(_05795_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__xnor2_4 _12634_ (.A(_05794_),
    .B(_05797_),
    .Y(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12635_ (.A1(_05794_),
    .A2(_05795_),
    .B1(_05796_),
    .X(_05798_));
 sky130_fd_sc_hd__nor2_1 _12636_ (.A(reg1_val[4]),
    .B(_05681_),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_1 _12637_ (.A(reg1_val[4]),
    .B(_05681_),
    .Y(_05800_));
 sky130_fd_sc_hd__and2b_1 _12638_ (.A_N(_05799_),
    .B(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__xnor2_4 _12639_ (.A(_05798_),
    .B(_05801_),
    .Y(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _12640_ (.A1(_05798_),
    .A2(_05799_),
    .B1(_05800_),
    .X(_05803_));
 sky130_fd_sc_hd__nor2_1 _12641_ (.A(reg1_val[5]),
    .B(_05528_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _12642_ (.A(reg1_val[5]),
    .B(_05528_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand2b_2 _12643_ (.A_N(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__xor2_4 _12644_ (.A(_05803_),
    .B(_05806_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _12645_ (.A1(_05803_),
    .A2(_05804_),
    .B1(_05805_),
    .X(_05807_));
 sky130_fd_sc_hd__nor2_1 _12646_ (.A(reg1_val[6]),
    .B(_05593_),
    .Y(_05808_));
 sky130_fd_sc_hd__and2_1 _12647_ (.A(reg1_val[6]),
    .B(_05593_),
    .X(_05809_));
 sky130_fd_sc_hd__or2_2 _12648_ (.A(_05808_),
    .B(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__xor2_4 _12649_ (.A(_05807_),
    .B(_05810_),
    .X(loadstore_address[6]));
 sky130_fd_sc_hd__o21ba_2 _12650_ (.A1(_05807_),
    .A2(_05808_),
    .B1_N(_05809_),
    .X(_05812_));
 sky130_fd_sc_hd__nor2_1 _12651_ (.A(reg1_val[7]),
    .B(_05453_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_1 _12652_ (.A(reg1_val[7]),
    .B(_05453_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand2b_2 _12653_ (.A_N(_05813_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__xor2_4 _12654_ (.A(_05812_),
    .B(_05815_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _12655_ (.A1(_05812_),
    .A2(_05813_),
    .B1(_05814_),
    .X(_05816_));
 sky130_fd_sc_hd__nor2_1 _12656_ (.A(reg1_val[8]),
    .B(_05388_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _12657_ (.A(reg1_val[8]),
    .B(_05388_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2b_2 _12658_ (.A_N(_05817_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__xor2_4 _12659_ (.A(_05816_),
    .B(_05819_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _12660_ (.A1(_05816_),
    .A2(_05817_),
    .B1(_05818_),
    .X(_05821_));
 sky130_fd_sc_hd__or2_1 _12661_ (.A(reg1_val[9]),
    .B(_05160_),
    .X(_05822_));
 sky130_fd_sc_hd__nand2_1 _12662_ (.A(reg1_val[9]),
    .B(_05160_),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2_2 _12663_ (.A(_05822_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__xor2_4 _12664_ (.A(_05821_),
    .B(_05824_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__nand2_1 _12665_ (.A(reg1_val[10]),
    .B(_05095_),
    .Y(_05825_));
 sky130_fd_sc_hd__or2_1 _12666_ (.A(reg1_val[10]),
    .B(_05095_),
    .X(_05826_));
 sky130_fd_sc_hd__nand2_1 _12667_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2b_1 _12668_ (.A_N(_05821_),
    .B(_05822_),
    .Y(_05828_));
 sky130_fd_sc_hd__a21o_1 _12669_ (.A1(_05823_),
    .A2(_05828_),
    .B1(_05827_),
    .X(_05830_));
 sky130_fd_sc_hd__nand3_1 _12670_ (.A(_05823_),
    .B(_05827_),
    .C(_05828_),
    .Y(_05831_));
 sky130_fd_sc_hd__and2_4 _12671_ (.A(_05830_),
    .B(_05831_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__nand2_1 _12672_ (.A(reg1_val[11]),
    .B(_05290_),
    .Y(_05832_));
 sky130_fd_sc_hd__or2_1 _12673_ (.A(reg1_val[11]),
    .B(_05290_),
    .X(_05833_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21o_1 _12675_ (.A1(_05825_),
    .A2(_05830_),
    .B1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__nand3_1 _12676_ (.A(_05825_),
    .B(_05830_),
    .C(_05834_),
    .Y(_05836_));
 sky130_fd_sc_hd__and2_4 _12677_ (.A(_05835_),
    .B(_05836_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__nand2_1 _12678_ (.A(reg1_val[12]),
    .B(_05019_),
    .Y(_05837_));
 sky130_fd_sc_hd__or2_1 _12679_ (.A(reg1_val[12]),
    .B(_05019_),
    .X(_05839_));
 sky130_fd_sc_hd__nand2_1 _12680_ (.A(_05837_),
    .B(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__a21o_1 _12681_ (.A1(_05832_),
    .A2(_05835_),
    .B1(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__nand3_1 _12682_ (.A(_05832_),
    .B(_05835_),
    .C(_05840_),
    .Y(_05842_));
 sky130_fd_sc_hd__and2_4 _12683_ (.A(_05841_),
    .B(_05842_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__nand2_1 _12684_ (.A(reg1_val[13]),
    .B(_04866_),
    .Y(_05843_));
 sky130_fd_sc_hd__or2_1 _12685_ (.A(reg1_val[13]),
    .B(_04866_),
    .X(_05844_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(_05843_),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__a21o_1 _12687_ (.A1(_05837_),
    .A2(_05841_),
    .B1(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__nand3_1 _12688_ (.A(_05837_),
    .B(_05841_),
    .C(_05845_),
    .Y(_05847_));
 sky130_fd_sc_hd__and2_4 _12689_ (.A(_05846_),
    .B(_05847_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__nand2_1 _12690_ (.A(reg1_val[14]),
    .B(_04779_),
    .Y(_05849_));
 sky130_fd_sc_hd__or2_1 _12691_ (.A(reg1_val[14]),
    .B(_04779_),
    .X(_05850_));
 sky130_fd_sc_hd__nand2_1 _12692_ (.A(_05849_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__a21o_1 _12693_ (.A1(_05843_),
    .A2(_05846_),
    .B1(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__nand3_1 _12694_ (.A(_05843_),
    .B(_05846_),
    .C(_05851_),
    .Y(_05853_));
 sky130_fd_sc_hd__and2_4 _12695_ (.A(_05852_),
    .B(_05853_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _12696_ (.A(reg1_val[15]),
    .B(_04942_),
    .Y(_05854_));
 sky130_fd_sc_hd__a21oi_4 _12697_ (.A1(_05849_),
    .A2(_05852_),
    .B1(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__and3_2 _12698_ (.A(_05849_),
    .B(_05852_),
    .C(_05854_),
    .X(_05856_));
 sky130_fd_sc_hd__nor2_8 _12699_ (.A(_05855_),
    .B(_05856_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__xor2_4 _12700_ (.A(reg1_val[16]),
    .B(net267),
    .X(_05858_));
 sky130_fd_sc_hd__a21o_2 _12701_ (.A1(reg1_val[15]),
    .A2(_04942_),
    .B1(_05855_),
    .X(_05859_));
 sky130_fd_sc_hd__nand2_1 _12702_ (.A(_05858_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__xor2_4 _12703_ (.A(_05858_),
    .B(_05859_),
    .X(loadstore_address[16]));
 sky130_fd_sc_hd__a21bo_1 _12704_ (.A1(reg1_val[16]),
    .A2(net267),
    .B1_N(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__xnor2_4 _12705_ (.A(reg1_val[17]),
    .B(net267),
    .Y(_05862_));
 sky130_fd_sc_hd__xnor2_4 _12706_ (.A(_05861_),
    .B(_05862_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__nand2_2 _12707_ (.A(reg1_val[18]),
    .B(net267),
    .Y(_05863_));
 sky130_fd_sc_hd__or2_1 _12708_ (.A(reg1_val[18]),
    .B(net267),
    .X(_05864_));
 sky130_fd_sc_hd__nand2_4 _12709_ (.A(_05863_),
    .B(_05864_),
    .Y(_05866_));
 sky130_fd_sc_hd__o2bb2a_2 _12710_ (.A1_N(net267),
    .A2_N(_00185_),
    .B1(_05860_),
    .B2(_05862_),
    .X(_05867_));
 sky130_fd_sc_hd__xor2_4 _12711_ (.A(_05866_),
    .B(_05867_),
    .X(loadstore_address[18]));
 sky130_fd_sc_hd__o21ai_4 _12712_ (.A1(_05866_),
    .A2(_05867_),
    .B1(_05863_),
    .Y(_05868_));
 sky130_fd_sc_hd__xnor2_4 _12713_ (.A(reg1_val[19]),
    .B(net267),
    .Y(_05869_));
 sky130_fd_sc_hd__xnor2_4 _12714_ (.A(_05868_),
    .B(_05869_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _12715_ (.A(reg1_val[20]),
    .B(net267),
    .Y(_05870_));
 sky130_fd_sc_hd__or4_2 _12716_ (.A(_05860_),
    .B(_05862_),
    .C(_05866_),
    .D(_05869_),
    .X(_05871_));
 sky130_fd_sc_hd__nand2_1 _12717_ (.A(net267),
    .B(_00186_),
    .Y(_05872_));
 sky130_fd_sc_hd__a21oi_4 _12718_ (.A1(_05871_),
    .A2(_05872_),
    .B1(_05870_),
    .Y(_05873_));
 sky130_fd_sc_hd__and3_2 _12719_ (.A(_05870_),
    .B(_05871_),
    .C(_05872_),
    .X(_05875_));
 sky130_fd_sc_hd__nor2_8 _12720_ (.A(_05873_),
    .B(_05875_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _12721_ (.A(reg1_val[21]),
    .B(net266),
    .Y(_05876_));
 sky130_fd_sc_hd__nand2_1 _12722_ (.A(reg1_val[21]),
    .B(net266),
    .Y(_05877_));
 sky130_fd_sc_hd__nand2b_2 _12723_ (.A_N(_05876_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21oi_4 _12724_ (.A1(reg1_val[20]),
    .A2(net267),
    .B1(_05873_),
    .Y(_05879_));
 sky130_fd_sc_hd__xor2_4 _12725_ (.A(_05878_),
    .B(_05879_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__nand2_2 _12726_ (.A(reg1_val[22]),
    .B(net266),
    .Y(_05880_));
 sky130_fd_sc_hd__or2_1 _12727_ (.A(reg1_val[22]),
    .B(net266),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_4 _12728_ (.A(_05880_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__o21a_2 _12729_ (.A1(_05876_),
    .A2(_05879_),
    .B1(_05877_),
    .X(_05884_));
 sky130_fd_sc_hd__xor2_4 _12730_ (.A(_05882_),
    .B(_05884_),
    .X(loadstore_address[22]));
 sky130_fd_sc_hd__o21ai_4 _12731_ (.A1(_05882_),
    .A2(_05884_),
    .B1(_05880_),
    .Y(_05885_));
 sky130_fd_sc_hd__xnor2_4 _12732_ (.A(reg1_val[23]),
    .B(net266),
    .Y(_05886_));
 sky130_fd_sc_hd__xnor2_4 _12733_ (.A(_05885_),
    .B(_05886_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__nand2_1 _12734_ (.A(reg1_val[24]),
    .B(net266),
    .Y(_05887_));
 sky130_fd_sc_hd__or2_1 _12735_ (.A(reg1_val[24]),
    .B(net266),
    .X(_05888_));
 sky130_fd_sc_hd__nand2_2 _12736_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__or4_1 _12737_ (.A(_05870_),
    .B(_05878_),
    .C(_05882_),
    .D(_05886_),
    .X(_05890_));
 sky130_fd_sc_hd__a2bb2o_2 _12738_ (.A1_N(_05871_),
    .A2_N(_05890_),
    .B1(net267),
    .B2(_00217_),
    .X(_05891_));
 sky130_fd_sc_hd__nand2b_1 _12739_ (.A_N(_05889_),
    .B(_05891_),
    .Y(_05893_));
 sky130_fd_sc_hd__xnor2_4 _12740_ (.A(_05889_),
    .B(_05891_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _12741_ (.A(_05887_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__xnor2_2 _12742_ (.A(reg1_val[25]),
    .B(net266),
    .Y(_05895_));
 sky130_fd_sc_hd__xnor2_4 _12743_ (.A(_05894_),
    .B(_05895_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__and2_1 _12744_ (.A(reg1_val[26]),
    .B(net266),
    .X(_05896_));
 sky130_fd_sc_hd__or2_1 _12745_ (.A(reg1_val[26]),
    .B(net266),
    .X(_05897_));
 sky130_fd_sc_hd__nand2b_2 _12746_ (.A_N(_05896_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__or2_1 _12747_ (.A(_05893_),
    .B(_05895_),
    .X(_05899_));
 sky130_fd_sc_hd__a21bo_2 _12748_ (.A1(net267),
    .A2(_00219_),
    .B1_N(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__xnor2_4 _12749_ (.A(_05898_),
    .B(_05900_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21o_1 _12750_ (.A1(_05897_),
    .A2(_05900_),
    .B1(_05896_),
    .X(_05902_));
 sky130_fd_sc_hd__xnor2_2 _12751_ (.A(reg1_val[27]),
    .B(net266),
    .Y(_05903_));
 sky130_fd_sc_hd__xnor2_4 _12752_ (.A(_05902_),
    .B(_05903_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__and2_1 _12753_ (.A(reg1_val[28]),
    .B(net266),
    .X(_05904_));
 sky130_fd_sc_hd__nor2_1 _12754_ (.A(reg1_val[28]),
    .B(net266),
    .Y(_05905_));
 sky130_fd_sc_hd__or2_1 _12755_ (.A(_05904_),
    .B(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__nand2_1 _12756_ (.A(net266),
    .B(_00439_),
    .Y(_05907_));
 sky130_fd_sc_hd__or3_1 _12757_ (.A(_05898_),
    .B(_05899_),
    .C(_05903_),
    .X(_05908_));
 sky130_fd_sc_hd__a21oi_2 _12758_ (.A1(_05907_),
    .A2(_05908_),
    .B1(_05906_),
    .Y(_05909_));
 sky130_fd_sc_hd__and3_2 _12759_ (.A(_05906_),
    .B(_05907_),
    .C(_05908_),
    .X(_05911_));
 sky130_fd_sc_hd__nor2_8 _12760_ (.A(_05909_),
    .B(_05911_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__or2_1 _12761_ (.A(reg1_val[29]),
    .B(net267),
    .X(_05912_));
 sky130_fd_sc_hd__nand2_1 _12762_ (.A(reg1_val[29]),
    .B(net267),
    .Y(_05913_));
 sky130_fd_sc_hd__nand2_2 _12763_ (.A(_05912_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__or2_2 _12764_ (.A(_05904_),
    .B(_05909_),
    .X(_05915_));
 sky130_fd_sc_hd__xnor2_4 _12765_ (.A(_05914_),
    .B(_05915_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__and2_1 _12766_ (.A(reg1_val[30]),
    .B(net266),
    .X(_05916_));
 sky130_fd_sc_hd__or2_1 _12767_ (.A(reg1_val[30]),
    .B(net267),
    .X(_05917_));
 sky130_fd_sc_hd__nand2b_2 _12768_ (.A_N(_05916_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a21bo_2 _12769_ (.A1(_05912_),
    .A2(_05915_),
    .B1_N(_05913_),
    .X(_05920_));
 sky130_fd_sc_hd__xnor2_4 _12770_ (.A(_05918_),
    .B(_05920_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21oi_1 _12771_ (.A1(_05917_),
    .A2(_05920_),
    .B1(_05916_),
    .Y(_05921_));
 sky130_fd_sc_hd__xnor2_2 _12772_ (.A(_04427_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__xnor2_4 _12773_ (.A(net266),
    .B(_05922_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__nand2_1 _12774_ (.A(net488),
    .B(net444),
    .Y(_05923_));
 sky130_fd_sc_hd__nand3_1 _12775_ (.A(net492),
    .B(net488),
    .C(net444),
    .Y(_05924_));
 sky130_fd_sc_hd__and4_1 _12776_ (.A(net449),
    .B(net492),
    .C(net488),
    .D(net444),
    .X(_05925_));
 sky130_fd_sc_hd__inv_2 _12777_ (.A(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_1 _12778_ (.A(net296),
    .B(_05925_),
    .Y(_05927_));
 sky130_fd_sc_hd__nor2_1 _12779_ (.A(_04383_),
    .B(net493),
    .Y(_05929_));
 sky130_fd_sc_hd__nor3_1 _12780_ (.A(rst),
    .B(net204),
    .C(_05929_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_2 _12781_ (.A(net260),
    .B(_06438_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_4 _12782_ (.A(_04383_),
    .B(_06437_),
    .Y(_05931_));
 sky130_fd_sc_hd__or2_1 _12783_ (.A(net304),
    .B(net182),
    .X(_05932_));
 sky130_fd_sc_hd__o211a_1 _12784_ (.A1(_02081_),
    .A2(net178),
    .B1(net305),
    .C1(net283),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _12785_ (.A(net210),
    .B(net180),
    .Y(_05933_));
 sky130_fd_sc_hd__o211a_1 _12786_ (.A1(net298),
    .A2(net180),
    .B1(_05933_),
    .C1(net282),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _12787_ (.A(net460),
    .B(net180),
    .X(_05934_));
 sky130_fd_sc_hd__o211a_1 _12788_ (.A1(_00225_),
    .A2(net177),
    .B1(net461),
    .C1(net282),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _12789_ (.A(net341),
    .B(net180),
    .X(_05936_));
 sky130_fd_sc_hd__o211a_1 _12790_ (.A1(_00250_),
    .A2(net177),
    .B1(net342),
    .C1(net282),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _12791_ (.A(net343),
    .B(net180),
    .X(_05937_));
 sky130_fd_sc_hd__o211a_1 _12792_ (.A1(_00243_),
    .A2(net177),
    .B1(net344),
    .C1(net282),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _12793_ (.A(net399),
    .B(net180),
    .X(_05938_));
 sky130_fd_sc_hd__o211a_1 _12794_ (.A1(_00211_),
    .A2(net177),
    .B1(net400),
    .C1(net282),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _12795_ (.A(net316),
    .B(net180),
    .X(_05939_));
 sky130_fd_sc_hd__o211a_1 _12796_ (.A1(_00198_),
    .A2(net177),
    .B1(net317),
    .C1(net282),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _12797_ (.A(net336),
    .B(net180),
    .X(_05940_));
 sky130_fd_sc_hd__o211a_1 _12798_ (.A1(_00360_),
    .A2(net177),
    .B1(net337),
    .C1(net282),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _12799_ (.A(net324),
    .B(net182),
    .X(_05942_));
 sky130_fd_sc_hd__o211a_1 _12800_ (.A1(_00299_),
    .A2(net178),
    .B1(net325),
    .C1(net283),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(net310),
    .B(net182),
    .X(_05943_));
 sky130_fd_sc_hd__o211a_1 _12802_ (.A1(_00293_),
    .A2(net178),
    .B1(net311),
    .C1(net283),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _12803_ (.A(net333),
    .B(net179),
    .X(_05944_));
 sky130_fd_sc_hd__o211a_1 _12804_ (.A1(_00315_),
    .A2(_05931_),
    .B1(net334),
    .C1(net283),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _12805_ (.A(net327),
    .B(net179),
    .X(_05945_));
 sky130_fd_sc_hd__o211a_1 _12806_ (.A1(_00309_),
    .A2(net176),
    .B1(net328),
    .C1(net278),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _12807_ (.A(net390),
    .B(_05930_),
    .X(_05946_));
 sky130_fd_sc_hd__o211a_1 _12808_ (.A1(_00276_),
    .A2(net176),
    .B1(net391),
    .C1(net278),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _12809_ (.A(net330),
    .B(net179),
    .X(_05948_));
 sky130_fd_sc_hd__o211a_1 _12810_ (.A1(_00272_),
    .A2(net176),
    .B1(net331),
    .C1(net275),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _12811_ (.A(net351),
    .B(net179),
    .X(_05949_));
 sky130_fd_sc_hd__o211a_1 _12812_ (.A1(_00352_),
    .A2(net176),
    .B1(net352),
    .C1(net275),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _12813_ (.A(net348),
    .B(net179),
    .X(_05950_));
 sky130_fd_sc_hd__o211a_1 _12814_ (.A1(_00347_),
    .A2(net176),
    .B1(net349),
    .C1(net276),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _12815_ (.A(net375),
    .B(net179),
    .X(_05951_));
 sky130_fd_sc_hd__o211a_1 _12816_ (.A1(_00340_),
    .A2(net176),
    .B1(net376),
    .C1(net276),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _12817_ (.A(net369),
    .B(net179),
    .X(_05952_));
 sky130_fd_sc_hd__o211a_1 _12818_ (.A1(_00334_),
    .A2(net176),
    .B1(net370),
    .C1(net277),
    .X(_00018_));
 sky130_fd_sc_hd__or2_1 _12819_ (.A(net345),
    .B(net179),
    .X(_05954_));
 sky130_fd_sc_hd__o211a_1 _12820_ (.A1(_00174_),
    .A2(_05931_),
    .B1(net346),
    .C1(net277),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _12821_ (.A(net434),
    .B(net179),
    .X(_05955_));
 sky130_fd_sc_hd__o211a_1 _12822_ (.A1(_00164_),
    .A2(_05931_),
    .B1(net435),
    .C1(net277),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _12823_ (.A(net354),
    .B(net179),
    .X(_05956_));
 sky130_fd_sc_hd__o211a_1 _12824_ (.A1(_00157_),
    .A2(net176),
    .B1(net355),
    .C1(net275),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _12825_ (.A(net381),
    .B(net179),
    .X(_05957_));
 sky130_fd_sc_hd__o211a_1 _12826_ (.A1(_00148_),
    .A2(net176),
    .B1(net382),
    .C1(net276),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _12827_ (.A(net360),
    .B(net179),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _12828_ (.A1(_06522_),
    .A2(net176),
    .B1(net361),
    .C1(net276),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _12829_ (.A(net372),
    .B(net179),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_1 _12830_ (.A1(_06515_),
    .A2(net176),
    .B1(net373),
    .C1(net276),
    .X(_00024_));
 sky130_fd_sc_hd__or2_1 _12831_ (.A(net396),
    .B(net179),
    .X(_05961_));
 sky130_fd_sc_hd__o211a_1 _12832_ (.A1(_06538_),
    .A2(_05931_),
    .B1(net397),
    .C1(net277),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _12833_ (.A(net403),
    .B(net179),
    .X(_05962_));
 sky130_fd_sc_hd__o211a_1 _12834_ (.A1(_06534_),
    .A2(net176),
    .B1(net404),
    .C1(net278),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _12835_ (.A(net415),
    .B(_05930_),
    .X(_05963_));
 sky130_fd_sc_hd__o211a_1 _12836_ (.A1(_06500_),
    .A2(net176),
    .B1(net416),
    .C1(net277),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _12837_ (.A(net393),
    .B(_05930_),
    .X(_05964_));
 sky130_fd_sc_hd__o211a_1 _12838_ (.A1(_06492_),
    .A2(net176),
    .B1(net394),
    .C1(net277),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _12839_ (.A(net366),
    .B(_05930_),
    .X(_05966_));
 sky130_fd_sc_hd__o211a_1 _12840_ (.A1(_06553_),
    .A2(net176),
    .B1(net367),
    .C1(net277),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _12841_ (.A(net409),
    .B(net179),
    .X(_05967_));
 sky130_fd_sc_hd__o211a_1 _12842_ (.A1(_00398_),
    .A2(net176),
    .B1(net410),
    .C1(net277),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _12843_ (.A(net424),
    .B(net182),
    .X(_05968_));
 sky130_fd_sc_hd__o211a_1 _12844_ (.A1(_00690_),
    .A2(net178),
    .B1(net425),
    .C1(net283),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _12845_ (.A(net363),
    .B(net182),
    .X(_05969_));
 sky130_fd_sc_hd__o211a_1 _12846_ (.A1(_01954_),
    .A2(net178),
    .B1(net364),
    .C1(net283),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12847_ (.A(net357),
    .B(net182),
    .X(_05970_));
 sky130_fd_sc_hd__o211a_1 _12848_ (.A1(_02069_),
    .A2(net178),
    .B1(net358),
    .C1(net283),
    .X(_00033_));
 sky130_fd_sc_hd__and2b_1 _12849_ (.A_N(net363),
    .B(\div_shifter[61] ),
    .X(_05972_));
 sky130_fd_sc_hd__and2b_1 _12850_ (.A_N(\div_shifter[61] ),
    .B(net363),
    .X(_05973_));
 sky130_fd_sc_hd__nor2_1 _12851_ (.A(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2b_1 _12852_ (.A_N(\div_shifter[60] ),
    .B(net424),
    .Y(_05975_));
 sky130_fd_sc_hd__and2b_1 _12853_ (.A_N(net409),
    .B(net596),
    .X(_05976_));
 sky130_fd_sc_hd__nand2b_1 _12854_ (.A_N(net586),
    .B(net366),
    .Y(_05977_));
 sky130_fd_sc_hd__and2b_1 _12855_ (.A_N(net393),
    .B(net564),
    .X(_05978_));
 sky130_fd_sc_hd__nand2b_1 _12856_ (.A_N(net564),
    .B(net393),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2b_1 _12857_ (.A_N(_05978_),
    .B(_05979_),
    .Y(_05980_));
 sky130_fd_sc_hd__nand2b_1 _12858_ (.A_N(\div_shifter[56] ),
    .B(net415),
    .Y(_05981_));
 sky130_fd_sc_hd__and2b_1 _12859_ (.A_N(net403),
    .B(net584),
    .X(_05983_));
 sky130_fd_sc_hd__nand2b_1 _12860_ (.A_N(\div_shifter[54] ),
    .B(net396),
    .Y(_05984_));
 sky130_fd_sc_hd__and2b_1 _12861_ (.A_N(net372),
    .B(net594),
    .X(_05985_));
 sky130_fd_sc_hd__nand2b_1 _12862_ (.A_N(net597),
    .B(net360),
    .Y(_05986_));
 sky130_fd_sc_hd__and2b_1 _12863_ (.A_N(net381),
    .B(net570),
    .X(_05987_));
 sky130_fd_sc_hd__nand2b_1 _12864_ (.A_N(net590),
    .B(net354),
    .Y(_05988_));
 sky130_fd_sc_hd__and2b_1 _12865_ (.A_N(net434),
    .B(net576),
    .X(_05989_));
 sky130_fd_sc_hd__nand2b_1 _12866_ (.A_N(net576),
    .B(net434),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2b_1 _12867_ (.A_N(\div_shifter[48] ),
    .B(net345),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2b_1 _12868_ (.A_N(net592),
    .B(net369),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2b_1 _12869_ (.A_N(net606),
    .B(net375),
    .Y(_05994_));
 sky130_fd_sc_hd__nand2b_1 _12870_ (.A_N(\div_shifter[45] ),
    .B(net348),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2b_1 _12871_ (.A_N(net572),
    .B(net351),
    .Y(_05996_));
 sky130_fd_sc_hd__nand2b_1 _12872_ (.A_N(net600),
    .B(net330),
    .Y(_05997_));
 sky130_fd_sc_hd__nand2b_1 _12873_ (.A_N(\div_shifter[42] ),
    .B(net390),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2b_1 _12874_ (.A_N(net598),
    .B(net327),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2b_1 _12875_ (.A_N(net578),
    .B(net333),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2b_1 _12876_ (.A_N(\div_shifter[39] ),
    .B(net310),
    .Y(_06001_));
 sky130_fd_sc_hd__nand2b_1 _12877_ (.A_N(net604),
    .B(net324),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2b_1 _12878_ (.A_N(net588),
    .B(net336),
    .Y(_06003_));
 sky130_fd_sc_hd__and2b_1 _12879_ (.A_N(net316),
    .B(\div_shifter[36] ),
    .X(_06005_));
 sky130_fd_sc_hd__nand2b_1 _12880_ (.A_N(\div_shifter[36] ),
    .B(net316),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2b_1 _12881_ (.A_N(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__and2b_1 _12882_ (.A_N(net399),
    .B(net566),
    .X(_06008_));
 sky130_fd_sc_hd__nand2b_1 _12883_ (.A_N(net566),
    .B(net399),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2b_1 _12884_ (.A_N(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2b_1 _12885_ (.A_N(\div_shifter[34] ),
    .B(net343),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2b_1 _12886_ (.A_N(net560),
    .B(net341),
    .Y(_06012_));
 sky130_fd_sc_hd__and2b_1 _12887_ (.A_N(net460),
    .B(\div_shifter[32] ),
    .X(_06013_));
 sky130_fd_sc_hd__xnor2_1 _12888_ (.A(\div_shifter[32] ),
    .B(net460),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2b_1 _12889_ (.A_N(net568),
    .B(net298),
    .Y(_06016_));
 sky130_fd_sc_hd__a21o_1 _12890_ (.A1(_06014_),
    .A2(_06016_),
    .B1(_06013_),
    .X(_06017_));
 sky130_fd_sc_hd__nand2b_1 _12891_ (.A_N(net341),
    .B(net560),
    .Y(_06018_));
 sky130_fd_sc_hd__a21bo_1 _12892_ (.A1(_06012_),
    .A2(_06017_),
    .B1_N(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__nand2b_1 _12893_ (.A_N(net343),
    .B(\div_shifter[34] ),
    .Y(_06020_));
 sky130_fd_sc_hd__a21bo_1 _12894_ (.A1(_06011_),
    .A2(_06019_),
    .B1_N(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__a21o_1 _12895_ (.A1(_06009_),
    .A2(_06021_),
    .B1(_06008_),
    .X(_06022_));
 sky130_fd_sc_hd__a21o_1 _12896_ (.A1(_06006_),
    .A2(_06022_),
    .B1(_06005_),
    .X(_06023_));
 sky130_fd_sc_hd__nand2b_1 _12897_ (.A_N(net336),
    .B(net588),
    .Y(_06024_));
 sky130_fd_sc_hd__a21bo_1 _12898_ (.A1(_06003_),
    .A2(_06023_),
    .B1_N(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__nand2b_1 _12899_ (.A_N(net324),
    .B(net604),
    .Y(_06027_));
 sky130_fd_sc_hd__a21bo_1 _12900_ (.A1(_06002_),
    .A2(_06025_),
    .B1_N(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2b_1 _12901_ (.A_N(net310),
    .B(\div_shifter[39] ),
    .Y(_06029_));
 sky130_fd_sc_hd__a21bo_1 _12902_ (.A1(_06001_),
    .A2(_06028_),
    .B1_N(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__nand2b_1 _12903_ (.A_N(net333),
    .B(net578),
    .Y(_06031_));
 sky130_fd_sc_hd__a21bo_1 _12904_ (.A1(_06000_),
    .A2(_06030_),
    .B1_N(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__nand2b_1 _12905_ (.A_N(net327),
    .B(net598),
    .Y(_06033_));
 sky130_fd_sc_hd__a21bo_1 _12906_ (.A1(_05999_),
    .A2(_06032_),
    .B1_N(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__nand2b_1 _12907_ (.A_N(net390),
    .B(\div_shifter[42] ),
    .Y(_06035_));
 sky130_fd_sc_hd__a21bo_1 _12908_ (.A1(_05998_),
    .A2(_06034_),
    .B1_N(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__nand2b_1 _12909_ (.A_N(net330),
    .B(net600),
    .Y(_06038_));
 sky130_fd_sc_hd__a21bo_1 _12910_ (.A1(_05997_),
    .A2(_06036_),
    .B1_N(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__nand2b_1 _12911_ (.A_N(net351),
    .B(net572),
    .Y(_06040_));
 sky130_fd_sc_hd__a21bo_1 _12912_ (.A1(_05996_),
    .A2(_06039_),
    .B1_N(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2b_1 _12913_ (.A_N(net348),
    .B(\div_shifter[45] ),
    .Y(_06042_));
 sky130_fd_sc_hd__a21bo_1 _12914_ (.A1(_05995_),
    .A2(_06041_),
    .B1_N(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__nand2b_1 _12915_ (.A_N(net375),
    .B(net606),
    .Y(_06044_));
 sky130_fd_sc_hd__a21bo_1 _12916_ (.A1(_05994_),
    .A2(_06043_),
    .B1_N(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__nand2b_1 _12917_ (.A_N(net369),
    .B(net592),
    .Y(_06046_));
 sky130_fd_sc_hd__a21bo_1 _12918_ (.A1(_05992_),
    .A2(_06045_),
    .B1_N(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__nand2b_1 _12919_ (.A_N(net345),
    .B(\div_shifter[48] ),
    .Y(_06049_));
 sky130_fd_sc_hd__a21bo_1 _12920_ (.A1(_05991_),
    .A2(_06047_),
    .B1_N(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__a21o_1 _12921_ (.A1(_05990_),
    .A2(_06050_),
    .B1(_05989_),
    .X(_06051_));
 sky130_fd_sc_hd__nand2b_1 _12922_ (.A_N(net354),
    .B(net590),
    .Y(_06052_));
 sky130_fd_sc_hd__a21bo_1 _12923_ (.A1(_05988_),
    .A2(_06051_),
    .B1_N(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__nand2b_1 _12924_ (.A_N(net570),
    .B(net381),
    .Y(_06054_));
 sky130_fd_sc_hd__nand2b_1 _12925_ (.A_N(_05987_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__a21o_1 _12926_ (.A1(_06053_),
    .A2(_06054_),
    .B1(_05987_),
    .X(_06056_));
 sky130_fd_sc_hd__nand2b_1 _12927_ (.A_N(net360),
    .B(net597),
    .Y(_06057_));
 sky130_fd_sc_hd__a21bo_1 _12928_ (.A1(_05986_),
    .A2(_06056_),
    .B1_N(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__nand2b_1 _12929_ (.A_N(net594),
    .B(net372),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2b_1 _12930_ (.A_N(_05985_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__a21o_1 _12931_ (.A1(_06058_),
    .A2(_06060_),
    .B1(_05985_),
    .X(_06062_));
 sky130_fd_sc_hd__nand2b_1 _12932_ (.A_N(net396),
    .B(\div_shifter[54] ),
    .Y(_06063_));
 sky130_fd_sc_hd__a21bo_1 _12933_ (.A1(_05984_),
    .A2(_06062_),
    .B1_N(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__nand2b_1 _12934_ (.A_N(net584),
    .B(net403),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2b_1 _12935_ (.A_N(_05983_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__a21o_1 _12936_ (.A1(_06064_),
    .A2(_06065_),
    .B1(_05983_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2b_1 _12937_ (.A_N(net415),
    .B(\div_shifter[56] ),
    .Y(_06068_));
 sky130_fd_sc_hd__a21bo_1 _12938_ (.A1(_05981_),
    .A2(_06067_),
    .B1_N(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__a21o_1 _12939_ (.A1(_05979_),
    .A2(_06069_),
    .B1(_05978_),
    .X(_06071_));
 sky130_fd_sc_hd__nand2b_1 _12940_ (.A_N(net366),
    .B(net586),
    .Y(_06072_));
 sky130_fd_sc_hd__a21bo_1 _12941_ (.A1(_05977_),
    .A2(_06071_),
    .B1_N(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__nand2b_1 _12942_ (.A_N(net596),
    .B(net409),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2b_1 _12943_ (.A_N(_05976_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__a21o_1 _12944_ (.A1(_06073_),
    .A2(_06074_),
    .B1(_05976_),
    .X(_06076_));
 sky130_fd_sc_hd__nand2b_1 _12945_ (.A_N(net424),
    .B(\div_shifter[60] ),
    .Y(_06077_));
 sky130_fd_sc_hd__a21boi_1 _12946_ (.A1(_05975_),
    .A2(_06076_),
    .B1_N(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__o21ba_1 _12947_ (.A1(_05973_),
    .A2(_06078_),
    .B1_N(_05972_),
    .X(_06079_));
 sky130_fd_sc_hd__nor2_1 _12948_ (.A(net357),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__a21boi_1 _12949_ (.A1(net357),
    .A2(_06079_),
    .B1_N(net574),
    .Y(_06082_));
 sky130_fd_sc_hd__or2_1 _12950_ (.A(_06080_),
    .B(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__a22o_1 _12951_ (.A1(net616),
    .A2(net202),
    .B1(net3),
    .B2(net257),
    .X(_06084_));
 sky130_fd_sc_hd__and2_1 _12952_ (.A(net279),
    .B(_06084_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _12953_ (.A1(\div_res[0] ),
    .A2(net256),
    .B1(net202),
    .B2(net580),
    .X(_06085_));
 sky130_fd_sc_hd__and2_1 _12954_ (.A(net279),
    .B(net581),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _12955_ (.A1(\div_res[1] ),
    .A2(net256),
    .B1(net202),
    .B2(net562),
    .X(_06086_));
 sky130_fd_sc_hd__and2_1 _12956_ (.A(net279),
    .B(net563),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _12957_ (.A1(net620),
    .A2(net256),
    .B1(net202),
    .B2(net525),
    .X(_06087_));
 sky130_fd_sc_hd__and2_1 _12958_ (.A(net279),
    .B(net526),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _12959_ (.A1(net525),
    .A2(net256),
    .B1(net202),
    .B2(net556),
    .X(_06089_));
 sky130_fd_sc_hd__and2_1 _12960_ (.A(net279),
    .B(net557),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _12961_ (.A1(\div_res[4] ),
    .A2(net256),
    .B1(net202),
    .B2(net517),
    .X(_06090_));
 sky130_fd_sc_hd__and2_1 _12962_ (.A(net279),
    .B(net518),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _12963_ (.A1(net517),
    .A2(net256),
    .B1(net202),
    .B2(net527),
    .X(_06091_));
 sky130_fd_sc_hd__and2_1 _12964_ (.A(net279),
    .B(net528),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _12965_ (.A1(net527),
    .A2(net256),
    .B1(net202),
    .B2(net542),
    .X(_06092_));
 sky130_fd_sc_hd__and2_1 _12966_ (.A(net279),
    .B(net543),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _12967_ (.A1(net542),
    .A2(net256),
    .B1(net202),
    .B2(net552),
    .X(_06093_));
 sky130_fd_sc_hd__and2_1 _12968_ (.A(net279),
    .B(net553),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _12969_ (.A1(\div_res[8] ),
    .A2(net256),
    .B1(net202),
    .B2(net508),
    .X(_06095_));
 sky130_fd_sc_hd__and2_1 _12970_ (.A(net279),
    .B(net509),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _12971_ (.A1(net508),
    .A2(net256),
    .B1(net202),
    .B2(net535),
    .X(_06096_));
 sky130_fd_sc_hd__and2_1 _12972_ (.A(net279),
    .B(net536),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _12973_ (.A1(\div_res[10] ),
    .A2(net256),
    .B1(net202),
    .B2(net502),
    .X(_06097_));
 sky130_fd_sc_hd__and2_1 _12974_ (.A(net279),
    .B(net503),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _12975_ (.A1(net502),
    .A2(net256),
    .B1(net202),
    .B2(net515),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _12976_ (.A(net279),
    .B(net516),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _12977_ (.A1(net515),
    .A2(net256),
    .B1(net202),
    .B2(net554),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _12978_ (.A(net279),
    .B(net555),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _12979_ (.A1(\div_res[13] ),
    .A2(net258),
    .B1(net200),
    .B2(net529),
    .X(_06101_));
 sky130_fd_sc_hd__and2_1 _12980_ (.A(net275),
    .B(net530),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _12981_ (.A1(\div_res[14] ),
    .A2(net258),
    .B1(net200),
    .B2(net505),
    .X(_06102_));
 sky130_fd_sc_hd__and2_1 _12982_ (.A(net275),
    .B(net506),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _12983_ (.A1(net505),
    .A2(net258),
    .B1(net200),
    .B2(net540),
    .X(_06103_));
 sky130_fd_sc_hd__and2_1 _12984_ (.A(net275),
    .B(net541),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _12985_ (.A1(net621),
    .A2(net258),
    .B1(net200),
    .B2(net511),
    .X(_06104_));
 sky130_fd_sc_hd__and2_1 _12986_ (.A(net275),
    .B(net512),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _12987_ (.A1(net511),
    .A2(net258),
    .B1(net200),
    .B2(net550),
    .X(_06105_));
 sky130_fd_sc_hd__and2_1 _12988_ (.A(net275),
    .B(net551),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _12989_ (.A1(\div_res[18] ),
    .A2(net258),
    .B1(net200),
    .B2(net532),
    .X(_06107_));
 sky130_fd_sc_hd__and2_1 _12990_ (.A(net275),
    .B(net533),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _12991_ (.A1(\div_res[19] ),
    .A2(net258),
    .B1(net200),
    .B2(net520),
    .X(_06108_));
 sky130_fd_sc_hd__and2_1 _12992_ (.A(net275),
    .B(net521),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _12993_ (.A1(net520),
    .A2(net258),
    .B1(net200),
    .B2(net513),
    .X(_06109_));
 sky130_fd_sc_hd__and2_1 _12994_ (.A(net275),
    .B(net545),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _12995_ (.A1(net513),
    .A2(net258),
    .B1(net200),
    .B2(net494),
    .X(_06110_));
 sky130_fd_sc_hd__and2_1 _12996_ (.A(net275),
    .B(net514),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _12997_ (.A1(net494),
    .A2(net259),
    .B1(net200),
    .B2(\div_res[23] ),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12998_ (.A(net275),
    .B(net495),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _12999_ (.A1(net499),
    .A2(net258),
    .B1(net201),
    .B2(\div_res[24] ),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _13000_ (.A(net275),
    .B(net500),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _13001_ (.A1(net523),
    .A2(net258),
    .B1(net201),
    .B2(net483),
    .X(_06114_));
 sky130_fd_sc_hd__and2_1 _13002_ (.A(net278),
    .B(net524),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _13003_ (.A1(net483),
    .A2(net258),
    .B1(net201),
    .B2(\div_res[26] ),
    .X(_06115_));
 sky130_fd_sc_hd__and2_1 _13004_ (.A(net278),
    .B(net484),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _13005_ (.A1(\div_res[26] ),
    .A2(net260),
    .B1(net201),
    .B2(net537),
    .X(_06116_));
 sky130_fd_sc_hd__and2_1 _13006_ (.A(net278),
    .B(net538),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _13007_ (.A1(net537),
    .A2(net260),
    .B1(net201),
    .B2(net546),
    .X(_06117_));
 sky130_fd_sc_hd__and2_1 _13008_ (.A(net278),
    .B(net547),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _13009_ (.A1(net546),
    .A2(net260),
    .B1(net204),
    .B2(net548),
    .X(_06119_));
 sky130_fd_sc_hd__and2_1 _13010_ (.A(net278),
    .B(net549),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _13011_ (.A1(net548),
    .A2(net261),
    .B1(net203),
    .B2(net558),
    .X(_06120_));
 sky130_fd_sc_hd__and2_1 _13012_ (.A(_04448_),
    .B(net559),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _13013_ (.A1(\div_res[30] ),
    .A2(net261),
    .B1(net203),
    .B2(net457),
    .X(_06121_));
 sky130_fd_sc_hd__and2_1 _13014_ (.A(net277),
    .B(net458),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _13015_ (.A1(net442),
    .A2(net203),
    .B1(net181),
    .B2(net293),
    .X(_06122_));
 sky130_fd_sc_hd__and2_1 _13016_ (.A(net281),
    .B(net443),
    .X(_00066_));
 sky130_fd_sc_hd__o221a_1 _13017_ (.A1(\div_shifter[0] ),
    .A2(net254),
    .B1(net198),
    .B2(net378),
    .C1(net281),
    .X(_06123_));
 sky130_fd_sc_hd__o21a_1 _13018_ (.A1(net240),
    .A2(net177),
    .B1(net379),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _13019_ (.A1(net378),
    .A2(net254),
    .B1(net198),
    .B2(net313),
    .C1(net281),
    .X(_06125_));
 sky130_fd_sc_hd__a21boi_1 _13020_ (.A1(_06527_),
    .A2(net180),
    .B1_N(net456),
    .Y(_00068_));
 sky130_fd_sc_hd__o221a_1 _13021_ (.A1(net313),
    .A2(net254),
    .B1(net198),
    .B2(\div_shifter[3] ),
    .C1(net280),
    .X(_06126_));
 sky130_fd_sc_hd__a21boi_1 _13022_ (.A1(net192),
    .A2(net180),
    .B1_N(net314),
    .Y(_00069_));
 sky130_fd_sc_hd__o221a_1 _13023_ (.A1(\div_shifter[3] ),
    .A2(net254),
    .B1(net198),
    .B2(net476),
    .C1(net280),
    .X(_06127_));
 sky130_fd_sc_hd__a21boi_1 _13024_ (.A1(_06510_),
    .A2(net180),
    .B1_N(net477),
    .Y(_00070_));
 sky130_fd_sc_hd__o221a_1 _13025_ (.A1(\div_shifter[4] ),
    .A2(net254),
    .B1(net198),
    .B2(net452),
    .C1(net280),
    .X(_06128_));
 sky130_fd_sc_hd__o21a_1 _13026_ (.A1(_06507_),
    .A2(net177),
    .B1(net453),
    .X(_00071_));
 sky130_fd_sc_hd__o221a_1 _13027_ (.A1(net452),
    .A2(net254),
    .B1(net198),
    .B2(net471),
    .C1(net280),
    .X(_06129_));
 sky130_fd_sc_hd__a21boi_1 _13028_ (.A1(_00142_),
    .A2(net180),
    .B1_N(net472),
    .Y(_00072_));
 sky130_fd_sc_hd__o221a_1 _13029_ (.A1(net471),
    .A2(net254),
    .B1(net198),
    .B2(net481),
    .C1(net280),
    .X(_06131_));
 sky130_fd_sc_hd__a21boi_1 _13030_ (.A1(net190),
    .A2(net180),
    .B1_N(net482),
    .Y(_00073_));
 sky130_fd_sc_hd__o221a_1 _13031_ (.A1(\div_shifter[7] ),
    .A2(net254),
    .B1(net198),
    .B2(net473),
    .C1(net280),
    .X(_06132_));
 sky130_fd_sc_hd__a21boi_1 _13032_ (.A1(_00166_),
    .A2(net180),
    .B1_N(net474),
    .Y(_00074_));
 sky130_fd_sc_hd__o221a_1 _13033_ (.A1(\div_shifter[8] ),
    .A2(net254),
    .B1(net198),
    .B2(net462),
    .C1(net280),
    .X(_06133_));
 sky130_fd_sc_hd__a21boi_1 _13034_ (.A1(net173),
    .A2(net181),
    .B1_N(net463),
    .Y(_00075_));
 sky130_fd_sc_hd__o221a_1 _13035_ (.A1(net462),
    .A2(net254),
    .B1(net198),
    .B2(net486),
    .C1(net280),
    .X(_06134_));
 sky130_fd_sc_hd__a21boi_1 _13036_ (.A1(_00373_),
    .A2(net181),
    .B1_N(net487),
    .Y(_00076_));
 sky130_fd_sc_hd__o221a_1 _13037_ (.A1(\div_shifter[10] ),
    .A2(net254),
    .B1(net198),
    .B2(net436),
    .C1(net281),
    .X(_06135_));
 sky130_fd_sc_hd__o21a_1 _13038_ (.A1(_00328_),
    .A2(net177),
    .B1(net437),
    .X(_00077_));
 sky130_fd_sc_hd__o221a_1 _13039_ (.A1(net436),
    .A2(net255),
    .B1(net198),
    .B2(net490),
    .C1(net280),
    .X(_06137_));
 sky130_fd_sc_hd__a21boi_1 _13040_ (.A1(_00330_),
    .A2(net181),
    .B1_N(net491),
    .Y(_00078_));
 sky130_fd_sc_hd__o221a_1 _13041_ (.A1(\div_shifter[12] ),
    .A2(net255),
    .B1(net199),
    .B2(net429),
    .C1(net281),
    .X(_06138_));
 sky130_fd_sc_hd__o21a_1 _13042_ (.A1(_00324_),
    .A2(net177),
    .B1(net430),
    .X(_00079_));
 sky130_fd_sc_hd__o221a_1 _13043_ (.A1(net429),
    .A2(net255),
    .B1(net199),
    .B2(net447),
    .C1(net280),
    .X(_06139_));
 sky130_fd_sc_hd__a21boi_1 _13044_ (.A1(_00343_),
    .A2(net181),
    .B1_N(net448),
    .Y(_00080_));
 sky130_fd_sc_hd__o221a_1 _13045_ (.A1(net447),
    .A2(net255),
    .B1(net199),
    .B2(net465),
    .C1(net280),
    .X(_06140_));
 sky130_fd_sc_hd__a21boi_1 _13046_ (.A1(net122),
    .A2(net181),
    .B1_N(net468),
    .Y(_00081_));
 sky130_fd_sc_hd__o221a_1 _13047_ (.A1(net465),
    .A2(net254),
    .B1(net198),
    .B2(net401),
    .C1(net280),
    .X(_06141_));
 sky130_fd_sc_hd__a21boi_1 _13048_ (.A1(_00265_),
    .A2(net181),
    .B1_N(net466),
    .Y(_00082_));
 sky130_fd_sc_hd__o221a_1 _13049_ (.A1(net401),
    .A2(net254),
    .B1(net198),
    .B2(net321),
    .C1(net280),
    .X(_06143_));
 sky130_fd_sc_hd__o21a_1 _13050_ (.A1(net126),
    .A2(net177),
    .B1(net402),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _13051_ (.A1(net321),
    .A2(net254),
    .B1(net198),
    .B2(\div_shifter[18] ),
    .C1(net280),
    .X(_06144_));
 sky130_fd_sc_hd__a21boi_1 _13052_ (.A1(_00305_),
    .A2(net181),
    .B1_N(net322),
    .Y(_00084_));
 sky130_fd_sc_hd__o221a_1 _13053_ (.A1(\div_shifter[18] ),
    .A2(net254),
    .B1(net198),
    .B2(net439),
    .C1(net280),
    .X(_06145_));
 sky130_fd_sc_hd__o21a_1 _13054_ (.A1(net88),
    .A2(net177),
    .B1(net440),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _13055_ (.A1(\div_shifter[19] ),
    .A2(net254),
    .B1(net199),
    .B2(net412),
    .C1(net281),
    .X(_06146_));
 sky130_fd_sc_hd__o21a_1 _13056_ (.A1(_00287_),
    .A2(net177),
    .B1(net413),
    .X(_00086_));
 sky130_fd_sc_hd__o221a_1 _13057_ (.A1(net412),
    .A2(net255),
    .B1(net199),
    .B2(net432),
    .C1(net280),
    .X(_06147_));
 sky130_fd_sc_hd__o21a_1 _13058_ (.A1(_00201_),
    .A2(net177),
    .B1(net433),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _13059_ (.A1(\div_shifter[21] ),
    .A2(net255),
    .B1(net199),
    .B2(net406),
    .C1(net281),
    .X(_06149_));
 sky130_fd_sc_hd__o21a_1 _13060_ (.A1(_00205_),
    .A2(net177),
    .B1(net407),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _13061_ (.A1(net406),
    .A2(net255),
    .B1(net199),
    .B2(net418),
    .C1(net281),
    .X(_06150_));
 sky130_fd_sc_hd__o21a_1 _13062_ (.A1(net95),
    .A2(net178),
    .B1(net419),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _13063_ (.A1(\div_shifter[23] ),
    .A2(net255),
    .B1(net199),
    .B2(net387),
    .C1(net281),
    .X(_06151_));
 sky130_fd_sc_hd__o21a_1 _13064_ (.A1(_00244_),
    .A2(net178),
    .B1(net388),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _13065_ (.A1(net387),
    .A2(net255),
    .B1(net199),
    .B2(net421),
    .C1(net281),
    .X(_06152_));
 sky130_fd_sc_hd__o21a_1 _13066_ (.A1(net89),
    .A2(net178),
    .B1(_06152_),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _13067_ (.A1(net421),
    .A2(net255),
    .B1(net199),
    .B2(net384),
    .C1(net281),
    .X(_06153_));
 sky130_fd_sc_hd__o21a_1 _13068_ (.A1(_00231_),
    .A2(net178),
    .B1(net422),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _13069_ (.A1(net384),
    .A2(net255),
    .B1(net199),
    .B2(net307),
    .C1(net281),
    .X(_06155_));
 sky130_fd_sc_hd__o21a_1 _13070_ (.A1(net93),
    .A2(net178),
    .B1(net385),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _13071_ (.A1(net307),
    .A2(net255),
    .B1(net199),
    .B2(\div_shifter[28] ),
    .C1(net281),
    .X(_06156_));
 sky130_fd_sc_hd__o21a_1 _13072_ (.A1(_00441_),
    .A2(net178),
    .B1(net308),
    .X(_00094_));
 sky130_fd_sc_hd__a221o_1 _13073_ (.A1(net339),
    .A2(net257),
    .B1(net203),
    .B2(net319),
    .C1(rst),
    .X(_06157_));
 sky130_fd_sc_hd__a21oi_1 _13074_ (.A1(net68),
    .A2(net180),
    .B1(net340),
    .Y(_00095_));
 sky130_fd_sc_hd__a221o_1 _13075_ (.A1(net319),
    .A2(net257),
    .B1(net203),
    .B2(net301),
    .C1(rst),
    .X(_06158_));
 sky130_fd_sc_hd__a21oi_1 _13076_ (.A1(_01967_),
    .A2(net180),
    .B1(net320),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _13077_ (.A1(net301),
    .A2(net257),
    .B1(rst),
    .Y(_06159_));
 sky130_fd_sc_hd__o221a_1 _13078_ (.A1(net568),
    .A2(_06440_),
    .B1(net21),
    .B2(net177),
    .C1(net302),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _13079_ (.A(net568),
    .B(net298),
    .C(net3),
    .Y(_06161_));
 sky130_fd_sc_hd__a21o_1 _13080_ (.A1(net298),
    .A2(net3),
    .B1(net568),
    .X(_06162_));
 sky130_fd_sc_hd__a32o_1 _13081_ (.A1(net257),
    .A2(_06161_),
    .A3(_06162_),
    .B1(net203),
    .B2(\div_shifter[32] ),
    .X(_06163_));
 sky130_fd_sc_hd__and2_1 _13082_ (.A(net282),
    .B(net569),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_1 _13083_ (.A(_06014_),
    .B(_06016_),
    .X(_06164_));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(\div_shifter[32] ),
    .A1(_06164_),
    .S(net3),
    .X(_06165_));
 sky130_fd_sc_hd__a22o_1 _13085_ (.A1(net560),
    .A2(net203),
    .B1(_06165_),
    .B2(net256),
    .X(_06166_));
 sky130_fd_sc_hd__and2_1 _13086_ (.A(net282),
    .B(net561),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_1 _13087_ (.A(_06012_),
    .B(_06018_),
    .Y(_06167_));
 sky130_fd_sc_hd__xnor2_1 _13088_ (.A(_06017_),
    .B(_06167_),
    .Y(_06168_));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(net560),
    .A1(_06168_),
    .S(net3),
    .X(_06170_));
 sky130_fd_sc_hd__a22o_1 _13090_ (.A1(net617),
    .A2(net203),
    .B1(_06170_),
    .B2(net256),
    .X(_06171_));
 sky130_fd_sc_hd__and2_1 _13091_ (.A(net282),
    .B(net618),
    .X(_00100_));
 sky130_fd_sc_hd__nand2_1 _13092_ (.A(_06011_),
    .B(_06020_),
    .Y(_06172_));
 sky130_fd_sc_hd__xnor2_1 _13093_ (.A(_06019_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(\div_shifter[34] ),
    .A1(_06173_),
    .S(net3),
    .X(_06174_));
 sky130_fd_sc_hd__a22o_1 _13095_ (.A1(net566),
    .A2(net203),
    .B1(_06174_),
    .B2(net256),
    .X(_06175_));
 sky130_fd_sc_hd__and2_1 _13096_ (.A(net282),
    .B(net567),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13097_ (.A(_06010_),
    .B(_06021_),
    .Y(_06176_));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(net566),
    .A1(_06176_),
    .S(net3),
    .X(_06177_));
 sky130_fd_sc_hd__a22o_1 _13099_ (.A1(net612),
    .A2(net203),
    .B1(_06177_),
    .B2(net257),
    .X(_06179_));
 sky130_fd_sc_hd__and2_1 _13100_ (.A(net282),
    .B(net613),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _13101_ (.A(_06007_),
    .B(_06022_),
    .Y(_06180_));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(\div_shifter[36] ),
    .A1(_06180_),
    .S(net3),
    .X(_06181_));
 sky130_fd_sc_hd__a22o_1 _13103_ (.A1(net588),
    .A2(net203),
    .B1(_06181_),
    .B2(net257),
    .X(_06182_));
 sky130_fd_sc_hd__and2_1 _13104_ (.A(net282),
    .B(net589),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _13105_ (.A(_06003_),
    .B(_06024_),
    .Y(_06183_));
 sky130_fd_sc_hd__xnor2_1 _13106_ (.A(_06023_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(net588),
    .A1(_06184_),
    .S(net3),
    .X(_06185_));
 sky130_fd_sc_hd__a22o_1 _13108_ (.A1(net604),
    .A2(net203),
    .B1(_06185_),
    .B2(net257),
    .X(_06186_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(net282),
    .B(net605),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _13110_ (.A(_06002_),
    .B(_06027_),
    .Y(_06188_));
 sky130_fd_sc_hd__xnor2_1 _13111_ (.A(_06025_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(net604),
    .A1(_06189_),
    .S(net2),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _13113_ (.A1(net608),
    .A2(net203),
    .B1(_06190_),
    .B2(net260),
    .X(_06191_));
 sky130_fd_sc_hd__and2_1 _13114_ (.A(net283),
    .B(_06191_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(_06001_),
    .B(_06029_),
    .Y(_06192_));
 sky130_fd_sc_hd__xnor2_1 _13116_ (.A(_06028_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\div_shifter[39] ),
    .A1(_06193_),
    .S(net2),
    .X(_06194_));
 sky130_fd_sc_hd__a22o_1 _13118_ (.A1(net578),
    .A2(net204),
    .B1(_06194_),
    .B2(net260),
    .X(_06195_));
 sky130_fd_sc_hd__and2_1 _13119_ (.A(net283),
    .B(net579),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_1 _13120_ (.A(_06000_),
    .B(_06031_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_1 _13121_ (.A(_06030_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__mux2_1 _13122_ (.A0(net578),
    .A1(_06198_),
    .S(net2),
    .X(_06199_));
 sky130_fd_sc_hd__a22o_1 _13123_ (.A1(net598),
    .A2(net204),
    .B1(_06199_),
    .B2(net260),
    .X(_06200_));
 sky130_fd_sc_hd__and2_1 _13124_ (.A(net278),
    .B(net599),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _13125_ (.A(_05999_),
    .B(_06033_),
    .Y(_06201_));
 sky130_fd_sc_hd__xnor2_1 _13126_ (.A(_06032_),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(net598),
    .A1(_06202_),
    .S(net2),
    .X(_06203_));
 sky130_fd_sc_hd__a22o_1 _13128_ (.A1(net603),
    .A2(net201),
    .B1(_06203_),
    .B2(net258),
    .X(_06204_));
 sky130_fd_sc_hd__and2_1 _13129_ (.A(net278),
    .B(_06204_),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(_05998_),
    .B(_06035_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13131_ (.A(_06034_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(\div_shifter[42] ),
    .A1(_06207_),
    .S(net1),
    .X(_06208_));
 sky130_fd_sc_hd__a22o_1 _13133_ (.A1(net600),
    .A2(net201),
    .B1(_06208_),
    .B2(net258),
    .X(_06209_));
 sky130_fd_sc_hd__and2_1 _13134_ (.A(net278),
    .B(net601),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _13135_ (.A(_05997_),
    .B(_06038_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _13136_ (.A(_06036_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__mux2_1 _13137_ (.A0(\div_shifter[43] ),
    .A1(_06211_),
    .S(net1),
    .X(_06212_));
 sky130_fd_sc_hd__a22o_1 _13138_ (.A1(net572),
    .A2(net200),
    .B1(_06212_),
    .B2(net258),
    .X(_06213_));
 sky130_fd_sc_hd__and2_1 _13139_ (.A(net275),
    .B(net573),
    .X(_00110_));
 sky130_fd_sc_hd__nand2_1 _13140_ (.A(_05996_),
    .B(_06040_),
    .Y(_06215_));
 sky130_fd_sc_hd__xnor2_1 _13141_ (.A(_06039_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(net572),
    .A1(_06216_),
    .S(net1),
    .X(_06217_));
 sky130_fd_sc_hd__a22o_1 _13143_ (.A1(net614),
    .A2(net200),
    .B1(_06217_),
    .B2(net258),
    .X(_06218_));
 sky130_fd_sc_hd__and2_1 _13144_ (.A(net275),
    .B(_06218_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _13145_ (.A(_05995_),
    .B(_06042_),
    .Y(_06219_));
 sky130_fd_sc_hd__xnor2_1 _13146_ (.A(_06041_),
    .B(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(\div_shifter[45] ),
    .A1(_06220_),
    .S(net2),
    .X(_06221_));
 sky130_fd_sc_hd__a22o_1 _13148_ (.A1(net606),
    .A2(net200),
    .B1(_06221_),
    .B2(net259),
    .X(_06222_));
 sky130_fd_sc_hd__and2_1 _13149_ (.A(net276),
    .B(net607),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _13150_ (.A(_05994_),
    .B(_06044_),
    .Y(_06224_));
 sky130_fd_sc_hd__xnor2_1 _13151_ (.A(_06043_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__mux2_1 _13152_ (.A0(\div_shifter[46] ),
    .A1(_06225_),
    .S(net1),
    .X(_06226_));
 sky130_fd_sc_hd__a22o_1 _13153_ (.A1(net592),
    .A2(net200),
    .B1(_06226_),
    .B2(net259),
    .X(_06227_));
 sky130_fd_sc_hd__and2_1 _13154_ (.A(net276),
    .B(net593),
    .X(_00113_));
 sky130_fd_sc_hd__nand2_1 _13155_ (.A(_05992_),
    .B(_06046_),
    .Y(_06228_));
 sky130_fd_sc_hd__xnor2_1 _13156_ (.A(_06045_),
    .B(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(net592),
    .A1(_06229_),
    .S(net1),
    .X(_06230_));
 sky130_fd_sc_hd__a22o_1 _13158_ (.A1(net615),
    .A2(net202),
    .B1(_06230_),
    .B2(net259),
    .X(_06231_));
 sky130_fd_sc_hd__and2_1 _13159_ (.A(net276),
    .B(_06231_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _13160_ (.A(_05991_),
    .B(_06049_),
    .Y(_06233_));
 sky130_fd_sc_hd__xnor2_1 _13161_ (.A(_06047_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__mux2_1 _13162_ (.A0(\div_shifter[48] ),
    .A1(_06234_),
    .S(net1),
    .X(_06235_));
 sky130_fd_sc_hd__a22o_1 _13163_ (.A1(net576),
    .A2(_06439_),
    .B1(_06235_),
    .B2(net259),
    .X(_06236_));
 sky130_fd_sc_hd__and2_1 _13164_ (.A(net276),
    .B(net577),
    .X(_00115_));
 sky130_fd_sc_hd__nand2b_1 _13165_ (.A_N(_05989_),
    .B(_05990_),
    .Y(_06237_));
 sky130_fd_sc_hd__xnor2_1 _13166_ (.A(_06050_),
    .B(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(net576),
    .A1(_06238_),
    .S(net1),
    .X(_06239_));
 sky130_fd_sc_hd__a22o_1 _13168_ (.A1(net590),
    .A2(net200),
    .B1(_06239_),
    .B2(net259),
    .X(_06240_));
 sky130_fd_sc_hd__and2_1 _13169_ (.A(net276),
    .B(net591),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _13170_ (.A(_05988_),
    .B(_06052_),
    .Y(_06242_));
 sky130_fd_sc_hd__xnor2_1 _13171_ (.A(_06051_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(\div_shifter[50] ),
    .A1(_06243_),
    .S(net1),
    .X(_06244_));
 sky130_fd_sc_hd__a22o_1 _13173_ (.A1(net570),
    .A2(net201),
    .B1(_06244_),
    .B2(net259),
    .X(_06245_));
 sky130_fd_sc_hd__and2_1 _13174_ (.A(net276),
    .B(net571),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13175_ (.A(_06053_),
    .B(_06055_),
    .Y(_06246_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(net570),
    .A1(_06246_),
    .S(net1),
    .X(_06247_));
 sky130_fd_sc_hd__a22o_1 _13177_ (.A1(net597),
    .A2(net201),
    .B1(_06247_),
    .B2(net259),
    .X(_06248_));
 sky130_fd_sc_hd__and2_1 _13178_ (.A(net276),
    .B(_06248_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _13179_ (.A(_05986_),
    .B(_06057_),
    .Y(_06250_));
 sky130_fd_sc_hd__xnor2_1 _13180_ (.A(_06056_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(\div_shifter[52] ),
    .A1(_06251_),
    .S(net1),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _13182_ (.A1(net594),
    .A2(net201),
    .B1(_06252_),
    .B2(net259),
    .X(_06253_));
 sky130_fd_sc_hd__and2_1 _13183_ (.A(net276),
    .B(net595),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13184_ (.A(_06058_),
    .B(_06061_),
    .Y(_06254_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(net594),
    .A1(_06254_),
    .S(net1),
    .X(_06255_));
 sky130_fd_sc_hd__a22o_1 _13186_ (.A1(net611),
    .A2(net200),
    .B1(_06255_),
    .B2(net259),
    .X(_06256_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(net276),
    .B(_06256_),
    .X(_00120_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_05984_),
    .B(_06063_),
    .Y(_06257_));
 sky130_fd_sc_hd__xnor2_1 _13189_ (.A(_06062_),
    .B(_06257_),
    .Y(_06259_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(\div_shifter[54] ),
    .A1(_06259_),
    .S(net1),
    .X(_06260_));
 sky130_fd_sc_hd__a22o_1 _13191_ (.A1(net584),
    .A2(net201),
    .B1(_06260_),
    .B2(net259),
    .X(_06261_));
 sky130_fd_sc_hd__and2_1 _13192_ (.A(net277),
    .B(net585),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13193_ (.A(_06064_),
    .B(_06066_),
    .Y(_06262_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(net584),
    .A1(_06262_),
    .S(net1),
    .X(_06263_));
 sky130_fd_sc_hd__a22o_1 _13195_ (.A1(net609),
    .A2(net201),
    .B1(_06263_),
    .B2(net259),
    .X(_06264_));
 sky130_fd_sc_hd__and2_1 _13196_ (.A(net277),
    .B(net610),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(_05981_),
    .B(_06068_),
    .Y(_06265_));
 sky130_fd_sc_hd__xnor2_1 _13198_ (.A(_06067_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(\div_shifter[56] ),
    .A1(_06266_),
    .S(net1),
    .X(_06268_));
 sky130_fd_sc_hd__a22o_1 _13200_ (.A1(net564),
    .A2(net201),
    .B1(_06268_),
    .B2(net259),
    .X(_06269_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(net277),
    .B(net565),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13202_ (.A(_05980_),
    .B(_06069_),
    .Y(_06270_));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(net564),
    .A1(_06270_),
    .S(net1),
    .X(_06271_));
 sky130_fd_sc_hd__a22o_1 _13204_ (.A1(net586),
    .A2(net201),
    .B1(_06271_),
    .B2(net259),
    .X(_06272_));
 sky130_fd_sc_hd__and2_1 _13205_ (.A(net277),
    .B(net587),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _13206_ (.A(_05977_),
    .B(_06072_),
    .Y(_06273_));
 sky130_fd_sc_hd__xnor2_1 _13207_ (.A(_06071_),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(net586),
    .A1(_06274_),
    .S(net1),
    .X(_06275_));
 sky130_fd_sc_hd__a22o_1 _13209_ (.A1(net596),
    .A2(net201),
    .B1(_06275_),
    .B2(net260),
    .X(_06277_));
 sky130_fd_sc_hd__and2_1 _13210_ (.A(net277),
    .B(_06277_),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _13211_ (.A(_06073_),
    .B(_06075_),
    .Y(_06278_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(net596),
    .A1(_06278_),
    .S(net2),
    .X(_06279_));
 sky130_fd_sc_hd__a22o_1 _13213_ (.A1(net602),
    .A2(net203),
    .B1(_06279_),
    .B2(net260),
    .X(_06280_));
 sky130_fd_sc_hd__and2_1 _13214_ (.A(net277),
    .B(_06280_),
    .X(_00126_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(_05975_),
    .B(_06077_),
    .Y(_06281_));
 sky130_fd_sc_hd__xnor2_1 _13216_ (.A(_06076_),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(\div_shifter[60] ),
    .A1(_06282_),
    .S(net2),
    .X(_06283_));
 sky130_fd_sc_hd__a22o_1 _13218_ (.A1(net582),
    .A2(net203),
    .B1(_06283_),
    .B2(net260),
    .X(_06284_));
 sky130_fd_sc_hd__and2_1 _13219_ (.A(_04448_),
    .B(net583),
    .X(_00127_));
 sky130_fd_sc_hd__xnor2_1 _13220_ (.A(_05974_),
    .B(_06078_),
    .Y(_06286_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(\div_shifter[61] ),
    .A1(_06286_),
    .S(net2),
    .X(_06287_));
 sky130_fd_sc_hd__a22o_1 _13222_ (.A1(net574),
    .A2(net203),
    .B1(_06287_),
    .B2(net260),
    .X(_06288_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(net283),
    .B(net575),
    .X(_00128_));
 sky130_fd_sc_hd__nand2b_1 _13224_ (.A_N(_06080_),
    .B(_06082_),
    .Y(_06289_));
 sky130_fd_sc_hd__a32o_1 _13225_ (.A1(net619),
    .A2(net260),
    .A3(_06289_),
    .B1(net204),
    .B2(net469),
    .X(_06290_));
 sky130_fd_sc_hd__and2_1 _13226_ (.A(net277),
    .B(net470),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _13227_ (.A(net444),
    .B(_06440_),
    .Y(_06291_));
 sky130_fd_sc_hd__o211a_1 _13228_ (.A1(net444),
    .A2(net260),
    .B1(net283),
    .C1(net445),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13229_ (.A1(net488),
    .A2(net204),
    .B1(_05923_),
    .B2(net261),
    .X(_06293_));
 sky130_fd_sc_hd__o211a_1 _13230_ (.A1(net488),
    .A2(net444),
    .B1(net283),
    .C1(_06293_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13231_ (.A1(net492),
    .A2(net204),
    .B1(net624),
    .B2(net261),
    .X(_06294_));
 sky130_fd_sc_hd__a21o_1 _13232_ (.A1(net488),
    .A2(net444),
    .B1(net492),
    .X(_06295_));
 sky130_fd_sc_hd__and3_1 _13233_ (.A(net283),
    .B(_06294_),
    .C(net498),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13234_ (.A1(net449),
    .A2(net204),
    .B1(_05926_),
    .B2(net260),
    .X(_06296_));
 sky130_fd_sc_hd__a31o_1 _13235_ (.A1(\div_counter[2] ),
    .A2(\div_counter[1] ),
    .A3(net444),
    .B1(net449),
    .X(_06297_));
 sky130_fd_sc_hd__and3_1 _13236_ (.A(net283),
    .B(_06296_),
    .C(net450),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13237_ (.A1(net296),
    .A2(net204),
    .B1(_05927_),
    .B2(net260),
    .X(_06298_));
 sky130_fd_sc_hd__o211a_1 _13238_ (.A1(net296),
    .A2(_05925_),
    .B1(_06298_),
    .C1(net283),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13239_ (.A1(net479),
    .A2(_05929_),
    .B1(net283),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00000_),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net306),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net299),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00003_),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00004_),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00005_),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00006_),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00007_),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net326),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net312),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net335),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net329),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net392),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net332),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net353),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net350),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net377),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net371),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net347),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00020_),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net356),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net383),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net362),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net374),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net398),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net405),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net417),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net395),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net368),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net411),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net426),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net365),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net359),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13274_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00035_),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00037_),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net519),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00040_),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00041_),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00042_),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net510),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00044_),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net504),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00046_),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00047_),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net531),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net507),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00051_),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00052_),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net534),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net522),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00055_),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00056_),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net496),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net501),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00059_),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net485),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net539),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00062_),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00063_),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00064_),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net459),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net380),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00068_),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net315),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net478),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net454),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00073_),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net475),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net464),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00076_),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net438),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00078_),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net431),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00080_),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00081_),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00082_),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00083_),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net323),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net441),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net414),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00087_),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net408),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net420),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net389),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net428),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net423),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net386),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net309),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00095_),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00096_),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net303),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13338_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00099_),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_2 _13340_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00129_),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net446),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net489),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00132_),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net451),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net297),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net480),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13376_ (.A(instruction[11]),
    .X(loadstore_dest[0]));
 sky130_fd_sc_hd__buf_12 _13377_ (.A(instruction[12]),
    .X(loadstore_dest[1]));
 sky130_fd_sc_hd__buf_12 _13378_ (.A(instruction[13]),
    .X(loadstore_dest[2]));
 sky130_fd_sc_hd__buf_12 _13379_ (.A(instruction[14]),
    .X(loadstore_dest[3]));
 sky130_fd_sc_hd__buf_12 _13380_ (.A(instruction[15]),
    .X(loadstore_dest[4]));
 sky130_fd_sc_hd__buf_12 _13381_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13382_ (.A(instruction[6]),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13383_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13384_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13385_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13386_ (.A(instruction[4]),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_6 fanout1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 fanout10 (.A(_01971_),
    .X(net10));
 sky130_fd_sc_hd__buf_6 fanout100 (.A(_00165_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(_00165_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(_00380_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(_00379_),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(_00361_),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_8 fanout11 (.A(_01955_),
    .X(net11));
 sky130_fd_sc_hd__buf_8 fanout110 (.A(_00310_),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(_00310_),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout113 (.A(_00298_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 fanout114 (.A(_00294_),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(_00275_),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(_01955_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 fanout120 (.A(_00271_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_16 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__buf_12 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_16 fanout123 (.A(_00264_),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_16 fanout124 (.A(_00261_),
    .X(net124));
 sky130_fd_sc_hd__buf_12 fanout125 (.A(_00260_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(_00260_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(_00212_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(_00212_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(_00197_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout13 (.A(_00689_),
    .X(net13));
 sky130_fd_sc_hd__buf_4 fanout130 (.A(_00197_),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(_00175_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(_00175_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_8 fanout134 (.A(_00169_),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_16 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(_00327_),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_16 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_12 fanout138 (.A(_00323_),
    .X(net138));
 sky130_fd_sc_hd__buf_6 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(_00249_),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(_00242_),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(_00226_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(_00151_),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(_00151_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(_00145_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(_06539_),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(_06539_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(_00678_),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(_06533_),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(_06533_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_8 fanout152 (.A(_06517_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(_06517_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_8 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(_06513_),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(net158),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(_06465_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 fanout159 (.A(_06464_),
    .X(net159));
 sky130_fd_sc_hd__buf_6 fanout16 (.A(_00399_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(_06464_),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(_06464_),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(_06464_),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(_06464_),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(_02250_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout17 (.A(_02082_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(_02249_),
    .X(net170));
 sky130_fd_sc_hd__buf_12 fanout171 (.A(net622),
    .X(net171));
 sky130_fd_sc_hd__buf_12 fanout172 (.A(_00163_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(_00163_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(_06471_),
    .X(net174));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(_06470_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(_05931_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(_05931_),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(_05930_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout18 (.A(_02082_),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_2 fanout182 (.A(_05930_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(_02335_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(_02335_),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(_02332_),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(_02322_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(_02246_),
    .X(net187));
 sky130_fd_sc_hd__buf_12 fanout188 (.A(_00140_),
    .X(net188));
 sky130_fd_sc_hd__buf_12 fanout189 (.A(_00140_),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(_00140_),
    .X(net190));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__buf_8 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_16 fanout193 (.A(_06509_),
    .X(net193));
 sky130_fd_sc_hd__buf_12 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(_06506_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_8 fanout196 (.A(_06449_),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(_06440_),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout2 (.A(net3),
    .X(net2));
 sky130_fd_sc_hd__buf_8 fanout20 (.A(_02082_),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_8 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(_06439_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 fanout203 (.A(_06439_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_06439_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net207),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(_06342_),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_8 fanout21 (.A(_02081_),
    .X(net21));
 sky130_fd_sc_hd__buf_6 fanout210 (.A(_06341_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(_06337_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(net216),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(_06331_),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(_06324_),
    .X(net218));
 sky130_fd_sc_hd__buf_6 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(net222),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(_06317_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(_06308_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(_04768_),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_2 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(_00443_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(_02516_),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(_02337_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_8 fanout233 (.A(_02329_),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(_02326_),
    .X(net234));
 sky130_fd_sc_hd__buf_2 fanout235 (.A(_02326_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(_02324_),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(_06495_),
    .X(net237));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_16 fanout239 (.A(_06469_),
    .X(net239));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(_00312_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 fanout241 (.A(_06461_),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(_06460_),
    .X(net242));
 sky130_fd_sc_hd__buf_6 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_6 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout245 (.A(_06433_),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_8 fanout246 (.A(_06433_),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(_06433_),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_16 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_6 fanout249 (.A(_06432_),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout25 (.A(_00312_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(_06307_),
    .X(net251));
 sky130_fd_sc_hd__buf_8 fanout252 (.A(_04746_),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(_04746_),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 fanout255 (.A(_04383_),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net261),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net261),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__buf_6 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(net427),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 fanout262 (.A(_06466_),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(_06466_),
    .X(net263));
 sky130_fd_sc_hd__buf_8 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(_04670_),
    .X(net265));
 sky130_fd_sc_hd__buf_8 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_16 fanout267 (.A(_04670_),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(net270),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_8 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout27 (.A(_00308_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(_04659_),
    .X(net270));
 sky130_fd_sc_hd__buf_8 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(_04648_),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(_04481_),
    .X(net273));
 sky130_fd_sc_hd__buf_2 fanout274 (.A(_04481_),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net279),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(_04448_),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(_04448_),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_8 fanout28 (.A(_00295_),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(_04448_),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout283 (.A(_04448_),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(_04438_),
    .X(net286));
 sky130_fd_sc_hd__buf_6 fanout287 (.A(_04405_),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(_04405_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_16 fanout289 (.A(reg1_val[1]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout29 (.A(_00295_),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(reg1_val[15]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(reg1_val[14]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(reg1_val[0]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_8 fanout294 (.A(instruction[7]),
    .X(net294));
 sky130_fd_sc_hd__buf_4 fanout295 (.A(instruction[7]),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout3 (.A(_06083_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 fanout31 (.A(_00290_),
    .X(net31));
 sky130_fd_sc_hd__buf_8 fanout32 (.A(_00278_),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(_00278_),
    .X(net33));
 sky130_fd_sc_hd__buf_6 fanout34 (.A(_00269_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(_00269_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_8 fanout37 (.A(_00251_),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_8 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_8 fanout39 (.A(_00247_),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout4 (.A(net5),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_6 fanout41 (.A(_00236_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_8 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_6 fanout43 (.A(_00234_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(_00214_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_8 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_6 fanout47 (.A(_00208_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_16 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_12 fanout49 (.A(_00202_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(_02084_),
    .X(net5));
 sky130_fd_sc_hd__buf_6 fanout50 (.A(_00156_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(_00156_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_8 fanout52 (.A(_00149_),
    .X(net52));
 sky130_fd_sc_hd__buf_4 fanout53 (.A(_00149_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(_06552_),
    .X(net55));
 sky130_fd_sc_hd__buf_8 fanout56 (.A(_06537_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_06537_),
    .X(net57));
 sky130_fd_sc_hd__buf_8 fanout58 (.A(_06535_),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(_06535_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 fanout6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(_06521_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_06521_),
    .X(net61));
 sky130_fd_sc_hd__buf_8 fanout62 (.A(_06516_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(_06516_),
    .X(net63));
 sky130_fd_sc_hd__buf_8 fanout64 (.A(_06499_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(_06499_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(_06493_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_16 fanout68 (.A(net70),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_6 fanout7 (.A(_02070_),
    .X(net7));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(_00669_),
    .X(net70));
 sky130_fd_sc_hd__buf_8 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_6 fanout72 (.A(_00351_),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(_00349_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_8 fanout76 (.A(_00348_),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(_00346_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(_00339_),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_8 fanout82 (.A(_00336_),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(_00335_),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(_00333_),
    .X(net86));
 sky130_fd_sc_hd__buf_12 fanout87 (.A(_00286_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 fanout88 (.A(_00286_),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_8 fanout91 (.A(_00230_),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_8 fanout94 (.A(_00223_),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_00193_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_12 fanout97 (.A(_00193_),
    .X(net97));
 sky130_fd_sc_hd__buf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(_00173_),
    .X(net99));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1 (.A(\div_counter[4] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_05932_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00028_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\divi2_l[23] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_05961_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_00025_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\divi2_l[4] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_05938_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\div_shifter[16] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_06143_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\divi2_l[24] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_05962_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_00001_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_00026_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\div_shifter[22] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_06149_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_00088_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\divi2_l[28] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_05967_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_00030_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\div_shifter[20] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_06146_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_00086_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\div_shifter[27] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\divi2_l[25] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_05963_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_00027_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\div_shifter[23] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_06150_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00089_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\div_shifter[25] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_06153_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_00092_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\divi2_l[29] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_06156_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_05968_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_00031_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(busy_l),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_00091_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\div_shifter[13] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_06138_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00079_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\div_shifter[21] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_06147_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\divi2_l[18] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00094_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_05955_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\div_shifter[11] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_06135_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_00077_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\div_shifter[19] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_06145_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_00085_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\div_shifter[0] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_06122_),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 hold149 (.A(net623),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\divi2_l[8] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_06291_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_00130_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\div_shifter[14] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_06139_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\div_counter[3] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_06297_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00133_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\div_shifter[5] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06128_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_00071_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_05943_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\div_shifter[2] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_06125_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\div_res[31] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_06121_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_00065_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\divi2_l[1] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_05934_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\div_shifter[9] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_06133_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_00075_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_00010_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net467),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_06141_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\div_shifter[15] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_06140_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\div_shifter[63] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_06290_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\div_shifter[6] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_06129_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\div_shifter[8] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_06132_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net455),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_00074_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\div_shifter[4] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_06127_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_00070_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(div_complete),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_00135_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\div_shifter[7] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_06131_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\div_res[25] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_06115_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_06126_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_00060_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\div_shifter[10] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_06134_),
    .X(net487));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold193 (.A(\div_counter[1] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_00131_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\div_shifter[12] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_06137_),
    .X(net491));
 sky130_fd_sc_hd__buf_1 hold197 (.A(net497),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_05927_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\div_res[22] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00134_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00069_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_06111_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_00057_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\div_counter[2] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_06295_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\div_res[23] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_06113_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_00058_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\div_res[11] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_06097_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_00045_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\divi2_l[5] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\div_res[15] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_06102_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_00049_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\div_res[9] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_06095_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_00043_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\div_res[17] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_06104_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net544),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_06110_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_05939_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\div_res[12] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_06098_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\div_res[5] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_06090_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_00039_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\div_res[20] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_06108_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_00054_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\div_res[24] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_06114_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\div_shifter[29] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\div_res[3] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_06087_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\div_res[6] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_06091_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\div_res[14] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_06101_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_00048_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\div_res[19] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_06107_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_00053_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_04361_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\div_res[10] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_06096_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\div_res[27] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_06116_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_00061_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\div_res[16] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_06103_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\div_res[7] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_06092_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\div_res[21] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_06158_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_06109_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\div_res[28] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_06117_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\div_res[29] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_06119_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\div_res[18] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_06105_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\div_res[8] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_06093_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\div_res[13] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\div_shifter[17] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_06099_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\div_res[4] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_06089_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\div_res[30] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_06120_),
    .X(net559));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold265 (.A(\div_shifter[33] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_06166_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\div_res[2] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_06086_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\div_shifter[57] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_06144_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_06269_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\div_shifter[35] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_06175_),
    .X(net567));
 sky130_fd_sc_hd__buf_1 hold273 (.A(\div_shifter[31] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_06163_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\div_shifter[51] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_06245_),
    .X(net571));
 sky130_fd_sc_hd__buf_1 hold277 (.A(net626),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_06213_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\div_shifter[62] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00084_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_06288_),
    .X(net575));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold281 (.A(\div_shifter[49] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_06236_),
    .X(net577));
 sky130_fd_sc_hd__buf_1 hold283 (.A(\div_shifter[40] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_06195_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\div_res[1] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_06085_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[61] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_06284_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\div_shifter[55] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\divi2_l[7] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_06261_),
    .X(net585));
 sky130_fd_sc_hd__buf_1 hold291 (.A(net625),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_06272_),
    .X(net587));
 sky130_fd_sc_hd__buf_1 hold293 (.A(\div_shifter[37] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_06182_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\div_shifter[50] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_06240_),
    .X(net591));
 sky130_fd_sc_hd__buf_1 hold297 (.A(net627),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_06227_),
    .X(net593));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold299 (.A(\div_shifter[53] ),
    .X(net594));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\divi2_l[0] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_05942_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_06253_),
    .X(net595));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold301 (.A(\div_shifter[59] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\div_shifter[52] ),
    .X(net597));
 sky130_fd_sc_hd__buf_1 hold303 (.A(\div_shifter[41] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_06200_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\div_shifter[43] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_06209_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\div_shifter[60] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\div_shifter[42] ),
    .X(net603));
 sky130_fd_sc_hd__buf_1 hold309 (.A(\div_shifter[38] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_00009_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_06186_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\div_shifter[46] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_06222_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\div_shifter[39] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\div_shifter[56] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_06264_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\div_shifter[54] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\div_shifter[36] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_06179_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\div_shifter[45] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\divi2_l[10] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\div_shifter[48] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\div_res[0] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\div_shifter[34] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_06171_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\div_shifter[62] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\div_res[2] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\div_res[16] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\div_counter[0] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_05924_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\div_shifter[58] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_05945_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\div_shifter[44] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\div_shifter[47] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_00012_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\divi2_l[12] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_05948_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_00014_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\divi2_l[9] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_05944_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00002_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_00011_),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\divi2_l[6] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_05940_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\div_shifter[28] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_04372_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_06157_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\divi2_l[2] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_05936_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\divi2_l[3] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_05937_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\div_shifter[30] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\divi2_l[17] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_05954_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_00019_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\divi2_l[14] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_05950_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_00016_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\divi2_l[13] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_05949_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00015_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\divi2_l[19] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_04350_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_05956_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_00021_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\divi2_l[31] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_05970_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_00033_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\divi2_l[21] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_05958_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_00023_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\divi2_l[30] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_05969_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_06159_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_00032_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\divi2_l[27] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_05966_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_00029_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\divi2_l[16] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_05952_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_00018_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\divi2_l[22] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_05960_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_00024_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00097_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\divi2_l[15] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_05951_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_00017_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\div_shifter[1] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_06123_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_00067_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\divi2_l[20] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_05957_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_00022_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\div_shifter[26] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(divi1_sign),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_06155_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_00093_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\div_shifter[24] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_06151_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00090_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\divi2_l[11] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_05946_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_00013_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\divi2_l[26] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_05964_),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_8 load_slew1 (.A(_00163_),
    .X(net622));
 sky130_fd_sc_hd__buf_4 max_cap102 (.A(_00164_),
    .X(net102));
 sky130_fd_sc_hd__buf_4 max_cap109 (.A(_00314_),
    .X(net109));
 sky130_fd_sc_hd__buf_6 max_cap112 (.A(_00299_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 max_cap115 (.A(_00276_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_8 max_cap117 (.A(_00275_),
    .X(net117));
 sky130_fd_sc_hd__buf_6 max_cap118 (.A(_00272_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 max_cap139 (.A(_00297_),
    .X(net139));
 sky130_fd_sc_hd__buf_4 max_cap197 (.A(_06448_),
    .X(net197));
 sky130_fd_sc_hd__buf_4 max_cap219 (.A(_06323_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 max_cap240 (.A(_06468_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_8 wire8 (.A(_02069_),
    .X(net8));
endmodule

